* NGSPICE file created from OQPSK_RCOSINE_ALL.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 D SETN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latrnq_1 D E RN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

.subckt OQPSK_RCOSINE_ALL ACK Bit_In EN I[0] I[10] I[11] I[12] I[1] I[2] I[3] I[4]
+ I[5] I[6] I[7] I[8] I[9] Q[0] Q[10] Q[11] Q[12] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7]
+ Q[8] Q[9] REQ_SAMPLE RST addI[0] addI[1] addI[2] addI[3] addI[4] addI[5] addQ[0]
+ addQ[1] addQ[2] addQ[3] addQ[4] addQ[5] vdd vss
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2106_ _1173_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1997__C _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2037_ _1071_ _1074_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2706__A1 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2182__A2 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2237__A3 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1996__A2 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2173__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1684__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1389__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1987__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1739__A2 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2724_ gen_sym.Reg_2M.data_in net52 net45 gen_sym.Reg_Sym.data_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2655_ _0439_ _0442_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1606_ p_shaping_Q.p_shaping_I.bit_in_2 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2586_ _0228_ _0146_ _0209_ _0331_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1537_ _0590_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_59_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1468_ _0548_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1399_ net51 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2683__I _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1978__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2351__C _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2440_ _0041_ _0209_ _0208_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2371_ _1319_ _1318_ _0055_ _0058_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__1672__I p_shaping_Q.p_shaping_I.bit_in_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2621__A3 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2385__A2 _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2707_ _0783_ net63 net3 _0864_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2638_ _0172_ _0516_ _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2569_ _0299_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1896__A1 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2073__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1820__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2128__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1940_ _0900_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1811__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1871_ _0943_ _0946_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2423_ _0160_ _0104_ _0142_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1878__A1 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2354_ _0119_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2285_ _0044_ _0045_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2166__C _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2055__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1802__A1 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2358__A2 _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1869__A1 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2530__A2 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2349__A2 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2521__A2 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2070_ _0521_ _1139_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2267__B _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2285__A1 _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1923_ _0907_ _0851_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1397__I _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1854_ _0929_ _0926_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1785_ _0700_ _0731_ _0861_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2406_ _0167_ _0175_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2337_ _0291_ _1330_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2268_ _1332_ _1340_ _0022_ _0026_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_55_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2276__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2733__CLK net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2199_ _1247_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2028__A1 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2579__A2 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2267__A1 _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2019__A1 p_shaping_Q.p_shaping_I.bit_in_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2106__I _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1570_ _0562_ _0591_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1950__B1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1680__I _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2122_ _0215_ _1161_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2053_ _1101_ _1123_ _1030_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1906_ _0977_ _0523_ _0980_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2430__A1 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1837_ _0909_ _0911_ _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1768_ _0706_ _0810_ _0699_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1699_ _0548_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2725__RN net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2249__A1 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1472__A2 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2421__A1 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput31 net31 Q[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput20 net20 Q[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput42 net42 addQ[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput7 net7 I[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2488__A1 _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2740_ _0015_ net52 net64 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__1766__A3 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2280__B _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2671_ _0453_ _0454_ _0457_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1622_ _0618_ _0698_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1553_ _0612_ _0623_ _0632_ _0633_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1484_ _0564_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2439__C _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2105_ _1172_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2036_ _1097_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_fanout49_I _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2651__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2706__A2 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1905__B1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1684__A2 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2633__A1 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2397__B1 _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2723_ _0007_ net56 net49 p_shaping_Q.p_shaping_I.counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2654_ _0415_ _0441_ _0412_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2585_ _0183_ _0515_ _0367_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1605_ _0683_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1536_ _0591_ _0600_ _0376_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1911__A3 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1467_ _0418_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1398_ _0355_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2019_ p_shaping_Q.p_shaping_I.bit_in_1 _1089_ _1090_ _0834_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__2624__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1363__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2370_ _1273_ _0126_ _0130_ _0136_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_37_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1657__A2 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1409__A2 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2706_ net48 _0784_ _0472_ _0486_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2637_ _0172_ _0289_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2568_ _0348_ _0349_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1896__A2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2499_ _0250_ _0275_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1519_ _0535_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1648__A2 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2553__B _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1811__A2 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1870_ _0944_ _0945_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2422_ _0162_ _0192_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2353_ _0150_ _0117_ _1204_ _1164_ _1294_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2284_ _1259_ _1305_ _1293_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2463__B _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1802__A2 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2182__C _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1999_ _1022_ _1029_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1869__A2 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2046__A2 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1922_ _0995_ _0996_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1853_ _0680_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1784_ _0860_ _0742_ _0674_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2405_ _0169_ _0170_ _0171_ _0174_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2336_ _0512_ _0097_ _0098_ _0099_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2267_ _0023_ _0024_ _1339_ _0025_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_37_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2198_ _1265_ _1272_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2028__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2193__B _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1787__A1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2368__B _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2267__A2 _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2019__A2 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1498__I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1950__B2 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1950__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1702__A1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2121_ _1189_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2052_ _1099_ _0688_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2258__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1769__A1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1905_ _0948_ _0484_ _0979_ _0924_ _0943_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__2430__A2 _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1836_ _0807_ _0852_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1767_ _0663_ _0777_ _0666_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2194__A1 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1941__A1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1698_ _0773_ _0774_ _0775_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2497__A2 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2319_ _1206_ _1207_ _1281_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1820__B _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2421__A2 _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput21 net21 Q[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput32 net32 addI[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput8 net8 I[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput43 net43 addQ[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput10 net10 I[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1766__A4 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2670_ _0445_ _0452_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1621_ _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2176__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2723__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1923__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1552_ _0561_ _0630_ _0397_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__1691__I _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1483_ _0545_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input3_I EN vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2104_ _1181_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2035_ _1098_ _1105_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2455__C _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1819_ _0753_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2706__A3 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1920__A4 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2330__A1 _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2556__B _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2275__C _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2633__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2722_ _0006_ net56 net49 p_shaping_Q.p_shaping_I.counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2653_ _0378_ _0380_ _0411_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2584_ _0288_ _0366_ _0183_ _0515_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1604_ net44 _0635_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1635__B _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1535_ _0547_ _0615_ _0555_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1466_ _0546_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2321__A1 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1397_ _0387_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout61_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2018_ _0875_ _0965_ _1089_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2624__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1596__I _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2388__B2 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2560__A1 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output42_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2130__I _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2551__A1 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2303__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2286__B p_shaping_I.p_shaping_I.bit_in vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2705_ _0883_ _0470_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2636_ _0062_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2567_ _0308_ _0310_ _0347_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__1896__A3 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2498_ _0252_ _0258_ _0273_ _0253_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_1518_ _0583_ _0567_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1449_ p_shaping_Q.p_shaping_I.counter\[1\] _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1812__C _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2196__B _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2421_ _0178_ _0191_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2352_ _1341_ _1276_ _1178_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1913__B _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1878__A3 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2283_ _0034_ _0035_ _0039_ _0042_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1998_ _1064_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1566__A2 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2619_ _0232_ _0279_ _0403_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2515__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1493__A1 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1921_ _0982_ _0983_ _0994_ _0532_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1796__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1852_ _0810_ _0654_ _0896_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1908__B _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1783_ _0721_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2404_ _0173_ _0023_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2335_ _0087_ _0075_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2266_ _0043_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2197_ _1239_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1787__A2 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1553__B _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2368__C _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1728__B _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1463__B _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2120_ _1236_ _1181_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2051_ _1121_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1904_ _0701_ _0593_ _0978_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_30_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1835_ _0907_ _0851_ _0838_ _0849_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_1766_ _0820_ _0843_ _0628_ _0681_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2313__I _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2718__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2194__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1941__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1697_ _0737_ _0749_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_66_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2318_ _1246_ _0078_ _0079_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2249_ _0508_ _0517_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput33 net33 addI[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput11 net11 I[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput9 net9 I[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput22 net22 Q[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1620_ _0699_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2176__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1551_ _0624_ _0627_ _0628_ _0631_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1482_ _0562_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2103_ _1165_ _1168_ _1169_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2509__S _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2034_ _1065_ _1101_ _1104_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_35_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1439__A1 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1818_ _0523_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1749_ _0819_ _0824_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__1678__A1 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1831__B _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1850__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1602__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1905__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1669__A1 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2330__A2 _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2721_ _0021_ _0497_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2397__A2 _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2652_ _0435_ _0438_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2583_ _0266_ _0251_ _0364_ _0147_ _0267_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1603_ _0648_ _0668_ _0675_ _0682_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1534_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1465_ _0545_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1396_ _0344_ _0365_ _0376_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_67_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2321__A2 _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2609__B1 _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout54_I net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2017_ _1084_ _1060_ _1087_ _1088_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_42_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2624__A3 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1832__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2388__A2 _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2411__I _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2704_ _0485_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2635_ _0394_ _0282_ _0402_ _0419_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__1646__B _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2566_ _0308_ _0310_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2497_ _0252_ _0258_ _0271_ _0253_ _0273_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1517_ _0539_ _0597_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1448_ _0529_ net49 _1448_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1379_ _0194_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2058__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2230__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2297__A1 _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2049__A1 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2221__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1980__B1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2141__I _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2420_ _0180_ _0190_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2351_ _0114_ _1237_ _1337_ _0115_ _1195_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_2282_ _1164_ _0040_ _1238_ _1163_ _0041_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__2288__A1 _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2460__A1 _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1997_ _1065_ _1068_ _1069_ _0532_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2618_ _0294_ _0401_ _0402_ _0394_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__2515__A2 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2549_ _0082_ _0165_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2279__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2451__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2203__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2506__A2 _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1493__A2 _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2136__I _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1920_ _0531_ _0982_ _0983_ _0994_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1851_ _0705_ _0612_ _0924_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1782_ _0612_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1924__B _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2403_ _0128_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2334_ _0077_ _0084_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2737__RN net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2265_ _1341_ _0258_ _1229_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2196_ _1269_ _1270_ _1271_ _1217_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1834__B _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1553__C _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2672__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1475__A2 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2424__A1 _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2050_ _1118_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1903_ _0674_ _0779_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1834_ _0910_ _0908_ _0873_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1765_ _0789_ _0592_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1696_ _0767_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2351__B1 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2317_ _1281_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2248_ _1328_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2179_ _1165_ _1250_ _1251_ _1252_ _1253_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_38_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2504__I _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput23 net23 Q[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput12 net12 I[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 addI[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2645__B2 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2645__A1 _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1448__A2 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1550_ _0629_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1384__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1481_ _0500_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2102_ _1162_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1687__A2 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2736__D p_shaping_I.p_shaping_I.bit_in vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2033_ _1101_ _1104_ _1030_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1439__A2 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1817_ _0634_ _0683_ _0746_ _0848_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__1375__A1 _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1748_ _0814_ _0815_ _0825_ _0641_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1679_ _0560_ _0579_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1678__A2 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1403__I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1850__A2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1905__A3 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2144__I _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2720_ _0218_ p_shaping_I.p_shaping_I.counter\[0\] _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2651_ _0400_ _0436_ _0437_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1602_ _0571_ _0677_ _0679_ _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2582_ _0205_ _1177_ _0268_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1533_ _0468_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1464_ net38 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1395_ net51 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2321__A3 _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2609__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2016_ _1031_ _0569_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_23_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout47_I _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1823__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1587__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1511__A1 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2703_ _0863_ _0469_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2634_ _0394_ _0402_ _0419_ _0281_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2565_ _0328_ _0346_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1516_ _0533_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2496_ _0272_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1447_ _0529_ net45 _1447_/ZN vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1378_ _1268_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1805__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2518__B1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2049__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2221__A2 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1980__B2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2350_ _1190_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2281_ _0065_ _0118_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1996_ _1065_ _0880_ _1030_ _1068_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2617_ _0292_ _0331_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2548_ _1212_ _0313_ _0327_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__1723__A1 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2479_ _0089_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2279__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2203__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1962__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2690__A2 _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2442__A2 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1850_ _0676_ _0925_ _0568_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1781_ _0799_ _0856_ _0857_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2402_ _1202_ _0057_ _0147_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2333_ _0093_ _0095_ _1210_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2264_ _1255_ _1174_ _1333_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2195_ _1312_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1979_ _1050_ _0698_ _1051_ _0984_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1944__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1944__B2 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1850__B _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2424__A2 _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1702__A4 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1902_ _0976_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1833_ _0906_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2179__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2179__B2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1764_ _0793_ _0673_ _0691_ _0692_ _0758_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__2610__I _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1695_ _0737_ _0749_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2351__A1 _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2316_ _1244_ _1266_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2351__B2 _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2247_ _1211_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2103__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2178_ _0065_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1917__A1 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput13 net13 I[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput24 net24 Q[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2590__A1 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput35 net35 addI[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2342__A1 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1480_ _0560_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2101_ _1167_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2032_ _1099_ _1103_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1816_ _0833_ _0891_ _0892_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1665__B _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1747_ _0819_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1678_ _0552_ _0333_ _0678_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1575__B _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2650_ _0405_ _0409_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1601_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2581_ _0356_ _0362_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1532_ _0584_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1463_ _0537_ _0540_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input1_I ACK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2747__D _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1394_ _0355_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1504__I _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2015_ _1085_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2545__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1899__A3 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2536__A1 _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2536__B2 _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2583__C _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2155__I _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2702_ _0479_ _0483_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2633_ _0316_ _0321_ _0272_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2564_ _0338_ _0345_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1515_ _0562_ _0564_ _0365_ _0376_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_59_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2495_ _1197_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1750__A2 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1446_ _0514_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1377_ _0032_ _0172_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2518__A1 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1741__A2 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output40_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1980__A2 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2280_ _1220_ _1231_ _0248_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1995_ _1031_ _1066_ _1067_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2616_ _0219_ _0272_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2547_ _0314_ _0325_ _0326_ _0203_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2478_ _0079_ _0090_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1723__A2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1429_ _0515_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1567__C _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1411__A1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1714__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1803__S _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2690__A3 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1650__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1780_ _0751_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1953__A2 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2401_ _1273_ _1238_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2332_ _0094_ _1282_ _1285_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2263_ _1342_ _1343_ _1295_ _1344_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_1_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2194_ _1190_ _1266_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1978_ _0810_ _0791_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1880__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1901_ _0894_ _0904_ _0940_ _0522_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1832_ _0873_ _0906_ _0908_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_30_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1763_ _0650_ _0739_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1926__A2 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1694_ _0639_ _0712_ _0770_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2315_ _0076_ _1270_ _1199_ _1222_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2351__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2246_ _1291_ _1325_ _1326_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2338__I _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2177_ _1162_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput25 net25 Q[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput14 net14 I[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput36 net36 addI[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2342__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1605__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2030__A1 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1384__A3 _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2100_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2031_ _0588_ _1102_ _0937_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2097__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1815_ _0835_ _0874_ _0890_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2021__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1746_ _0822_ _0823_ _0703_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1677_ _0669_ _0586_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2229_ _1307_ _1259_ _1305_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2088__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1835__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2260__A1 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2315__A2 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1826__B2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1600_ _0533_ _0579_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2580_ _0314_ _0360_ _0361_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1357__A3 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1531_ _0539_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1462_ _0542_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1393_ net41 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2014_ _1032_ _0588_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1520__I _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1729_ _0799_ _0805_ _0806_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_58_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2701_ _0390_ _0480_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2632_ _0417_ net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2563_ _0289_ _0343_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1735__B1 _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1514_ _0590_ _0592_ _0594_ _0560_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_4_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2494_ _0266_ _0267_ _0270_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1445_ _0528_ gen_sym.Reg_2M.enable vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1376_ _0085_ _0161_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2463__A1 _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1741__A3 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1425__I _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2256__I _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout60 net62 net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2693__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1994_ _0568_ _1014_ _1032_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2615_ _0396_ _0399_ _0356_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2546_ _0512_ _0325_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2477_ _1342_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1428_ _0508_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1487__A2 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1359_ net36 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2436__A1 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2690__A4 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1774__B _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2400_ _1271_ _0168_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2331_ _0025_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2262_ _1226_ _1190_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2193_ _1206_ _1266_ _1267_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2418__A1 _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1977_ _0883_ _0887_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2529_ _0307_ net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2409__A1 _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1632__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1900_ _0833_ _0973_ _0974_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_15_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1831_ _0907_ _0851_ _0893_ _0905_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_30_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1762_ _0746_ _0747_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1693_ _0716_ _0768_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2314_ _1202_ _0057_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2639__A1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2245_ _1309_ _1321_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2176_ _1218_ _1158_ _0043_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1862__A2 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1917__A3 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput15 net15 I[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput37 net37 addI[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput26 net26 Q[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2342__A3 _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1550__A1 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2529__I _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2030__A2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1608__I _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1541__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2030_ _0887_ _0692_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2097__A2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2174__I _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1814_ _0835_ _0875_ _0890_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2021__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1745_ _0790_ _0791_ _0779_ _0604_ _0699_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_7_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1375__A4 _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1962__B _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1676_ _0550_ _0549_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1681__C _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2228_ p_shaping_I.p_shaping_I.bit_in_2 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2159_ _1220_ _1231_ _1173_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2743__SETN net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1599__A1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2260__A2 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1428__I _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2208__B _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1530_ _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1762__A1 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1461_ _0541_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1392_ net39 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1801__I _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2013_ _0783_ _0784_ _0925_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1817__A2 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2632__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1728_ _0799_ _0805_ _0530_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1659_ _0726_ _0673_ _0727_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2481__A2 _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2542__I _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2698__B _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1621__I _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2472__A2 _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2224__A2 _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2700_ _0479_ _0482_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1983__A1 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2631_ _0413_ _0416_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2562_ _0161_ _1270_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1735__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1735__B2 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1513_ _0536_ _0593_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2493_ _0268_ _0254_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1444_ _0291_ net48 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1375_ _0096_ _0107_ _0118_ _0150_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_67_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout45_I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2463__A2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1687__B p_shaping_Q.p_shaping_I.counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1974__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1706__I _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout61 net62 net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout50 net42 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__2205__C _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2447__I _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2693__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1993_ _0695_ _0627_ _0938_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2614_ _0087_ _0398_ _0203_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1708__A1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2381__A1 _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2545_ _1332_ _0315_ _0320_ _0324_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2476_ _1338_ _0089_ _0220_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1427_ net53 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1358_ _1225_ _1290_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2436__A2 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2092__I _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1436__I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1938__A1 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2363__A1 _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1346__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2330_ _0074_ _0092_ _0034_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2363__B2 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2261_ _1275_ _1249_ _0194_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2192_ _1221_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2177__I _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1874__B1 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2418__A2 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2126__B _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1976_ _0728_ _1048_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2528_ _0303_ _0306_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2459_ _0232_ _0176_ _0163_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2409__A2 _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2593__A1 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2345__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1830_ _0607_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1761_ p_shaping_Q.p_shaping_I.bit_in _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1692_ _0716_ _0768_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2313_ _0027_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2244_ _1309_ _1321_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2175_ _1225_ _1249_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1959_ _0985_ _0886_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2575__A1 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput38 net38 addQ[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2327__A1 _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput16 net16 I[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput27 net27 Q[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_29_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2318__A1 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1624__I _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1541__A2 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1813_ _0876_ _0880_ _0882_ _0759_ _0889_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__2557__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2190__I _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2021__A3 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1744_ _0820_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2309__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1675_ _0613_ _0645_ _0571_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2227_ _1293_ _1259_ _1305_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_53_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2158_ _1175_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_38_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2089_ _1156_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1599__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2548__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1771__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2208__C _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1460_ _0468_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1354__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1391_ _0322_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2711__A1 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1514__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2012_ _0876_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1817__A3 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1727_ _0686_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1658_ _0609_ _0736_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2702__A1 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1589_ _0542_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2044__B _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1441__A1 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2224__A3 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1432__A1 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1983__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2630_ _0414_ _0415_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1793__B _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2561_ _0339_ _1228_ _0341_ _0181_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1735__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2492_ _0207_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2742__SETN net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1512_ _0344_ _0376_ _0365_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_4_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1443_ _0527_ gen_sym.Reg_2M.data_in vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1374_ _0129_ _0140_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1974__A2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2151__A2 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1662__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout62 net5 net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout51 net40 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2142__A2 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1653__A1 _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1992_ _0857_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1405__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2613_ _0390_ _0393_ _0395_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1708__A2 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2544_ _0321_ _0323_ _0269_ _0250_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2381__A2 _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2475_ _0181_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1426_ _0512_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1357_ _1247_ _1268_ _1279_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2133__A2 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1644__A1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2372__A2 _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1452__I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1938__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2363__A2 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2260_ _1341_ _1188_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2115__A2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2191_ _1163_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1874__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2407__B _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1975_ _0695_ _0677_ _0843_ _1047_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2527_ _0304_ _0305_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2458_ _0231_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1409_ _0450_ _0387_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2389_ _0075_ _0098_ _0511_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1865__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1617__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2290__A1 _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2042__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2345__A2 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2281__A1 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1760_ _0834_ _0836_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2584__A2 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1691_ _0769_ net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2336__A2 _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2312_ _0072_ _0068_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2639__A3 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2243_ _1263_ _1264_ _1322_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2174_ _1279_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2272__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2024__A1 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1958_ _0985_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1889_ _0964_ net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput39 net39 addQ[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput28 net28 Q[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput17 net17 I[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2327__A2 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2098__I _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1730__I _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1829__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1812_ _0883_ _0885_ _0886_ _0888_ _0728_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_30_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1743_ _0789_ _0592_ _0699_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2557__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1674_ _0561_ _0580_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2226_ _1295_ _1296_ _1300_ _1199_ _1304_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA_fanout68_I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1835__A4 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2157_ _1226_ _1228_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2088_ _0639_ _0712_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2330__B _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1508__B1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1460__I _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2236__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2539__A2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1390_ _0311_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2011_ _1064_ _1070_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1370__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1817__A4 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output9_I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1726_ _0577_ _0803_ _0765_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1657_ _0718_ _0734_ _0735_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1588_ _0534_ _0618_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2209_ _1273_ _1282_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2218__A1 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1441__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2209__A1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2235__B _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2560_ _0207_ _0340_ _0024_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2491_ _0228_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1511_ _0591_ _0585_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_4_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1442_ net3 net2 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_67_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1373_ net34 _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1709_ _0628_ _0681_ _0730_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1726__A3 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2689_ net47 _0056_ _0472_ _0473_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_48_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2439__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1662__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2611__A1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout63 net68 net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout52 net54 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1894__B _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1991_ _1058_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1405__A2 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2612_ _0390_ _0393_ _0395_ _0314_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2543_ _0182_ _0251_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2474_ _0249_ net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1425_ _0511_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1356_ _1181_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1892__A2 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout50_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1644__A2 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1580__A1 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2060__A2 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2190_ _0074_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1874__A2 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2474__I _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1974_ _0703_ _0925_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2526_ _0193_ _0196_ _0197_ _0199_ _0202_ _0245_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
X_2457_ _1307_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1408_ net43 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2388_ _0146_ _0149_ _0152_ _1332_ _0155_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1865__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2290__A2 _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2294__I _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1792__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1690_ _0713_ _0716_ _0768_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2311_ _0062_ _0046_ _0060_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1373__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1544__A1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2242_ _1291_ _1309_ _1321_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_65_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2173_ _1178_ _1227_ _1246_ _1180_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2272__A2 _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1957_ _0719_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1888_ _0961_ _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput29 net29 Q[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput18 net18 I[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2379__I _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2509_ _0187_ _0286_ _0094_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1535__A1 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2328__B _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2263__A2 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1458__I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1811_ _0809_ _0887_ _0884_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1742_ _0721_ _0663_ _0742_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1673_ _0750_ _0709_ _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2225_ _1302_ _1303_ _1194_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2156_ _1180_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2087_ _1150_ _1152_ _1155_ _1114_ _0907_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_53_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1508__B2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2181__A1 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2484__A2 _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1897__B _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2236__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1747__A1 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2010_ _1058_ _1063_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1986__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1738__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1725_ _0703_ _0801_ _0707_ _0598_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_7_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1656_ _0606_ _0649_ _0659_ _0520_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_1587_ _0663_ _0665_ _0666_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2163__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2208_ _1267_ _1283_ _1284_ _1229_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2139_ _1183_ _1196_ _1200_ _1209_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2218__A2 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1977__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2325__C _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1729__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1901__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2490_ _0182_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1510_ _0545_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1441_ _0521_ _0505_ _0526_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2145__A1 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2696__A2 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1372_ net33 _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1381__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2448__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2384__A1 _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2161__B _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1708_ _0618_ _0785_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2688_ _0266_ _0472_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1639_ _0506_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_58_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2439__A2 _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1662__A3 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout64 net68 net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout53 net54 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2611__A2 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1894__C _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1653__A3 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1990_ _0523_ _0504_ _0977_ _1062_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2611_ _0394_ _0366_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2366__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2542_ _0267_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2473_ _0202_ _0245_ _0247_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1424_ p_shaping_I.p_shaping_I.bit_in_1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1355_ _1258_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1644__A3 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1580__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2596__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1571__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2520__A1 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1973_ _1046_ net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2490__I _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2525_ _0202_ _0245_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2456_ _0223_ _0229_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__1562__A2 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1407_ _0440_ _0484_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2387_ _1278_ _1283_ _0153_ _0154_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1945__S _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1553__A2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1792__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2310_ _1324_ _0066_ _0070_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2241_ _1318_ _1320_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_2_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2172_ _1231_ _0237_ _1235_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1603__B _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2434__B _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1956_ _0993_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1887_ _0915_ _0920_ _0962_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput19 net19 Q[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2508_ _1182_ _0188_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1535__A2 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2439_ _1338_ _0151_ _1280_ _0173_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_56_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1675__S _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1526__A2 p_shaping_Q.p_shaping_I.counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1810_ _0794_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1741_ _0689_ _0628_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_7_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1765__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1672_ p_shaping_Q.p_shaping_I.bit_in_2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2714__A1 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2224_ _1221_ _0248_ _1158_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2155_ _1227_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2086_ _1153_ _1154_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1939_ _0885_ _0791_ _1012_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2705__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1508__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2181__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2484__A3 _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1444__A1 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1469__I _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1747__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1683__A1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2227__A3 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1986__A2 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1738__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1724_ _0476_ _0650_ _0757_ _0794_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1655_ _0719_ _0725_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1586_ _0625_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2163__A2 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2159__B _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2207_ _1187_ _1290_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2138_ _1202_ _1204_ _1208_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1674__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2069_ _0574_ _1138_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1977__A2 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1901__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1665__A1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2090__A1 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1440_ _0505_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2145__A2 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1371_ net37 _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2696__A3 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1656__A1 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1959__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2384__A2 _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2687_ _0469_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1707_ _0783_ _0784_ _0429_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1638_ _0522_ _0524_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1569_ _0643_ _0647_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__1895__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2072__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout54 net55 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout65 net66 net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_6_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2352__B _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1482__I _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1638__A1 _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2610_ _0290_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2366__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2541_ _0154_ _0317_ _0319_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2472_ _0197_ _0199_ _0246_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1423_ _0510_ mapper.bit_Q\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1392__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1354_ net32 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2739_ _0014_ net55 net63 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_59_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2347__B _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2045__A1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2045__B2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2596__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2101__I _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2520__A2 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2257__B _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1972_ _1041_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2587__A2 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2524_ _0299_ _0302_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2455_ _0225_ _0131_ _0227_ _0228_ _0094_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_2386_ _1295_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1406_ _0450_ _0476_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2275__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2578__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2732__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2240_ p_shaping_I.p_shaping_I.bit_in _1319_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2171_ _1191_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2733__RN net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2257__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1955_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1886_ _0909_ _0911_ _0913_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1845__I _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2507_ _0277_ _0281_ _0284_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2438_ _0131_ _0206_ _0208_ _0209_ _1313_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_2369_ _0132_ _0133_ _0025_ _0135_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__2724__RN net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1829__A4 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1740_ _0795_ _0816_ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1671_ _0570_ _0576_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2714__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2223_ _1233_ _0248_ _1235_ _1187_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_38_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2154_ _1247_ _1268_ _1192_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2085_ _1127_ _1142_ _1120_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2650__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1938_ _0816_ _0698_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1869_ _0694_ _0756_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2166__B1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2705__A2 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2641__A1 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1444__A2 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1485__I _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1683__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2265__B _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1723_ _0720_ _0723_ _0800_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1654_ _0729_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1585_ _0664_ _0615_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2206_ _1275_ _1276_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout66_I net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2137_ _1206_ _1202_ _1207_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2068_ _0929_ _0945_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2623__A1 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2139__B1 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1901__A3 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1665__A2 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2085__B _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2614__A1 _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2090__A2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1370_ net36 _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1656__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2605__A1 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output7_I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1592__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2686_ _0471_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1706_ _0582_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1853__I _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1637_ _0714_ _0711_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1568_ _0630_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1499_ _0579_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2684__I _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout55 net62 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout44 p_shaping_Q.p_shaping_I.bit_in net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout66 net67 net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2063__A2 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2540_ _0057_ _0318_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2471_ _0193_ _0196_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1422_ _0507_ gen_sym.Reg_Sym.data_out\[0\] _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1353_ _1236_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1622__B _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2009__I _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2738_ _0002_ _2738_/E _2738_/RN p_shaping_Q.p_shaping_I.ctl_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XANTENNA__1583__I _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1565__A1 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2679__I _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2669_ _0456_ net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2520__A3 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2257__C _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2284__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1971_ _1043_ _1044_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2587__A3 _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1547__A1 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2523_ _0217_ _0300_ _0301_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1617__B _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2454_ _1271_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2385_ _0048_ _0204_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1405_ _0460_ _0468_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput1 ACK net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2275__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1578__I _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2578__A3 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1529__A1 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1701__A1 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2170_ _1160_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1954_ _0976_ _1027_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1768__A1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1885_ _0959_ _0960_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2193__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2506_ _0282_ _0277_ _0283_ _0218_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2437_ _1310_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2368_ _1226_ _0134_ _1246_ _1281_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_56_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2299_ _1243_ _0046_ _0060_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_56_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2641__B _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2420__A2 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2184__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1720__B _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2107__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1670_ _0746_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2175__A1 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2222_ _1201_ _1169_ _1297_ _1299_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2153_ _1221_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2084_ _1127_ _1142_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1989__A1 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2650__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1937_ _0874_ _0965_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2402__A2 _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1868_ _0440_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1799_ _0859_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2166__B2 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2166__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2722__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2687__I _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1591__I _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2469__A2 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2157__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1904__A1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1683__A3 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2745__CLK net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1722_ _0624_ _0617_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1653_ _0573_ _0724_ _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_7_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1584_ _0562_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2300__I _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2205_ _1186_ _1277_ _1280_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2136_ _1173_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_26_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout59_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2067_ _1122_ _1127_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1586__I _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2387__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2139__A1 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1535__B _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1656__A3 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1705_ _0777_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2685_ _1338_ _0470_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1592__A2 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1636_ _0007_ _0661_ _0685_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1567_ _0555_ _0557_ _0644_ _0646_ _0620_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1498_ net43 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2119_ _1187_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout45 net47 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout56 net58 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout67 net68 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2532__A1 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2470_ _0217_ _0235_ _0244_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_1421_ _0509_ p_shaping_I.p_shaping_I.bit_in vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1877__A3 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1352_ net33 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2737_ p_shaping_Q.p_shaping_I.bit_in_1 net59 net48 p_shaping_Q.p_shaping_I.bit_in_2
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2668_ _0445_ _0452_ _0455_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_59_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1619_ _0560_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2599_ _0352_ _0348_ _0382_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2554__B _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1970_ _1002_ _1006_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1795__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2522_ _0235_ _0244_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_5_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2453_ _0056_ _1186_ _1234_ _1204_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2384_ _0048_ _0151_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1404_ net51 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput2 Bit_In net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2464__B _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1859__I _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1710__A2 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2502__A4 _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1718__B _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1529__A2 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1701__A2 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1953_ _0948_ _0877_ _1025_ _1026_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1884_ _0910_ _0922_ _0958_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1768__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2717__A1 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2193__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2505_ _0122_ _0108_ _0278_ _0230_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2436_ _0207_ _1343_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1363__B _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2367_ _1275_ _1168_ _1336_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2298_ _0047_ _0059_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1589__I _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2708__A1 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2369__B _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1998__A2 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1499__I _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2175__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2221_ _1203_ _1298_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2152_ _1215_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2083_ _1147_ _1151_ _1144_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1438__A1 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1936_ _1009_ _0975_ _0981_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2402__A3 _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1867_ _0896_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1610__A1 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1798_ _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1872__I _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2166__A2 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2419_ _0181_ _0187_ _0189_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1677__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2157__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1904__A2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1840__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1957__I _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1721_ _0782_ _0788_ _0798_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_11_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1652_ _0538_ _0602_ _0582_ _0730_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1583_ _0566_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2204_ _1312_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1659__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2135_ _1205_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2066_ _1118_ _1120_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1831__A1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1867__I _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1919_ _0990_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2387__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2139__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1551__B _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2311__A2 _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2382__B _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1813__B2 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1813__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1704_ _0631_ _0780_ _0781_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2684_ _0469_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1635_ _0007_ _0661_ _0685_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1566_ _0557_ _0645_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1497_ _0532_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2118_ _0226_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2049_ _0839_ _0503_ _0633_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_42_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1804__A1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout46 _0004_ net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout68 net4 net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout57 net58 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1546__B _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2296__A1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2048__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1420_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1351_ _1214_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2211__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2736_ p_shaping_I.p_shaping_I.bit_in net60 net46 p_shaping_I.p_shaping_I.bit_in_1
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2667_ _0453_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1618_ _0697_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2598_ _0349_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2514__A2 _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1549_ _0498_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2278__A1 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2450__A1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2745__RN net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2269__A1 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2521_ _0235_ _0244_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1547__A3 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2452_ _1232_ _0224_ _0079_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2383_ _1250_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1403_ net41 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput3 EN net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2719_ _0492_ _0496_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2499__A1 _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2727__RN net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1734__B _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1952_ _0719_ _0502_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2414__A1 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1883_ _0910_ _0922_ _0958_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2504_ _1307_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2435_ _1244_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2366_ _1253_ _1197_ _1299_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_56_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2297_ _0055_ _0058_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2405__A1 _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2708__A2 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1695__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2644__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2220_ _1247_ _1161_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2151_ _1217_ _1219_ _1180_ _1222_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2082_ _1136_ _1137_ _1143_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__2635__A1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1935_ _1008_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1866_ _0940_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1797_ _0814_ _0819_ _0824_ _0520_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__1374__A1 _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2418_ _0109_ _0188_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2349_ _1217_ _1219_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1677__A2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1668__A2 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2617__A1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1720_ _0792_ _0797_ _0759_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1973__I _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1651_ _0564_ _0587_ _0614_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1582_ _0640_ _0661_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2203_ _1278_ _1204_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1659__A2 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2134_ _0054_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2065_ _1135_ net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2608__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1918_ _0751_ _0992_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1849_ _0581_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1551__C _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2311__A3 _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1822__A2 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2066__A2 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1813__A2 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1577__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1703_ _0670_ _0672_ _0779_ _0778_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_8_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2683_ _0467_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1634_ _0640_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1565_ _0591_ _0585_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1652__B _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1496_ _0570_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout64_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1501__A1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2117_ _1185_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2048_ _0503_ _0977_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout47 _0004_ net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout58 net61 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_8_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1740__A1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2296__A2 _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2412__I _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1350_ net35 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2734__D _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2735_ _0013_ net57 net66 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2666_ _0415_ _0441_ _0439_ _0412_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1617_ _0549_ _0666_ _0572_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2597_ _0378_ _0380_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1548_ _0450_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1722__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1479_ _0559_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2269__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2520_ _0265_ _0285_ _0298_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__1952__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2451_ _1252_ _0036_ _1244_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_5_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1402_ net50 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1704__A1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2382_ _0114_ _0148_ _1198_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput4 REQ_SAMPLE net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2680__A2 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2317__I _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2718_ _1084_ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1943__A1 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2649_ _0405_ _0409_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_59_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1934__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1951_ _0876_ _1024_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2414__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1882_ _0934_ _0942_ _0957_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2503_ _0231_ _0279_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2434_ _0205_ _0153_ _1316_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2365_ _1245_ _0131_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2296_ _1295_ _0057_ _1219_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1916__A1 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2644__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2332__A1 _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2150_ _1220_ _1221_ _1216_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_38_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2081_ _1131_ _1134_ _1146_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_19_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1934_ _0609_ _0923_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2399__A1 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1865_ _0894_ _0904_ _0522_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1796_ _0858_ _0871_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2417_ _1297_ _0117_ _1299_ _0050_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2348_ _0110_ _0112_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2279_ _1278_ _1294_ _0037_ _0038_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_25_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2562__A1 _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1650_ _0726_ _0580_ _0727_ _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_7_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1581_ _0642_ _0660_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2202_ _1161_ _0237_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2133_ _0054_ _1279_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2737__D p_shaping_Q.p_shaping_I.bit_in_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2064_ _1131_ _1134_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_19_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1917_ _0953_ _0804_ _0871_ _0991_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_1848_ _0793_ _0603_ _0697_ _0739_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__2544__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1779_ _0577_ _0803_ _0765_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_57_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1702_ _0778_ _0670_ _0672_ _0779_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_2682_ net67 net3 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1577__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1633_ _0639_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1564_ _0548_ _0625_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2526__B2 _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1495_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1501__A2 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2116_ _0096_ _1184_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2047_ _0640_ _1117_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout59 net61 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout48 _0005_ net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1740__A2 _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2296__A3 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2453__B1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1803__I0 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2508__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1753__B _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1472__C _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2734_ _0012_ net57 net65 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2665_ _0435_ _0438_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1616_ _0691_ _0692_ _0693_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2596_ _0335_ _0337_ _0345_ _0379_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1547_ _0552_ _0601_ _0615_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1722__A2 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1478_ net50 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2278__A3 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2513__I _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1573__B _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2505__A4 _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2388__C _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1477__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1799__I _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1401__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1952__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2450_ _0173_ _0222_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2579__B _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1401_ _0408_ _0429_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2381_ _0081_ _0147_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput5 RST net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__2745__D net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2196__A2 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2717_ _1099_ _0493_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1943__A2 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2648_ _0428_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2579_ _0513_ _0360_ _1331_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1459__A1 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1631__A1 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2399__B _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2111__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1870__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1950_ _0944_ _1023_ _0886_ _0885_ _0812_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_1881_ _0530_ _0955_ _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1622__A1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1992__I _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2502_ _0122_ _0108_ _0278_ _0230_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2433_ _1207_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2364_ _0194_ _1276_ _1201_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_56_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2295_ _1174_ _0056_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1613__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1852__A1 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1604__A1 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1745__C _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2580__A2 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2576__C _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2080_ _1149_ net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2148__I _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1933_ _1007_ net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2399__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1864_ _0859_ _0936_ _0938_ _0598_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1795_ _0858_ _0871_ _0531_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2416_ _0182_ _0169_ _0186_ _0079_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2347_ _1168_ _1249_ _0111_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2278_ _1201_ _1336_ _1177_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2087__B2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2562__A2 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2314__A2 _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1825__A1 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1580_ _0649_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2201_ _1275_ _1168_ _1276_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2132_ _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2069__A1 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2063_ _1083_ _1108_ _1133_ _1110_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2606__I _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1916_ _0704_ _0949_ _0950_ _0943_ _0946_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_30_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1847_ _0836_ _0837_ _0833_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1778_ _0855_ net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1420__I _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2232__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1576__B _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2251__I _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2299__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2223__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1701_ _0602_ _0625_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2681_ _0007_ _0466_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1632_ _0662_ _0685_ _0711_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__2526__A2 _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1563_ _0573_ _0397_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1494_ _0571_ _0537_ _0574_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2115_ _1175_ _1192_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2046_ _1114_ _1116_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_54_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout49 _0005_ net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1725__B1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2453__A1 _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2453__B2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2205__A1 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2508__A2 _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2692__A1 _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2156__I _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2733_ _0011_ net59 net67 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2664_ _0428_ _0451_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1615_ _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2595_ _0328_ _0346_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1546_ _0602_ _0625_ _0626_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1477_ _0333_ _0555_ _0557_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_39_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2029_ _1031_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1477__A2 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1400_ _0344_ _0311_ _0418_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2380_ _0089_ _1298_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2417__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2716_ _0492_ _0494_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2647_ _1212_ _0433_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2578_ _0154_ _1164_ _1343_ _0357_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__2353__B1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1529_ _0606_ _0609_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_59_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2647__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1622__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1880_ _0857_ _0954_ _0952_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1925__A3 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2501_ _0167_ _0175_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1494__B _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2432_ _0102_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2363_ _0040_ _1316_ _0127_ _1238_ _0128_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1689__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2294_ _1333_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2638__A1 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2344__I _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1613__A2 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1916__A3 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1852__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output13_I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1368__A1 _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2096__A2 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2635__A4 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1932_ _1002_ _1006_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1863_ _0884_ _0592_ _0644_ _0937_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1794_ _0859_ _0862_ _0867_ _0870_ _0723_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_2415_ _0184_ _0185_ _0078_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2346_ _1162_ _1157_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2277_ _1249_ _0036_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2011__A2 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1522__A1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1825__A2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2200_ _1172_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2131_ _1170_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2062_ _1071_ _1074_ _1132_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1915_ _0948_ _0986_ _0989_ _0944_ _0943_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1846_ _0873_ _0910_ _0908_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1777_ _0772_ _0854_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2329_ _0049_ _0090_ _0091_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2018__B _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2232__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2299__A2 _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2471__A2 _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2223__A2 _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1700_ _0726_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2680_ p_shaping_Q.p_shaping_I.counter\[0\] _1098_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1631_ _0531_ _0710_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1734__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1562_ _0641_ _0606_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1493_ _0572_ _0573_ _0539_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input4_I REQ_SAMPLE vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2114_ _1159_ _1164_ _1171_ _1179_ _1182_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2045_ _0929_ _0946_ _1115_ _1084_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2462__A2 _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1829_ _0607_ _0832_ _0893_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__1725__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2301__B _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1725__B2 _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2150__A1 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2453__A2 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2205__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1606__I p_shaping_Q.p_shaping_I.bit_in_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2692__A2 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2437__I _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2732_ _0010_ net56 net65 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2663_ _0356_ _0449_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1614_ _0663_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2594_ _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1707__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1545_ _0600_ _0322_ _0585_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_59_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2380__A1 _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1476_ _0556_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout62_I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2028_ _1099_ _1014_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1946__A1 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2031__B _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2123__A1 _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output43_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1764__C _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2362__A1 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2114__A1 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2417__A2 _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2715_ _0701_ _0493_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_10_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2646_ _0430_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2577_ _0081_ _0318_ _0358_ _0290_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__2353__A1 _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2353__B2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1528_ _0608_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1459_ _0538_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_67_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1864__B1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1616__B1 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1865__B _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2592__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1386__A2 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2500_ _0219_ _0109_ _0274_ _0276_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2583__B2 _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2431_ _0162_ _0192_ _0201_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2335__A1 _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2362_ _1229_ _1239_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1689__A3 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2293_ _0051_ _0053_ _1182_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2638__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2574__A1 _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1377__A2 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2360__I _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2629_ _0383_ _0384_ _0381_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1595__B _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1368__A2 _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1907__A4 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1614__I _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2445__I _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1931_ _1003_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1862_ _0866_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1793_ _0868_ _0869_ _0631_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2308__A1 _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2414_ _1188_ _1197_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1906__I1 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2345_ _1160_ _1314_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2276_ _1205_ _1231_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1770__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1434__I p_shaping_Q.p_shaping_I.bit_in_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2483__B1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2538__A1 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1513__A2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2130_ _1199_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2061_ _1083_ _1108_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2226__B1 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1914_ _0987_ _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1845_ _0921_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1776_ _0776_ _0807_ _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_2328_ _1207_ _0056_ _1271_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2701__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2259_ _1268_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1440__A1 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1991__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1743__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2299__A3 _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1431__A1 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1982__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1630_ _0687_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1561_ _0520_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1492_ _0450_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2113_ _1180_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2044_ _0937_ _1023_ _0701_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1670__A1 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1422__A1 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1828_ _0895_ _0904_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1759_ _0835_ _0827_ _0828_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1489__A1 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1489__B2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1661__A1 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1652__A1 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2731_ _0009_ net56 net65 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2662_ _0203_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1613_ _0671_ _0676_ _0543_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2593_ _0363_ _0375_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1707__A2 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1544_ _0500_ _0545_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2380__A2 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1475_ _0535_ _0468_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1532__I _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout55_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2027_ _1032_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1643__A1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2123__A2 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2362__A2 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2114__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1352__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1873__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2183__I _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2714_ _0679_ _0467_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2645_ _0041_ _0222_ _0431_ _0390_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1527__I _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2353__A2 _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2576_ _0316_ _0115_ _1245_ _0165_ _0292_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_1527_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1458_ net43 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1864__A1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1389_ net38 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1864__B2 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1616__A1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2592__A2 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1437__I _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2280__A1 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2032__A1 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1347__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2430_ _0178_ _0191_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_51_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1791__B _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2361_ _1343_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2292_ _1267_ _1297_ _0052_ _1278_ _1334_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2178__I _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1846__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1810__I _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2271__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2628_ _0378_ _0380_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2559_ _0182_ _0205_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2262__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1525__B1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1930_ _0960_ _1004_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2253__A1 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1861_ _0755_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1792_ _0783_ _0619_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1764__B1 _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2413_ _0048_ _1252_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2344_ _1345_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2275_ _1226_ _1232_ _1185_ _1253_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_52_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2547__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1715__I _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1522__A3 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1450__I _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2483__A1 _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2483__B2 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2235__A1 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2538__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1625__I _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2060_ _1128_ _1130_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_19_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1360__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2226__B2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2226__A1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1913_ _0860_ _0878_ _0877_ _0984_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2191__I _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1844_ _0916_ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1775_ _0850_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2327_ _0089_ _1245_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2258_ _1335_ _1337_ _1339_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2189_ _1213_ _1261_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2465__A1 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2315__B _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1873__C _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2208__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1431__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1560_ _0608_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1491_ _0554_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2112_ _0107_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2043_ _1021_ _1113_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_47_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1827_ _0896_ _0897_ _0899_ _0903_ _0859_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_1758_ _0835_ _0828_ _0827_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1689_ _0737_ _0749_ _0767_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__2150__A3 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2438__A1 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1661__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1413__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1964__A3 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1652__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2730_ _0008_ net54 net64 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2661_ _0513_ _0446_ _0447_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1612_ _0537_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2592_ _0368_ _0374_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1543_ _0601_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1474_ _0554_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1891__A2 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2026_ _0532_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_fanout48_I _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1643__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2371__A3 _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2659__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1882__A2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1945__I0 p_shaping_Q.p_shaping_I.bit_in_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1570__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1873__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1808__I _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2050__A2 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2713_ _0505_ _0470_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2644_ _0391_ _1228_ _0294_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2575_ _1200_ _0319_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1526_ p_shaping_Q.p_shaping_I.counter\[0\] p_shaping_Q.p_shaping_I.counter\[1\]
+ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1457_ _0365_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1388_ _0291_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1616__A2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2009_ _1081_ net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1552__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1855__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1791__A1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2360_ _0269_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2291_ _1341_ _1235_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2271__A2 _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1538__I _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2627_ _0411_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2558_ _0220_ _1290_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2489_ _0102_ _0264_ _0160_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1509_ _0587_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2262__A2 _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2014__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1525__B2 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1828__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2253__A2 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1860_ _0935_ _0613_ _0865_ _0705_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_14_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1791_ _0664_ _0333_ _0572_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1764__B2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2412_ _1206_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2343_ _0106_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2274_ _1334_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1989_ _0504_ _1061_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2483__A2 _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2235__A2 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1994__A1 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1641__I _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1912_ _0743_ _0645_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1843_ _0918_ _0919_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1737__A1 _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1774_ _0808_ _0851_ _0838_ _0849_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_57_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2326_ _1169_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2257_ _1338_ _1174_ _1178_ _1165_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2188_ _1242_ _1260_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2465__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1976__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2315__C _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1728__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2208__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1719__A1 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1490_ _0355_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1371__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2111_ _1174_ _1177_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2042_ _0830_ _1011_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1826_ _0821_ _0901_ _0902_ _0809_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2151__B _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1757_ _0735_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1688_ _0752_ _0765_ _0766_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2309_ _1327_ _0068_ _0069_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1489__A3 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2374__A1 _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2126__A1 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2287__I _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1652__A3 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2660_ _0314_ _0446_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1611_ _0690_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2591_ _0218_ _0372_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1366__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2365__A1 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1542_ _0613_ _0616_ _0618_ _0619_ _0622_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_4_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1473_ _0460_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input2_I Bit_In vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2197__I _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2025_ _1092_ _1096_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1891__A3 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1809_ _0599_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_2_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2108__A1 _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1882__A3 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2292__B1 _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1570__A2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2586__A1 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2712_ _0490_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2643_ _1331_ _0263_ _0313_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2574_ _0021_ _0103_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1525_ _0580_ _0589_ _0595_ _0598_ _0605_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1456_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1387_ _0280_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout60_I net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2510__A1 _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2008_ _1075_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_23_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2577__A1 _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2329__A1 _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output41_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1909__I _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2514__B _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1791__A2 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2290_ _0049_ _0050_ _1284_ _0025_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_37_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2559__A1 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2626_ _0388_ _0389_ _0410_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2557_ _0335_ _0337_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2488_ _0261_ _0263_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1508_ _0581_ _0582_ _0584_ _0588_ _0533_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1439_ _0514_ _0523_ _0524_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1503__B _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1464__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1790_ _0694_ _0864_ _0865_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__1764__A2 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2411_ _0094_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2342_ _1257_ _1305_ _0044_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2713__A1 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1516__A2 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2273_ _1329_ _0031_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2154__B _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1988_ _0839_ _1060_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2609_ _0321_ _0209_ _0091_ _0392_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1507__A2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2329__B _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2235__A3 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1994__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1911_ _0883_ _0985_ _0691_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_15_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1842_ _0772_ _0854_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1737__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1773_ _0831_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2325_ _0075_ _0029_ _0086_ _0087_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2256_ _1167_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2187_ _1262_ net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1898__B _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2573__I _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2519__I1 p_shaping_I.p_shaping_I.bit_in vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2110_ _0096_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2041_ _1112_ net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1655__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1407__A1 _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1825_ _0720_ _0593_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1756_ _0833_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2151__C _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1687_ _0752_ _0765_ p_shaping_Q.p_shaping_I.counter\[1\] _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1894__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2308_ _0021_ _0031_ _0061_ _0063_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2239_ _1215_ _1223_ _1230_ _1240_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1646__A1 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2374__A2 _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1647__I _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1610_ _0566_ _0548_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2590_ _1307_ _0371_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2365__A2 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1541_ _0620_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1472_ _0547_ _0549_ _0550_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_67_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2024_ _0839_ _1094_ _1095_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1628__A1 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1557__I _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1808_ _0884_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1739_ _0549_ _0537_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2292__B2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2292__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2044__A1 _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1467__I _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2347__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1858__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2283__A1 _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2035__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2711_ _0885_ _0487_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2642_ _0426_ _0427_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2573_ _0354_ net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1524_ _0599_ _0603_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1455_ _0535_ _0311_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_67_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1386_ _0183_ _0269_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2510__A2 _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2007_ _1077_ _1079_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2157__B _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1552__A3 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2741__RN net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2265__A1 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2017__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2731__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2491__I _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2559__A2 _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2625_ _0388_ _0389_ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2556_ _0282_ _0283_ _0336_ _1292_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2487_ _0157_ _0262_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1507_ _0585_ _0586_ _0587_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1438_ net59 p_shaping_Q.p_shaping_I.ctl_1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1369_ _1214_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2486__A1 _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2238__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2410__A1 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2410_ _0508_ _0179_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2341_ _1329_ _0103_ _0104_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_35_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2713__A2 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1921__B1 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2272_ _1331_ _0027_ _0030_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2229__A1 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1987_ _0985_ _0553_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2401__A1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2608_ _0391_ _0340_ _0224_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2539_ _0254_ _1159_ _0268_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2396__I _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1514__B _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2255__B _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1910_ _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1841_ _0776_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1772_ _0808_ _0832_ _0838_ _0849_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__1737__A3 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2324_ p_shaping_I.p_shaping_I.bit_in_1 _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2255_ _0194_ _1336_ _1218_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2186_ _1213_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_65_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1673__A2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2689__A1 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1664__A2 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2613__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1933__I _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2040_ _1083_ _1108_ _1111_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_35_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1655__A2 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2604__A1 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1407__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1824_ _0886_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1755_ _0718_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1686_ _0753_ _0754_ _0760_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_38_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2307_ _1329_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2238_ _1345_ _1311_ _1315_ _1317_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__1894__A2 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2169_ p_shaping_I.p_shaping_I.counter\[1\] _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1582__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1540_ _0564_ _0614_ _0587_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1471_ _0551_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2708__B _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2023_ _0977_ _1094_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1807_ _0789_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1738_ _0543_ _0706_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2669__I _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1669_ net44 _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2292__A2 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2263__B _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2710_ _0489_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1794__A1 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1794__B2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2641_ _0420_ _0422_ _0424_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1546__A1 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2572_ _0350_ _0353_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1393__I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1523_ _0583_ _0567_ _0538_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1454_ net39 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1385_ _0204_ _0258_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2006_ _1043_ _1040_ _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout46_I _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2173__B _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1785__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2265__A2 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1478__I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2102__I _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1700__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1388__I _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1767__A1 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2624_ _0400_ _0405_ _0409_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__2012__I _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2555_ _0334_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2486_ _0087_ _0213_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1506_ _0355_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1437_ _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1368_ _0043_ _0074_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1761__I p_shaping_Q.p_shaping_I.bit_in vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2486__A2 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1749__A1 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2340_ _0101_ _0088_ _0100_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__1921__B2 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2271_ _0511_ _0029_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1988__A1 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1986_ _0756_ _0877_ _0695_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2401__A2 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2451__B _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2607_ _0316_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2538_ _0316_ _1266_ _0184_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1912__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2469_ _0236_ _0243_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_24_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1667__B1 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1840_ _0807_ _0853_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_30_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2395__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1771_ _0840_ _0848_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2147__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2323_ _0077_ _0084_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2254_ _1172_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2185_ _1242_ _1260_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_25_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1969_ _1042_ _1001_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2181__B _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2744__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2689__A2 _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2310__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1486__I _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2129__A1 _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2110__I _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2604__A2 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1812__B1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1823_ _0690_ _0868_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2368__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1754_ _0831_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1685_ _0693_ _0681_ _0762_ _0763_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_2306_ _1329_ _0031_ _0061_ _0063_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__2540__A1 _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2237_ _1195_ _1284_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_26_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2168_ _1224_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2176__B _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2099_ _1258_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2359__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2531__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1573__A2 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1470_ _0535_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2522__A1 _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2022_ _1026_ _0633_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1806_ _0809_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1564__A2 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1737_ _0606_ _0649_ _0659_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1668_ _0635_ _0683_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_49_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1599_ _0678_ _0626_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2618__C _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2353__C _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2544__B _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2640_ _0425_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2571_ _0304_ _0303_ _0305_ _0352_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1546__A2 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1522_ _0600_ _0601_ _0602_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_4_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1453_ _0533_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1384_ _0215_ _0237_ _0248_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_67_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2438__C _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2510__A4 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2005_ _1039_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2173__C _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1785__A2 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1584__I _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1537__A2 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2364__B _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1776__A2 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2623_ _0516_ _0406_ _0407_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2554_ _0232_ _0279_ _0334_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1505_ _0344_ _0311_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2485_ _0250_ _0257_ _0259_ _0260_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1436_ net44 _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1367_ _0054_ _1170_ _1279_ _0065_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_55_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2707__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1694__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1749__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2113__I _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2270_ _1200_ _1209_ _1274_ _1286_ _0028_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__1901__B _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1685__A1 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1985_ _1008_ _1057_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2606_ _0290_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2537_ _0268_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1912__A2 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2468_ _0239_ _0241_ _0242_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_57_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1419_ gen_sym.Reg_Sym.data_out\[1\] _0507_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2399_ _1165_ _1252_ _1188_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1811__B _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1979__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1903__A2 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1667__B2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1667__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1770_ _0841_ _0842_ _0844_ _0847_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__2395__A2 _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2322_ _0034_ _0080_ _0083_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2253_ _1169_ _1333_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2184_ _1243_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1658__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2462__B _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1968_ _0997_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1899_ _0875_ _0965_ _0972_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2138__A2 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2689__A3 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1897__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1649__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1821__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2129__A2 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2301__A2 _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1812__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1822_ _0898_ _0743_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2368__A2 _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1753_ _0826_ _0829_ _0830_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1684_ _0624_ _0645_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2305_ _0067_ net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2236_ _1205_ _1233_ _1187_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_53_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2167_ _1230_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2098_ _0215_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1567__B1 _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2531__A2 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2047__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2522__A2 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2021_ _1084_ _0944_ _0691_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2734__CLK net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2589__A2 _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1805_ _0860_ _0603_ _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1736_ _0612_ _0813_ _0729_ _0732_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_1667_ _0728_ _0738_ _0740_ _0705_ _0745_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_1598_ _0566_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2277__A1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2219_ _1205_ _1167_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1960__B1 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2744__RN net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2268__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2544__C _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2440__A1 _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2560__B _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2570_ _0351_ _0302_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1521_ _0541_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1452_ net50 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1703__B1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1383_ _0140_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_67_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2004_ _1003_ _1005_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2026__I _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1719_ _0692_ _0796_ _0665_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2699_ _0480_ _0481_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1814__B _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2726__RN net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1536__I0 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2661__A1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2413__A1 _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2290__B _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2622_ _0289_ _0406_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2553_ _0330_ _0332_ _0250_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1504_ _0418_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2484_ _0220_ _0150_ _0052_ _0109_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1435_ _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1366_ net36 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout51_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2404__A1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1915__B1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2643__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1685__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2634__A1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1984_ _0834_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2605_ _0363_ _0375_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2536_ _0115_ _0165_ _0185_ _0111_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2467_ _0041_ _0151_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1418_ net1 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2179__C _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2398_ _1313_ _0166_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_28_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1676__A2 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1349_ _1170_ _1192_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_24_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1600__A2 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2616__A1 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1419__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2321_ _1222_ _0081_ _0082_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_2_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2252_ _1236_ _1258_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_65_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2183_ _1257_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1967_ _1039_ _1040_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1594__A1 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1898_ _0875_ _0965_ _0972_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2519_ _0289_ p_shaping_I.p_shaping_I.bit_in _0297_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1821__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1585__A1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1783__I _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1812__A2 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1821_ _0676_ _0543_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2282__C _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1752_ _0506_ _0717_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1683_ _0761_ _0726_ _0476_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2304_ _1324_ _0066_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2235_ _1255_ _1313_ _1314_ _0161_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2166_ _1232_ _1234_ _1237_ _1238_ _1239_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_53_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2097_ _1160_ _1163_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__1868__I _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1567__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2295__A2 _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1778__I _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2020_ _1009_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2293__B _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1797__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1804_ _0761_ _0860_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1735_ _0809_ _0810_ _0811_ _0571_ _0812_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_1666_ _0741_ _0744_ _0658_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1597_ _0671_ _0676_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2218_ _1255_ _1159_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2149_ _1214_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1598__I _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1788__A1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1960__B2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1712__A1 _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2132__I _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1951__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1520_ _0408_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1451_ _0531_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1382_ _0226_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1703__B2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2288__B _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2003_ _1002_ _1041_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1367__B _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1718_ _0793_ _0794_ _0795_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2698_ _0270_ _0474_ _0292_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1942__A1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1649_ _0620_ _0630_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_58_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2198__B _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2498__A2 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2217__I _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2186__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1536__I1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2413__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2290__C _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2621_ _0146_ _1203_ _0219_ _0172_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2552_ _0267_ _0184_ _0050_ _0331_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1503_ _0583_ _0322_ _0542_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2483_ _0204_ _0115_ _1283_ _1284_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1434_ p_shaping_Q.p_shaping_I.bit_in_1 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1365_ _1236_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1650__B _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout44_I p_shaping_Q.p_shaping_I.bit_in vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2404__A2 _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2707__A3 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2340__A1 _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1786__I _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2159__A1 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1983_ _0521_ _1054_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2398__A1 _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1696__I _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2604_ _0368_ _0374_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2535_ _0263_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2466_ _1344_ _0154_ _0240_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1417_ _0506_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2322__A1 _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2397_ _0164_ _0052_ _0082_ _0165_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1348_ _1181_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1675__I0 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2552__A1 _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2320_ _1335_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2251_ _1195_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2304__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2182_ _1244_ _1245_ _1248_ _1254_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_18_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1966_ _1010_ _0995_ _1038_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_21_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1897_ _0876_ _0968_ _0970_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1594__A2 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2518_ _0290_ _0293_ _0294_ _0173_ _0296_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__2543__A1 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2449_ _0219_ _0221_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_56_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1585__A2 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2534__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1820_ _0756_ _0817_ _0884_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2135__I _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1576__A2 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1751_ _0735_ _0827_ _0828_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1682_ _0583_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2303_ _1327_ _0033_ _0064_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2234_ _1167_ _1172_ _0215_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2165_ _0118_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1500__A2 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2096_ _1161_ _1162_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1949_ _0878_ _0898_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2516__A1 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2507__A1 _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1743__B _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1494__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1797__A2 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1803_ _0688_ _0879_ _0700_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1734_ _0652_ _0590_ _0501_ _0629_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_1665_ _0721_ _0742_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1596_ _0652_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2217_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_38_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2148_ _0129_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2484__B _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2079_ _1146_ _1148_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1788__A2 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1960__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2659__B _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1789__I _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1450_ _0530_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1381_ net35 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2002_ _1071_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2697_ _0391_ _0321_ _0477_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1717_ _0590_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1942__A2 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1648_ _0554_ _0556_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1579_ _0654_ _0656_ _0657_ _0603_ _0658_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1402__I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2389__B _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2620_ _0232_ _0403_ _0404_ _0062_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__2143__I _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2551_ _0207_ _0272_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2482_ _0251_ _0091_ _0256_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1502_ _0551_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1433_ _0513_ net45 _0519_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1364_ net37 _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2519__S _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1860__A1 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2707__A4 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1851__A1 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1735__C _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2634__A3 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1982_ _1011_ _1054_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2603_ _0386_ net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2534_ _1331_ _0312_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2465_ _1186_ _1277_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2396_ _1337_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1416_ _0505_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2322__A2 _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1347_ net34 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1661__B _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2561__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1824__A1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1675__I1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1746__B _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2250_ _0280_ _1330_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2181_ _1255_ _1253_ _1239_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2737__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2068__A1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1965_ _1010_ _0995_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2240__A1 p_shaping_I.p_shaping_I.bit_in vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1896_ _0935_ _0816_ _0929_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2331__I _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2517_ _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2448_ _0220_ _1228_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2379_ _0034_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1410__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2231__A1 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2222__A1 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1750_ _0641_ _0814_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1681_ _0619_ _0755_ _0756_ _0757_ _0759_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2302_ _0061_ _0063_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_2_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2233_ _1312_ _1323_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2164_ _0096_ _1176_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_26_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2095_ _0140_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2326__I _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2213__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1948_ _0834_ _1019_ _1021_ _0640_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1879_ _0751_ _0952_ _0954_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2452__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1494__A2 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2443__A1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1797__A3 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1802_ _0694_ _0785_ _0877_ _0878_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1733_ _0615_ _0666_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1664_ _0563_ _0565_ _0538_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1595_ _0670_ _0672_ _0534_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1721__A3 _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2216_ _0107_ _0118_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_fanout67_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2147_ _1173_ _1176_ _1218_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2682__A1 net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2078_ _1131_ _1134_ _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2434__A1 _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1960__A3 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1779__A3 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1380_ _0129_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2001_ _1072_ _1037_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_35_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2416__A1 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2696_ _0183_ _0269_ _0469_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1664__B _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1716_ _0669_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1647_ _0565_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1578_ _0579_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_58_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1630__A2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1697__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2550_ _0329_ _0294_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1385__A1 _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2481_ _0252_ _0040_ _0253_ _0255_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1501_ _0500_ net38 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1432_ _0291_ _0518_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1363_ _1203_ _1301_ _1345_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1688__A2 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2637__A1 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2739__SETN net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1860__A2 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1376__A1 _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2679_ _0465_ net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1679__A2 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1981_ _1049_ _1052_ _1053_ _0719_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_60_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2602_ _0381_ _0385_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2533_ _0075_ _0030_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1358__A1 _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2103__B _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2464_ _0151_ _0238_ _1200_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2395_ _1267_ _0150_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1415_ _0333_ _0397_ _0504_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1346_ net35 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1597__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2010__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2013__B _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1408__I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1852__B _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2077__A2 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1588__A1 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2001__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2552__A3 _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1762__B _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1760__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2577__C _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2180_ _1170_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1964_ _1022_ _1029_ _1037_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__1579__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1579__B2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1895_ _0863_ _0674_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2516_ _0131_ _0206_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2447_ _1225_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2378_ _0145_ net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2231__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1990__A1 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1742__A1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1601__I _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2470__A2 _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2222__A2 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1680_ _0758_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1981__B2 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2301_ _0062_ _0046_ _0060_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1733__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2232_ _1310_ _1302_ _1303_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2289__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2163_ _1233_ _1216_ _1235_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2607__I _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2094_ _1258_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1947_ _0718_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1878_ _0953_ _0804_ _0871_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1724__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1724__B2 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2452__A2 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1577__B _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2727__CLK net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2443__A2 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1801_ _0673_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1487__B _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1732_ _0621_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1663_ _0557_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1594_ _0572_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2111__B _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2215_ p_shaping_I.p_shaping_I.bit_in_2 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2146_ _0226_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2682__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2077_ _1128_ _1130_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1416__I _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2370__A1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2122__A1 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2247__I _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2425__A2 _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2189__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1400__A3 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2000_ _1022_ _1029_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2416__A2 _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1715_ _0565_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2695_ _0478_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1646_ _0720_ _0722_ _0723_ _0724_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1577_ _0555_ _0626_ _0561_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_58_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2352__A1 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2129_ _0043_ _1198_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2646__A2 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1385__A2 _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2582__A1 _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2480_ _0254_ _0252_ _0253_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1500_ _0554_ _0556_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1431_ _0514_ _0516_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1362_ _1312_ _1334_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2747_ _0021_ net60 net46 p_shaping_I.p_shaping_I.counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2678_ _1322_ _0464_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1376__A2 _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2350__I _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1629_ _0689_ _0696_ _0702_ _0708_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1851__A3 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2316__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1980_ _0984_ _0688_ _0816_ _0698_ _1051_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_60_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2435__I _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2601_ _0383_ _0384_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2532_ _0265_ _0308_ _0309_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1358__A2 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2170__I _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2463_ _0205_ _1159_ _0117_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2394_ _0122_ _0108_ _1293_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1414_ _0491_ _0499_ _0503_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_24_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1597__A2 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1349__A2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1588__A2 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1815__A3 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1963_ _1030_ _1035_ _1036_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1894_ _0863_ _0604_ _0896_ _0626_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2515_ _0228_ _1203_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2446_ _1301_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2377_ _0071_ _0144_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2700__A1 _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1990__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1863__B _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1742__A2 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2470__A3 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2222__A3 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2300_ _1243_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2231_ _1225_ _1227_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2162_ _1189_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1497__A1 _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2093_ _0226_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1948__B _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1667__C _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1946_ _0734_ _0735_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1877_ _0782_ _0788_ _0798_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1724__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2429_ _0200_ net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1488__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1412__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1612__I _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1768__B _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1800_ _0817_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1731_ _0563_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1662_ _0671_ _0547_ _0678_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1593_ _0501_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1950__C _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2214_ p_shaping_I.p_shaping_I.counter\[1\] _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2145_ _1216_ _1158_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2076_ _1144_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1678__B _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1929_ _0962_ _0959_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2370__A2 _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1860__C _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1881__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1633__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1714_ _0790_ _0791_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2694_ _0391_ _0477_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1645_ _0664_ _0621_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1576_ _0655_ _0584_ _0629_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1863__A1 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2128_ _0237_ _1197_ _0065_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2059_ _1009_ _1091_ _1096_ _1129_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1427__I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1854__A1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2031__A1 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2582__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1430_ p_shaping_I.p_shaping_I.ctl_1 _0514_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1781__B _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1361_ _1323_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1542__B1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2270__A1 _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2746_ _0020_ net60 net46 p_shaping_I.p_shaping_I.counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2677_ _1263_ _1264_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1628_ _0704_ _0707_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2325__A2 _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1559_ _0578_ _0636_ _0638_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1836__A1 _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2013__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1367__A3 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2316__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1827__A1 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1827__B2 _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1620__I _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2600_ _0304_ _0303_ _0305_ _0350_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_2531_ _0285_ _0298_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2462_ _0179_ _0190_ _0516_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2393_ _0102_ _0159_ _0160_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1413_ _0498_ _0502_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1818__A1 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2361__I _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2546__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2729_ _0000_ _2729_/E _2729_/RN p_shaping_I.p_shaping_I.ctl_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
XFILLER_3_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2234__A1 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1588__A3 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1745__B1 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1615__I _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1350__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1962_ _0857_ _0992_ _1035_ _0530_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2225__A1 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1893_ _0966_ _0967_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2114__C _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2514_ _0164_ _0082_ _0292_ _0168_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2445_ _1292_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2376_ _0073_ _0143_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_56_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2356__I _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2464__A1 _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1863__C _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1742__A3 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2266__I _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2455__B2 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1430__A2 _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2230_ _1292_ _1306_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2161_ _1233_ _1216_ _1160_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2694__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2092_ _1158_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1948__C _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1945_ p_shaping_Q.p_shaping_I.bit_in_1 _1011_ _1018_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1876_ _0947_ _0951_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2428_ _0197_ _0199_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2359_ _1292_ _0123_ _0124_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__2685__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1488__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2019__C _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1412__A2 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1730_ _0607_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1661_ _0739_ _0599_ _0644_ _0658_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_1592_ _0671_ _0652_ _0550_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2213_ _1211_ _1289_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2144_ _1192_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2075_ _1136_ _1137_ _1143_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__1890__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1928_ _0918_ _0919_ _0916_ _0961_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1859_ _0739_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1936__A3 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2649__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2454__I _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1713_ _0653_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2693_ _1290_ _0467_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1644_ _0678_ _0669_ _0706_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1575_ _0546_ _0614_ _0408_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1533__I _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1863__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2127_ _0054_ _1175_ _0140_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2058_ _1098_ _1097_ _1105_ _1106_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_54_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2576__B1 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2040__A2 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1551__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1790__A1 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1360_ net37 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1542__B2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1542__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2022__A2 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2745_ net44 net59 net49 p_shaping_Q.p_shaping_I.bit_in_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2676_ _0458_ _0462_ _0463_ net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1781__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1627_ _0624_ _0705_ _0706_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1558_ _0611_ _0635_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1489_ _0534_ _0544_ _0553_ _0558_ _0569_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2261__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2013__A2 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1524__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2530_ _0285_ _0298_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1763__A1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2461_ _0218_ _0234_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1412_ _0460_ net50 _0501_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2392_ _1328_ _0103_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1515__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1818__A2 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2128__B _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2728_ p_shaping_I.p_shaping_I.bit_in_1 net60 net46 p_shaping_I.p_shaping_I.bit_in_2
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2659_ _1332_ _0221_ _1256_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2089__I _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2482__A2 _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1745__B2 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1681__B1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1961_ _1031_ _1034_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1892_ _0866_ _0693_ _0817_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1984__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2513_ _1182_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1806__I _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2444_ _0203_ _0216_ _0160_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2375_ _0105_ _0142_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_29_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2161__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1716__I _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1451__I _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2455__A2 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2207__A2 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1626__I _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2160_ _1166_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2457__I _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2091_ _1157_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1944_ _0759_ _1013_ _1015_ _0787_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1875_ _0948_ _0949_ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1709__A1 _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2382__A1 _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2427_ _0071_ _0144_ _0198_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2509__I0 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2358_ p_shaping_I.p_shaping_I.bit_in_2 _0121_ _0106_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2685__A2 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2289_ _1336_ _1177_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1948__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1874__C _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1446__I _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2373__A1 _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2428__A2 _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1939__A1 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1660_ _0655_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_7_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1591_ _0600_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2116__A1 _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2212_ _1287_ _1288_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2143_ _0085_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2074_ _1136_ _1137_ _1143_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2419__A2 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1975__B _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1927_ _0997_ _1001_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1858_ _0609_ _0923_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1789_ _0573_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2355__A1 _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2740__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2346__A1 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2649__A2 _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2282__B1 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1795__B _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1712_ _0552_ _0777_ _0789_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2692_ _0050_ _0472_ _0475_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1643_ _0721_ _0397_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2337__A1 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1574_ _0651_ _0653_ _0550_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2126_ _1186_ _1193_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout58_I net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2057_ _1122_ _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2576__A1 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1551__A2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2500__A1 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output39_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2555__I _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2319__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1790__A2 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1634__I _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1809__I _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2744_ _0019_ net53 net64 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2675_ _0459_ _0461_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1626_ _0582_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1557_ _0637_ net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1488_ _0561_ _0568_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2109_ _1176_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2549__A1 _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2721__A1 _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1454__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1524__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2485__B1 _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2234__B _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2460_ _0230_ _0233_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1763__A2 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1411_ _0500_ net51 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_47_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1364__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2391_ _0156_ _0158_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_24_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2727_ mapper.bit_Q\[1\] net53 net48 p_shaping_Q.p_shaping_I.bit_in vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2658_ _0444_ _0434_ _0426_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1609_ _0534_ _0688_ _0648_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2589_ _0282_ _0149_ _0281_ _0371_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2703__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2319__B _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1442__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1449__I p_shaping_Q.p_shaping_I.counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1993__A2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1745__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2229__B _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1681__A1 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1960_ _1032_ _0476_ _0731_ _0869_ _1014_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
X_1891_ _0793_ _0795_ _0794_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__1359__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1433__A1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2512_ _0181_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1736__A2 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2443_ _0513_ _0213_ _0214_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2374_ _0125_ _0141_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2161__A2 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1732__I _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2049__B _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1415__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1718__A2 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2090_ net33 net32 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_48_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1943_ _0704_ _0812_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_14_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1874_ _0925_ _0784_ _0594_ _0878_ _0700_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__1709__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2426_ _0073_ _0143_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2357_ _1293_ _0108_ _0122_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1893__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2288_ _0048_ _1184_ _1218_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1645__A1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2070__A1 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1462__I _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1939__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1590_ _0664_ _0669_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2211_ _0511_ _1210_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1372__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2142_ _1210_ _1212_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2073_ _1120_ _1126_ _1142_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1627__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2052__A1 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1926_ _0999_ _0957_ _1000_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1857_ _0830_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1788_ _0795_ _0742_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2409_ _0137_ _0138_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1866__A1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2291__A1 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2043__A1 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1857__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1609__A1 _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2282__A1 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2282__B2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1711_ _0601_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2691_ _0254_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1642_ _0322_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1573_ _0563_ _0652_ _0542_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1848__B2 _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2125_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1830__I _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2056_ _1126_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2147__B _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1909_ _0720_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2576__A2 _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2328__A2 _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2500__A2 _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2740__RN net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2264__A1 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2558__A2 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2743_ _0018_ net52 net64 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
XFILLER_8_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2674_ _0445_ _0452_ _0459_ _0461_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1625_ _0620_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1556_ _0578_ _0636_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1487_ _0563_ _0565_ _0566_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2656__I _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2108_ _0129_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_54_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2039_ _1109_ _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2730__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1524__A3 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2485__A1 _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2237__A1 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1410_ net39 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2390_ _0030_ _0157_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2476__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1380__I _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2400__A1 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2726_ gen_sym.Reg_2M.data_in net52 gen_sym.Reg_2M.enable gen_sym.Reg_2M.data_out
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2657_ _0426_ _0427_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1608_ _0596_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2588_ _0242_ _0369_ _0370_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2703__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1539_ _0559_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2467__A1 _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2386__I _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2219__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1442__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1414__B _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1890_ _0927_ _0928_ _0930_ _0641_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2511_ _0515_ _0288_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2442_ _0157_ _0213_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2373_ _0137_ _0139_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2697__A1 _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2449__A1 _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2709_ _0487_ _0488_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2612__A1 _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1415__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1942_ _0761_ _0935_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1406__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1873_ _0613_ _0588_ _0866_ _0935_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__1709__A3 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1590__A1 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2425_ _0193_ _0196_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2356_ _0121_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2287_ _1220_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1645__A2 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2061__A2 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2210_ _1274_ _1286_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2141_ _1211_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2072_ _0830_ _1141_ _1009_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_53_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1602__B _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2417__C _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1627__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1925_ _0998_ _0933_ _0942_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2052__A2 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1856_ _0521_ _0874_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1787_ _0761_ _0863_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__1563__A1 _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2408_ _0163_ _0176_ _0177_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2339_ _0088_ _0100_ _0102_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2608__B _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1473__I _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1609__A2 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2282__A2 _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1710_ _0786_ _0787_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2690_ _0266_ _0204_ net65 net3 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__1793__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1641_ _0629_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2479__I _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1572_ _0546_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1545__A1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I RST vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1848__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2124_ _0107_ _1323_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2055_ _1098_ _1124_ _1125_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1908_ _0808_ _0832_ _0975_ _0981_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1839_ _0914_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2016__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput40 net40 addQ[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_36_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2742_ _0017_ net55 net63 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffsnq_1
X_2673_ _0427_ _0451_ _0425_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1624_ _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1555_ _0611_ _0635_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1486_ _0418_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout63_I net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2494__A2 _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2107_ net32 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2038_ _1077_ _1079_ _1075_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2621__B _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1772__A4 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2182__A1 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2237__A2 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1748__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2173__A1 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1920__A1 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2476__A2 _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2492__I _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1739__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2725_ gen_sym.Reg_2M.data_out net53 net45 gen_sym.Reg_Sym.data_out\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2656_ _0443_ net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1607_ _0686_ _0577_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2164__A1 _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2587_ _0146_ _0224_ _0091_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1911__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1538_ _0586_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1469_ _0408_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2467__A2 _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2219__A2 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1978__A1 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1481__I _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2510_ _0137_ _0138_ _0287_ _0243_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_5_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2441_ _0210_ _0211_ _0212_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2372_ _0509_ _0138_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2697__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2621__A2 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2385__A1 _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2708_ _0619_ _0470_ _0887_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2137__A1 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2639_ _0420_ _0422_ _0424_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_58_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2688__A2 _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1415__A3 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1476__I _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2743__CLK net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1941_ _0811_ _1014_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1872_ _0704_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1590__A2 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2424_ _0125_ _0141_ _0195_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2355_ _0109_ _0113_ _0116_ _0120_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2286_ _1319_ _1318_ p_shaping_I.p_shaping_I.bit_in _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1802__B1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2530__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1636__A3 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2521__A1 _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1875__A3 _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ p_shaping_I.p_shaping_I.counter\[1\] p_shaping_I.p_shaping_I.counter\[0\]
+ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2071_ _1011_ _1139_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1602__C _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1627__A3 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1924_ _0998_ _0933_ _0942_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1855_ _0927_ _0928_ _0930_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1786_ _0547_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1563__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2407_ _0163_ _0176_ _1243_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2338_ _0101_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2269_ _1183_ _1196_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_55_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2579__A1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1793__A2 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1640_ _0648_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1571_ _0567_ _0650_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1613__B _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2123_ _1188_ _1190_ _1191_ _1334_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2495__I _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2054_ _1065_ _1101_ _1123_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__1856__I0 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1907_ _0808_ _0832_ _0975_ _0981_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__1784__A2 _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1838_ _0909_ _0911_ _0913_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1769_ _0845_ _0846_ _0658_ _0722_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_66_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1523__B _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1472__A1 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2264__A3 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput6 net6 I[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput30 net30 Q[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput41 net41 addQ[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_48_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1463__A1 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2741_ _0016_ net55 net63 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__1766__A2 _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2672_ _1212_ _0430_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2715__A1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1623_ _0580_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1554_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1485_ _0460_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

