magic
tech gf180mcuC
magscale 1 5
timestamp 1670198986
<< obsm1 >>
rect 672 1538 29288 28321
<< metal2 >>
rect 672 29600 728 29900
rect 3360 29600 3416 29900
rect 6048 29600 6104 29900
rect 9072 29600 9128 29900
rect 11760 29600 11816 29900
rect 14448 29600 14504 29900
rect 17472 29600 17528 29900
rect 20160 29600 20216 29900
rect 23184 29600 23240 29900
rect 25872 29600 25928 29900
rect 28560 29600 28616 29900
rect 0 100 56 400
rect 2688 100 2744 400
rect 5376 100 5432 400
rect 8400 100 8456 400
rect 11088 100 11144 400
rect 13776 100 13832 400
rect 16800 100 16856 400
rect 19488 100 19544 400
rect 22176 100 22232 400
rect 25200 100 25256 400
rect 27888 100 27944 400
<< obsm2 >>
rect 14 29570 642 29600
rect 758 29570 3330 29600
rect 3446 29570 6018 29600
rect 6134 29570 9042 29600
rect 9158 29570 11730 29600
rect 11846 29570 14418 29600
rect 14534 29570 17442 29600
rect 17558 29570 20130 29600
rect 20246 29570 23154 29600
rect 23270 29570 25842 29600
rect 25958 29570 28530 29600
rect 28646 29570 29722 29600
rect 14 430 29722 29570
rect 86 400 2658 430
rect 2774 400 5346 430
rect 5462 400 8370 430
rect 8486 400 11058 430
rect 11174 400 13746 430
rect 13862 400 16770 430
rect 16886 400 19458 430
rect 19574 400 22146 430
rect 22262 400 25170 430
rect 25286 400 27858 430
rect 27974 400 29722 430
<< metal3 >>
rect 29600 28560 29900 28616
rect 100 27888 400 27944
rect 29600 25872 29900 25928
rect 100 25200 400 25256
rect 29600 23184 29900 23240
rect 100 22176 400 22232
rect 29600 20160 29900 20216
rect 100 19488 400 19544
rect 29600 17472 29900 17528
rect 100 16800 400 16856
rect 29600 14448 29900 14504
rect 100 13776 400 13832
rect 29600 11760 29900 11816
rect 100 11088 400 11144
rect 29600 9072 29900 9128
rect 100 8400 400 8456
rect 29600 6048 29900 6104
rect 100 5376 400 5432
rect 29600 3360 29900 3416
rect 100 2688 400 2744
rect 29600 672 29900 728
<< obsm3 >>
rect 9 28646 29727 29274
rect 9 28530 29570 28646
rect 9 27974 29727 28530
rect 9 27858 70 27974
rect 430 27858 29727 27974
rect 9 25958 29727 27858
rect 9 25842 29570 25958
rect 9 25286 29727 25842
rect 9 25170 70 25286
rect 430 25170 29727 25286
rect 9 23270 29727 25170
rect 9 23154 29570 23270
rect 9 22262 29727 23154
rect 9 22146 70 22262
rect 430 22146 29727 22262
rect 9 20246 29727 22146
rect 9 20130 29570 20246
rect 9 19574 29727 20130
rect 9 19458 70 19574
rect 430 19458 29727 19574
rect 9 17558 29727 19458
rect 9 17442 29570 17558
rect 9 16886 29727 17442
rect 9 16770 70 16886
rect 430 16770 29727 16886
rect 9 14534 29727 16770
rect 9 14418 29570 14534
rect 9 13862 29727 14418
rect 9 13746 70 13862
rect 430 13746 29727 13862
rect 9 11846 29727 13746
rect 9 11730 29570 11846
rect 9 11174 29727 11730
rect 9 11058 70 11174
rect 430 11058 29727 11174
rect 9 9158 29727 11058
rect 9 9042 29570 9158
rect 9 8486 29727 9042
rect 9 8370 70 8486
rect 430 8370 29727 8486
rect 9 6134 29727 8370
rect 9 6018 29570 6134
rect 9 5462 29727 6018
rect 9 5346 70 5462
rect 430 5346 29727 5462
rect 9 3446 29727 5346
rect 9 3330 29570 3446
rect 9 2774 29727 3330
rect 9 2658 70 2774
rect 430 2658 29727 2774
rect 9 758 29727 2658
rect 9 686 29570 758
<< metal4 >>
rect 2224 1538 2384 28254
rect 9904 1538 10064 28254
rect 17584 1538 17744 28254
rect 25264 1538 25424 28254
<< obsm4 >>
rect 1078 28284 28602 29279
rect 1078 1508 2194 28284
rect 2414 1508 9874 28284
rect 10094 1508 17554 28284
rect 17774 1508 25234 28284
rect 25454 1508 28602 28284
rect 1078 737 28602 1508
<< labels >>
rlabel metal2 s 14448 29600 14504 29900 6 ACK
port 1 nsew signal input
rlabel metal2 s 672 29600 728 29900 6 Bit_In
port 2 nsew signal input
rlabel metal2 s 22176 100 22232 400 6 EN
port 3 nsew signal input
rlabel metal3 s 29600 3360 29900 3416 6 I[0]
port 4 nsew signal output
rlabel metal3 s 100 22176 400 22232 6 I[10]
port 5 nsew signal output
rlabel metal3 s 29600 672 29900 728 6 I[11]
port 6 nsew signal output
rlabel metal2 s 27888 100 27944 400 6 I[12]
port 7 nsew signal output
rlabel metal3 s 29600 20160 29900 20216 6 I[1]
port 8 nsew signal output
rlabel metal2 s 11088 100 11144 400 6 I[2]
port 9 nsew signal output
rlabel metal2 s 16800 100 16856 400 6 I[3]
port 10 nsew signal output
rlabel metal2 s 23184 29600 23240 29900 6 I[4]
port 11 nsew signal output
rlabel metal3 s 100 11088 400 11144 6 I[5]
port 12 nsew signal output
rlabel metal3 s 29600 23184 29900 23240 6 I[6]
port 13 nsew signal output
rlabel metal3 s 100 16800 400 16856 6 I[7]
port 14 nsew signal output
rlabel metal2 s 5376 100 5432 400 6 I[8]
port 15 nsew signal output
rlabel metal3 s 100 19488 400 19544 6 I[9]
port 16 nsew signal output
rlabel metal3 s 100 8400 400 8456 6 Q[0]
port 17 nsew signal output
rlabel metal2 s 17472 29600 17528 29900 6 Q[10]
port 18 nsew signal output
rlabel metal2 s 25872 29600 25928 29900 6 Q[11]
port 19 nsew signal output
rlabel metal3 s 29600 9072 29900 9128 6 Q[12]
port 20 nsew signal output
rlabel metal3 s 29600 25872 29900 25928 6 Q[1]
port 21 nsew signal output
rlabel metal2 s 6048 29600 6104 29900 6 Q[2]
port 22 nsew signal output
rlabel metal2 s 0 100 56 400 6 Q[3]
port 23 nsew signal output
rlabel metal3 s 100 5376 400 5432 6 Q[4]
port 24 nsew signal output
rlabel metal3 s 29600 17472 29900 17528 6 Q[5]
port 25 nsew signal output
rlabel metal2 s 3360 29600 3416 29900 6 Q[6]
port 26 nsew signal output
rlabel metal3 s 100 2688 400 2744 6 Q[7]
port 27 nsew signal output
rlabel metal2 s 25200 100 25256 400 6 Q[8]
port 28 nsew signal output
rlabel metal2 s 20160 29600 20216 29900 6 Q[9]
port 29 nsew signal output
rlabel metal3 s 29600 6048 29900 6104 6 REQ_SAMPLE
port 30 nsew signal input
rlabel metal2 s 2688 100 2744 400 6 RST
port 31 nsew signal input
rlabel metal2 s 8400 100 8456 400 6 addI[0]
port 32 nsew signal output
rlabel metal3 s 100 25200 400 25256 6 addI[1]
port 33 nsew signal output
rlabel metal3 s 29600 11760 29900 11816 6 addI[2]
port 34 nsew signal output
rlabel metal2 s 13776 100 13832 400 6 addI[3]
port 35 nsew signal output
rlabel metal3 s 29600 28560 29900 28616 6 addI[4]
port 36 nsew signal output
rlabel metal2 s 28560 29600 28616 29900 6 addI[5]
port 37 nsew signal output
rlabel metal2 s 9072 29600 9128 29900 6 addQ[0]
port 38 nsew signal output
rlabel metal2 s 11760 29600 11816 29900 6 addQ[1]
port 39 nsew signal output
rlabel metal2 s 19488 100 19544 400 6 addQ[2]
port 40 nsew signal output
rlabel metal3 s 100 13776 400 13832 6 addQ[3]
port 41 nsew signal output
rlabel metal3 s 100 27888 400 27944 6 addQ[4]
port 42 nsew signal output
rlabel metal3 s 29600 14448 29900 14504 6 addQ[5]
port 43 nsew signal output
rlabel metal4 s 2224 1538 2384 28254 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 28254 6 vdd
port 44 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 28254 6 vss
port 45 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 28254 6 vss
port 45 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3565500
string GDS_FILE /home/urielcho/Proyectos_caravel/gf180nm/modulador_a/openlane/modulador_a/runs/22_12_04_18_07/results/signoff/OQPSK_RCOSINE_ALL.magic.gds
string GDS_START 337848
<< end >>

