VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OQPSK_RCOSINE_ALL
  CLASS BLOCK ;
  FOREIGN OQPSK_RCOSINE_ALL ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN ACK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 296.000 145.040 299.000 ;
    END
  END ACK
  PIN Bit_In
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 296.000 7.280 299.000 ;
    END
  END Bit_In
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 1.000 222.320 4.000 ;
    END
  END EN
  PIN I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 33.600 299.000 34.160 ;
    END
  END I[0]
  PIN I[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 221.760 4.000 222.320 ;
    END
  END I[10]
  PIN I[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 6.720 299.000 7.280 ;
    END
  END I[11]
  PIN I[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 1.000 279.440 4.000 ;
    END
  END I[12]
  PIN I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 201.600 299.000 202.160 ;
    END
  END I[1]
  PIN I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 1.000 111.440 4.000 ;
    END
  END I[2]
  PIN I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 1.000 168.560 4.000 ;
    END
  END I[3]
  PIN I[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 296.000 232.400 299.000 ;
    END
  END I[4]
  PIN I[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 110.880 4.000 111.440 ;
    END
  END I[5]
  PIN I[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 231.840 299.000 232.400 ;
    END
  END I[6]
  PIN I[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 168.000 4.000 168.560 ;
    END
  END I[7]
  PIN I[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 1.000 54.320 4.000 ;
    END
  END I[8]
  PIN I[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 194.880 4.000 195.440 ;
    END
  END I[9]
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 84.000 4.000 84.560 ;
    END
  END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 296.000 175.280 299.000 ;
    END
  END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 296.000 259.280 299.000 ;
    END
  END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 90.720 299.000 91.280 ;
    END
  END Q[12]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 258.720 299.000 259.280 ;
    END
  END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 296.000 61.040 299.000 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 53.760 4.000 54.320 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 174.720 299.000 175.280 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 296.000 34.160 299.000 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 26.880 4.000 27.440 ;
    END
  END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 1.000 252.560 4.000 ;
    END
  END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 296.000 202.160 299.000 ;
    END
  END Q[9]
  PIN REQ_SAMPLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 60.480 299.000 61.040 ;
    END
  END REQ_SAMPLE
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 1.000 27.440 4.000 ;
    END
  END RST
  PIN addI[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 1.000 84.560 4.000 ;
    END
  END addI[0]
  PIN addI[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 252.000 4.000 252.560 ;
    END
  END addI[1]
  PIN addI[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 117.600 299.000 118.160 ;
    END
  END addI[2]
  PIN addI[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 137.760 1.000 138.320 4.000 ;
    END
  END addI[3]
  PIN addI[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 285.600 299.000 286.160 ;
    END
  END addI[4]
  PIN addI[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 296.000 286.160 299.000 ;
    END
  END addI[5]
  PIN addQ[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 296.000 91.280 299.000 ;
    END
  END addQ[0]
  PIN addQ[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 296.000 118.160 299.000 ;
    END
  END addQ[1]
  PIN addQ[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 1.000 195.440 4.000 ;
    END
  END addQ[2]
  PIN addQ[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 137.760 4.000 138.320 ;
    END
  END addQ[3]
  PIN addQ[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 278.880 4.000 279.440 ;
    END
  END addQ[4]
  PIN addQ[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 144.480 299.000 145.040 ;
    END
  END addQ[5]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 292.880 283.210 ;
      LAYER Metal2 ;
        RECT 0.140 295.700 6.420 296.000 ;
        RECT 7.580 295.700 33.300 296.000 ;
        RECT 34.460 295.700 60.180 296.000 ;
        RECT 61.340 295.700 90.420 296.000 ;
        RECT 91.580 295.700 117.300 296.000 ;
        RECT 118.460 295.700 144.180 296.000 ;
        RECT 145.340 295.700 174.420 296.000 ;
        RECT 175.580 295.700 201.300 296.000 ;
        RECT 202.460 295.700 231.540 296.000 ;
        RECT 232.700 295.700 258.420 296.000 ;
        RECT 259.580 295.700 285.300 296.000 ;
        RECT 286.460 295.700 297.220 296.000 ;
        RECT 0.140 4.300 297.220 295.700 ;
        RECT 0.860 4.000 26.580 4.300 ;
        RECT 27.740 4.000 53.460 4.300 ;
        RECT 54.620 4.000 83.700 4.300 ;
        RECT 84.860 4.000 110.580 4.300 ;
        RECT 111.740 4.000 137.460 4.300 ;
        RECT 138.620 4.000 167.700 4.300 ;
        RECT 168.860 4.000 194.580 4.300 ;
        RECT 195.740 4.000 221.460 4.300 ;
        RECT 222.620 4.000 251.700 4.300 ;
        RECT 252.860 4.000 278.580 4.300 ;
        RECT 279.740 4.000 297.220 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 286.460 297.270 292.740 ;
        RECT 0.090 285.300 295.700 286.460 ;
        RECT 0.090 279.740 297.270 285.300 ;
        RECT 0.090 278.580 0.700 279.740 ;
        RECT 4.300 278.580 297.270 279.740 ;
        RECT 0.090 259.580 297.270 278.580 ;
        RECT 0.090 258.420 295.700 259.580 ;
        RECT 0.090 252.860 297.270 258.420 ;
        RECT 0.090 251.700 0.700 252.860 ;
        RECT 4.300 251.700 297.270 252.860 ;
        RECT 0.090 232.700 297.270 251.700 ;
        RECT 0.090 231.540 295.700 232.700 ;
        RECT 0.090 222.620 297.270 231.540 ;
        RECT 0.090 221.460 0.700 222.620 ;
        RECT 4.300 221.460 297.270 222.620 ;
        RECT 0.090 202.460 297.270 221.460 ;
        RECT 0.090 201.300 295.700 202.460 ;
        RECT 0.090 195.740 297.270 201.300 ;
        RECT 0.090 194.580 0.700 195.740 ;
        RECT 4.300 194.580 297.270 195.740 ;
        RECT 0.090 175.580 297.270 194.580 ;
        RECT 0.090 174.420 295.700 175.580 ;
        RECT 0.090 168.860 297.270 174.420 ;
        RECT 0.090 167.700 0.700 168.860 ;
        RECT 4.300 167.700 297.270 168.860 ;
        RECT 0.090 145.340 297.270 167.700 ;
        RECT 0.090 144.180 295.700 145.340 ;
        RECT 0.090 138.620 297.270 144.180 ;
        RECT 0.090 137.460 0.700 138.620 ;
        RECT 4.300 137.460 297.270 138.620 ;
        RECT 0.090 118.460 297.270 137.460 ;
        RECT 0.090 117.300 295.700 118.460 ;
        RECT 0.090 111.740 297.270 117.300 ;
        RECT 0.090 110.580 0.700 111.740 ;
        RECT 4.300 110.580 297.270 111.740 ;
        RECT 0.090 91.580 297.270 110.580 ;
        RECT 0.090 90.420 295.700 91.580 ;
        RECT 0.090 84.860 297.270 90.420 ;
        RECT 0.090 83.700 0.700 84.860 ;
        RECT 4.300 83.700 297.270 84.860 ;
        RECT 0.090 61.340 297.270 83.700 ;
        RECT 0.090 60.180 295.700 61.340 ;
        RECT 0.090 54.620 297.270 60.180 ;
        RECT 0.090 53.460 0.700 54.620 ;
        RECT 4.300 53.460 297.270 54.620 ;
        RECT 0.090 34.460 297.270 53.460 ;
        RECT 0.090 33.300 295.700 34.460 ;
        RECT 0.090 27.740 297.270 33.300 ;
        RECT 0.090 26.580 0.700 27.740 ;
        RECT 4.300 26.580 297.270 27.740 ;
        RECT 0.090 7.580 297.270 26.580 ;
        RECT 0.090 6.860 295.700 7.580 ;
      LAYER Metal4 ;
        RECT 10.780 282.840 286.020 292.790 ;
        RECT 10.780 15.080 21.940 282.840 ;
        RECT 24.140 15.080 98.740 282.840 ;
        RECT 100.940 15.080 175.540 282.840 ;
        RECT 177.740 15.080 252.340 282.840 ;
        RECT 254.540 15.080 286.020 282.840 ;
        RECT 10.780 7.370 286.020 15.080 ;
  END
END OQPSK_RCOSINE_ALL
END LIBRARY

