// This is the unpowered netlist.
module OQPSK_RCOSINE_ALL (ACK,
    Bit_In,
    EN,
    REQ_SAMPLE,
    RST,
    I,
    Q,
    addI,
    addQ);
 input ACK;
 input Bit_In;
 input EN;
 input REQ_SAMPLE;
 input RST;
 output [12:0] I;
 output [12:0] Q;
 output [5:0] addI;
 output [5:0] addQ;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire \gen_sym.Reg_2M.data_in ;
 wire \gen_sym.Reg_2M.data_out ;
 wire \gen_sym.Reg_2M.enable ;
 wire \gen_sym.Reg_Sym.data_out[0] ;
 wire \gen_sym.Reg_Sym.data_out[1] ;
 wire \mapper.bit_Q[1] ;
 wire \p_shaping_I.p_shaping_I.bit_in ;
 wire \p_shaping_I.p_shaping_I.bit_in_1 ;
 wire \p_shaping_I.p_shaping_I.bit_in_2 ;
 wire \p_shaping_I.p_shaping_I.counter[0] ;
 wire \p_shaping_I.p_shaping_I.counter[1] ;
 wire \p_shaping_I.p_shaping_I.ctl_1 ;
 wire \p_shaping_Q.p_shaping_I.bit_in ;
 wire \p_shaping_Q.p_shaping_I.bit_in_1 ;
 wire \p_shaping_Q.p_shaping_I.bit_in_2 ;
 wire \p_shaping_Q.p_shaping_I.counter[0] ;
 wire \p_shaping_Q.p_shaping_I.counter[1] ;
 wire \p_shaping_Q.p_shaping_I.ctl_1 ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1346_ (.I(net35),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1347_ (.I(net34),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1348_ (.I(_1181_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1349_ (.A1(_1170_),
    .A2(_1192_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1350_ (.I(net35),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1351_ (.I(_1214_),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1352_ (.I(net33),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1353_ (.I(_1236_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1354_ (.I(net32),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1355_ (.I(_1258_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1356_ (.I(_1181_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1357_ (.A1(_1247_),
    .A2(_1268_),
    .A3(_1279_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1358_ (.A1(_1225_),
    .A2(_1290_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1359_ (.I(net36),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1360_ (.I(net37),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1361_ (.I(_1323_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1362_ (.A1(_1312_),
    .A2(_1334_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1363_ (.A1(_1203_),
    .A2(_1301_),
    .B(_1345_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1364_ (.I(net37),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1365_ (.I(_1236_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1366_ (.I(net36),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1367_ (.A1(_0054_),
    .A2(_1170_),
    .A3(_1279_),
    .B(_0065_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1368_ (.A1(_0043_),
    .A2(_0074_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1369_ (.I(_1214_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1370_ (.I(net36),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1371_ (.I(net37),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1372_ (.I(net33),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1373_ (.I(net34),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1374_ (.A1(_0129_),
    .A2(_0140_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1375_ (.A1(_0096_),
    .A2(_0107_),
    .A3(_0118_),
    .A4(_0150_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1376_ (.A1(_0085_),
    .A2(_0161_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1377_ (.A1(_0032_),
    .A2(_0172_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1378_ (.I(_1268_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1379_ (.I(_0194_),
    .Z(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1380_ (.I(_0129_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1381_ (.I(net35),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1382_ (.I(_0226_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1383_ (.I(_0140_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1384_ (.A1(_0215_),
    .A2(_0237_),
    .A3(_0248_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1385_ (.A1(_0204_),
    .A2(_0258_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1386_ (.A1(_0183_),
    .A2(_0269_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1387_ (.I(_0280_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1388_ (.I(_0291_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1389_ (.I(net38),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1390_ (.I(_0311_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1391_ (.I(_0322_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1392_ (.I(net39),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1393_ (.I(net41),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1394_ (.I(_0355_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1395_ (.I(net51),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1396_ (.A1(_0344_),
    .A2(_0365_),
    .A3(_0376_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1397_ (.I(_0387_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1398_ (.I(_0355_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1399_ (.I(net51),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1400_ (.A1(_0344_),
    .A2(_0311_),
    .A3(_0418_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1401_ (.A1(_0408_),
    .A2(_0429_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1402_ (.I(net50),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1403_ (.I(net41),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1404_ (.I(net51),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1405_ (.A1(_0460_),
    .A2(_0468_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1406_ (.A1(_0450_),
    .A2(_0476_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1407_ (.A1(_0440_),
    .A2(_0484_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1408_ (.I(net43),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1409_ (.A1(_0450_),
    .A2(_0387_),
    .B(_0498_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1410_ (.I(net39),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1411_ (.A1(_0500_),
    .A2(net51),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1412_ (.A1(_0460_),
    .A2(net50),
    .A3(_0501_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1413_ (.A1(_0498_),
    .A2(_0502_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1414_ (.A1(_0491_),
    .A2(_0499_),
    .B(_0503_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1415_ (.A1(_0333_),
    .A2(_0397_),
    .A3(_0504_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1416_ (.I(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1417_ (.I(_0506_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1418_ (.I(net1),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1419_ (.A1(\gen_sym.Reg_Sym.data_out[1] ),
    .A2(_0507_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1420_ (.I(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1421_ (.I(_0509_),
    .Z(\p_shaping_I.p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1422_ (.A1(_0507_),
    .A2(\gen_sym.Reg_Sym.data_out[0] ),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1423_ (.I(_0510_),
    .Z(\mapper.bit_Q[1] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1424_ (.I(\p_shaping_I.p_shaping_I.bit_in_1 ),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1425_ (.I(_0511_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1426_ (.I(_0512_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1427_ (.I(net53),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1428_ (.I(_0508_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1429_ (.I(_0515_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1430_ (.A1(\p_shaping_I.p_shaping_I.ctl_1 ),
    .A2(_0514_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1431_ (.A1(_0514_),
    .A2(_0516_),
    .B(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1432_ (.A1(_0291_),
    .A2(_0518_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1433_ (.A1(_0513_),
    .A2(net45),
    .B(_0519_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1434_ (.I(\p_shaping_Q.p_shaping_I.bit_in_1 ),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1435_ (.I(_0520_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1436_ (.I(net44),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1437_ (.I(_0522_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1438_ (.A1(net59),
    .A2(\p_shaping_Q.p_shaping_I.ctl_1 ),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1439_ (.A1(_0514_),
    .A2(_0523_),
    .B(_0524_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1440_ (.A1(_0505_),
    .A2(_0525_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1441_ (.A1(_0521_),
    .A2(_0505_),
    .B(_0526_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1442_ (.A1(net3),
    .A2(net2),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1443_ (.I(_0527_),
    .Z(\gen_sym.Reg_2M.data_in ));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1444_ (.A1(_0291_),
    .A2(net48),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1445_ (.I(_0528_),
    .Z(\gen_sym.Reg_2M.enable ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1446_ (.I(_0514_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1447_ (.A1(_0529_),
    .A2(net45),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1448_ (.A1(_0529_),
    .A2(net49),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1449_ (.I(\p_shaping_Q.p_shaping_I.counter[1] ),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1450_ (.I(_0530_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1451_ (.I(_0531_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1452_ (.I(net50),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1453_ (.I(_0533_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1454_ (.I(net39),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1455_ (.A1(_0535_),
    .A2(_0311_),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1456_ (.I(_0536_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1457_ (.I(_0365_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1458_ (.I(net43),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1459_ (.A1(_0538_),
    .A2(_0539_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1460_ (.I(_0468_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1461_ (.I(_0541_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1462_ (.I(_0542_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1463_ (.A1(_0537_),
    .A2(_0540_),
    .B(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1464_ (.I(net38),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1465_ (.I(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1466_ (.I(_0546_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1467_ (.I(_0418_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1468_ (.I(_0548_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1469_ (.I(_0408_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1470_ (.I(_0535_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1471_ (.I(_0551_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1472_ (.A1(_0547_),
    .A2(_0549_),
    .B(_0550_),
    .C(_0552_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1473_ (.I(_0460_),
    .Z(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1474_ (.I(_0554_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1475_ (.A1(_0535_),
    .A2(_0468_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1476_ (.I(_0556_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1477_ (.A1(_0333_),
    .A2(_0555_),
    .A3(_0557_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1478_ (.I(net50),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1479_ (.I(_0559_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1480_ (.I(_0560_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1481_ (.I(_0500_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1482_ (.I(_0562_),
    .Z(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1483_ (.I(_0545_),
    .Z(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1484_ (.I(_0564_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1485_ (.I(_0460_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1486_ (.I(_0418_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1487_ (.A1(_0563_),
    .A2(_0565_),
    .B(_0566_),
    .C(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1488_ (.A1(_0561_),
    .A2(_0568_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1489_ (.A1(_0534_),
    .A2(_0544_),
    .A3(_0553_),
    .B1(_0558_),
    .B2(_0569_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1490_ (.I(_0355_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1491_ (.I(_0554_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1492_ (.I(_0450_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1493_ (.A1(_0572_),
    .A2(_0573_),
    .B(_0539_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1494_ (.A1(_0571_),
    .A2(_0537_),
    .B(_0574_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1495_ (.I(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1496_ (.A1(_0570_),
    .A2(_0576_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1497_ (.A1(_0532_),
    .A2(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1498_ (.I(net43),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1499_ (.I(_0579_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1500_ (.A1(_0554_),
    .A2(_0556_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1501_ (.A1(_0500_),
    .A2(net38),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1502_ (.I(_0551_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1503_ (.A1(_0583_),
    .A2(_0322_),
    .B(_0542_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1504_ (.I(_0418_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1505_ (.A1(_0344_),
    .A2(_0311_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1506_ (.I(_0355_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1507_ (.A1(_0585_),
    .A2(_0586_),
    .B(_0587_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1508_ (.A1(_0581_),
    .A2(_0582_),
    .B1(_0584_),
    .B2(_0588_),
    .C(_0533_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1509_ (.I(_0587_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1510_ (.I(_0545_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1511_ (.A1(_0591_),
    .A2(_0585_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1512_ (.A1(_0344_),
    .A2(_0376_),
    .B(_0365_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1513_ (.A1(_0536_),
    .A2(_0593_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1514_ (.A1(_0590_),
    .A2(_0592_),
    .B(_0594_),
    .C(_0560_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1515_ (.A1(_0562_),
    .A2(_0564_),
    .A3(_0365_),
    .A4(_0376_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1516_ (.A1(_0533_),
    .A2(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1517_ (.A1(_0539_),
    .A2(_0597_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1518_ (.A1(_0583_),
    .A2(_0567_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1519_ (.I(_0535_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1520_ (.I(_0408_),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1521_ (.I(_0541_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _1522_ (.A1(_0600_),
    .A2(_0601_),
    .A3(_0602_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1523_ (.A1(_0583_),
    .A2(_0567_),
    .B(_0538_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1524_ (.A1(_0599_),
    .A2(_0603_),
    .A3(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1525_ (.A1(_0580_),
    .A2(_0589_),
    .A3(_0595_),
    .B1(_0598_),
    .B2(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1526_ (.A1(\p_shaping_Q.p_shaping_I.counter[0] ),
    .A2(\p_shaping_Q.p_shaping_I.counter[1] ),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1527_ (.I(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1528_ (.I(_0608_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1529_ (.A1(_0606_),
    .A2(_0609_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1530_ (.I(_0610_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1531_ (.I(_0539_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1532_ (.I(_0584_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1533_ (.I(_0468_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1534_ (.I(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1535_ (.A1(_0547_),
    .A2(_0615_),
    .B(_0555_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1536_ (.I0(_0591_),
    .I1(_0600_),
    .S(_0376_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1537_ (.A1(_0590_),
    .A2(_0617_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1538_ (.I(_0586_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1539_ (.I(_0559_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1540_ (.A1(_0564_),
    .A2(_0614_),
    .B(_0587_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1541_ (.A1(_0620_),
    .A2(_0621_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1542_ (.A1(_0613_),
    .A2(_0616_),
    .B1(_0618_),
    .B2(_0619_),
    .C(_0622_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1543_ (.I(_0601_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1544_ (.A1(_0500_),
    .A2(_0545_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1545_ (.A1(_0600_),
    .A2(_0322_),
    .A3(_0585_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1546_ (.A1(_0602_),
    .A2(_0625_),
    .B(_0626_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1547_ (.A1(_0552_),
    .A2(_0601_),
    .A3(_0615_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1548_ (.I(_0450_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1549_ (.I(_0498_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1550_ (.A1(_0629_),
    .A2(_0630_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1551_ (.A1(_0624_),
    .A2(_0627_),
    .B(_0628_),
    .C(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1552_ (.A1(_0561_),
    .A2(_0630_),
    .A3(_0397_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1553_ (.A1(_0612_),
    .A2(_0623_),
    .B(_0632_),
    .C(_0633_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1554_ (.I(_0634_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1555_ (.A1(_0611_),
    .A2(_0635_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1556_ (.A1(_0578_),
    .A2(_0636_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1557_ (.I(_0637_),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1558_ (.A1(_0611_),
    .A2(_0635_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1559_ (.A1(_0578_),
    .A2(_0636_),
    .B(_0638_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1560_ (.I(_0608_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1561_ (.I(_0520_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1562_ (.A1(_0641_),
    .A2(_0606_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1563_ (.A1(_0573_),
    .A2(_0397_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1564_ (.A1(_0548_),
    .A2(_0625_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1565_ (.A1(_0591_),
    .A2(_0585_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1566_ (.A1(_0557_),
    .A2(_0645_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1567_ (.A1(_0555_),
    .A2(_0557_),
    .B1(_0644_),
    .B2(_0646_),
    .C(_0620_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1568_ (.I(_0630_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1569_ (.A1(_0643_),
    .A2(_0647_),
    .B(_0648_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1570_ (.A1(_0562_),
    .A2(_0591_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1571_ (.A1(_0567_),
    .A2(_0650_),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1572_ (.I(_0546_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1573_ (.A1(_0563_),
    .A2(_0652_),
    .B(_0542_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1574_ (.A1(_0651_),
    .A2(_0653_),
    .B(_0550_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1575_ (.A1(_0546_),
    .A2(_0614_),
    .B(_0408_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1576_ (.A1(_0655_),
    .A2(_0584_),
    .B(_0629_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1577_ (.A1(_0555_),
    .A2(_0626_),
    .B(_0561_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1578_ (.I(_0579_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1579_ (.A1(_0654_),
    .A2(_0656_),
    .B1(_0657_),
    .B2(_0603_),
    .C(_0658_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1580_ (.A1(_0649_),
    .A2(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1581_ (.A1(_0642_),
    .A2(_0660_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1582_ (.A1(_0640_),
    .A2(_0661_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1583_ (.I(_0566_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1584_ (.I(_0562_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1585_ (.A1(_0664_),
    .A2(_0615_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1586_ (.I(_0625_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1587_ (.A1(_0663_),
    .A2(_0665_),
    .A3(_0666_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1588_ (.A1(_0534_),
    .A2(_0618_),
    .A3(_0667_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1589_ (.I(_0542_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1590_ (.A1(_0664_),
    .A2(_0669_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1591_ (.I(_0600_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1592_ (.A1(_0671_),
    .A2(_0652_),
    .B(_0550_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1593_ (.I(_0501_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1594_ (.A1(_0572_),
    .A2(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1595_ (.A1(_0670_),
    .A2(_0672_),
    .B(_0534_),
    .C(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1596_ (.I(_0652_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1597_ (.A1(_0671_),
    .A2(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1598_ (.I(_0566_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1599_ (.A1(_0678_),
    .A2(_0626_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1600_ (.A1(_0533_),
    .A2(_0579_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1601_ (.I(_0680_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1602_ (.A1(_0571_),
    .A2(_0677_),
    .B(_0679_),
    .C(_0681_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1603_ (.A1(_0648_),
    .A2(_0668_),
    .B(_0675_),
    .C(_0682_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1604_ (.A1(net44),
    .A2(_0635_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1605_ (.A1(_0683_),
    .A2(_0684_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1606_ (.I(\p_shaping_Q.p_shaping_I.bit_in_2 ),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1607_ (.A1(_0686_),
    .A2(_0577_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1608_ (.I(_0596_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1609_ (.A1(_0534_),
    .A2(_0688_),
    .B(_0648_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1610_ (.A1(_0566_),
    .A2(_0548_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1611_ (.I(_0690_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1612_ (.I(_0537_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1613_ (.A1(_0671_),
    .A2(_0676_),
    .B(_0543_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1614_ (.I(_0663_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1615_ (.I(_0694_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1616_ (.A1(_0691_),
    .A2(_0692_),
    .B1(_0693_),
    .B2(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1617_ (.A1(_0549_),
    .A2(_0666_),
    .B(_0572_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1618_ (.I(_0697_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1619_ (.I(_0560_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1620_ (.I(_0699_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1621_ (.I(_0700_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1622_ (.A1(_0618_),
    .A2(_0698_),
    .B(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1623_ (.I(_0580_),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1624_ (.I(_0703_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1625_ (.I(_0620_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1626_ (.I(_0582_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1627_ (.A1(_0624_),
    .A2(_0705_),
    .A3(_0706_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1628_ (.A1(_0704_),
    .A2(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1629_ (.A1(_0689_),
    .A2(_0696_),
    .B1(_0702_),
    .B2(_0708_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1630_ (.A1(_0687_),
    .A2(_0709_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1631_ (.A1(_0531_),
    .A2(_0710_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1632_ (.A1(_0662_),
    .A2(_0685_),
    .A3(_0711_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1633_ (.A1(_0639_),
    .A2(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1634_ (.I(_0640_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1635_ (.A1(_0007_),
    .A2(_0661_),
    .B(_0685_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1636_ (.A1(_0007_),
    .A2(_0661_),
    .A3(_0685_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1637_ (.A1(_0714_),
    .A2(_0711_),
    .B(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1638_ (.A1(_0522_),
    .A2(_0524_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1639_ (.A1(_0506_),
    .A2(_0717_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1640_ (.I(_0648_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1641_ (.I(_0629_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1642_ (.I(_0322_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1643_ (.A1(_0721_),
    .A2(_0397_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1644_ (.A1(_0678_),
    .A2(_0669_),
    .A3(_0706_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1645_ (.A1(_0664_),
    .A2(_0621_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1646_ (.A1(_0720_),
    .A2(_0722_),
    .B(_0723_),
    .C(_0724_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1647_ (.I(_0565_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1648_ (.A1(_0554_),
    .A2(_0556_),
    .Z(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1649_ (.A1(_0620_),
    .A2(_0630_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1650_ (.A1(_0726_),
    .A2(_0580_),
    .A3(_0727_),
    .B(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1651_ (.A1(_0564_),
    .A2(_0587_),
    .A3(_0614_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1652_ (.A1(_0538_),
    .A2(_0602_),
    .A3(_0582_),
    .B(_0730_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1653_ (.A1(_0573_),
    .A2(_0724_),
    .A3(_0731_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1654_ (.A1(_0729_),
    .A2(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1655_ (.A1(_0719_),
    .A2(_0725_),
    .B(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1656_ (.A1(_0606_),
    .A2(_0649_),
    .A3(_0659_),
    .B(_0520_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1657_ (.A1(_0718_),
    .A2(_0734_),
    .A3(_0735_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1658_ (.A1(_0609_),
    .A2(_0736_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1659_ (.A1(_0726_),
    .A2(_0673_),
    .A3(_0727_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1660_ (.I(_0655_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1661_ (.A1(_0739_),
    .A2(_0599_),
    .B(_0644_),
    .C(_0658_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1662_ (.A1(_0671_),
    .A2(_0547_),
    .A3(_0678_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1663_ (.I(_0557_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1664_ (.A1(_0563_),
    .A2(_0565_),
    .B(_0538_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1665_ (.A1(_0721_),
    .A2(_0742_),
    .B(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1666_ (.A1(_0741_),
    .A2(_0744_),
    .B(_0658_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1667_ (.A1(_0728_),
    .A2(_0738_),
    .B1(_0740_),
    .B2(_0705_),
    .C(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1668_ (.A1(_0635_),
    .A2(_0683_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1669_ (.A1(net44),
    .A2(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1670_ (.A1(_0746_),
    .A2(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1671_ (.A1(_0570_),
    .A2(_0576_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1672_ (.I(\p_shaping_Q.p_shaping_I.bit_in_2 ),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1673_ (.A1(_0750_),
    .A2(_0709_),
    .B(_0751_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1674_ (.A1(_0561_),
    .A2(_0580_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1675_ (.I0(_0613_),
    .I1(_0645_),
    .S(_0571_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1676_ (.A1(_0550_),
    .A2(_0549_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1677_ (.A1(_0669_),
    .A2(_0586_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1678_ (.A1(_0552_),
    .A2(_0333_),
    .B(_0678_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1679_ (.A1(_0560_),
    .A2(_0579_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1680_ (.I(_0758_),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1681_ (.A1(_0619_),
    .A2(_0755_),
    .B1(_0756_),
    .B2(_0757_),
    .C(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1682_ (.I(_0583_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1683_ (.A1(_0761_),
    .A2(_0726_),
    .A3(_0476_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1684_ (.A1(_0624_),
    .A2(_0645_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1685_ (.A1(_0693_),
    .A2(_0681_),
    .A3(_0762_),
    .A4(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1686_ (.A1(_0753_),
    .A2(_0754_),
    .B(_0760_),
    .C(_0764_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1687_ (.A1(_0752_),
    .A2(_0765_),
    .B(\p_shaping_Q.p_shaping_I.counter[1] ),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1688_ (.A1(_0752_),
    .A2(_0765_),
    .B(_0766_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1689_ (.A1(_0737_),
    .A2(_0749_),
    .A3(_0767_),
    .Z(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1690_ (.A1(_0713_),
    .A2(_0716_),
    .A3(_0768_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1691_ (.I(_0769_),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1692_ (.A1(_0716_),
    .A2(_0768_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1693_ (.A1(_0716_),
    .A2(_0768_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1694_ (.A1(_0639_),
    .A2(_0712_),
    .A3(_0770_),
    .B(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1695_ (.A1(_0737_),
    .A2(_0749_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1696_ (.I(_0767_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1697_ (.A1(_0737_),
    .A2(_0749_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1698_ (.A1(_0773_),
    .A2(_0774_),
    .B(_0775_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1699_ (.I(_0548_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1700_ (.A1(_0726_),
    .A2(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1701_ (.A1(_0602_),
    .A2(_0625_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1702_ (.A1(_0778_),
    .A2(_0670_),
    .A3(_0672_),
    .A4(_0779_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1703_ (.A1(_0670_),
    .A2(_0672_),
    .B1(_0779_),
    .B2(_0778_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1704_ (.A1(_0631_),
    .A2(_0780_),
    .A3(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1705_ (.I(_0777_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1706_ (.I(_0582_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1707_ (.A1(_0783_),
    .A2(_0784_),
    .B(_0429_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1708_ (.A1(_0618_),
    .A2(_0785_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1709_ (.A1(_0628_),
    .A2(_0681_),
    .A3(_0730_),
    .Z(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1710_ (.A1(_0786_),
    .A2(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1711_ (.I(_0601_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1712_ (.A1(_0552_),
    .A2(_0777_),
    .B(_0789_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1713_ (.I(_0653_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1714_ (.A1(_0790_),
    .A2(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1715_ (.I(_0565_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1716_ (.I(_0669_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1717_ (.I(_0590_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1718_ (.A1(_0793_),
    .A2(_0794_),
    .B(_0795_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1719_ (.A1(_0692_),
    .A2(_0796_),
    .B(_0665_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1720_ (.A1(_0792_),
    .A2(_0797_),
    .B(_0759_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1721_ (.A1(_0782_),
    .A2(_0788_),
    .A3(_0798_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1722_ (.A1(_0624_),
    .A2(_0617_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1723_ (.A1(_0720_),
    .A2(_0723_),
    .A3(_0800_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1724_ (.A1(_0476_),
    .A2(_0650_),
    .B1(_0757_),
    .B2(_0794_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1725_ (.A1(_0703_),
    .A2(_0801_),
    .A3(_0707_),
    .B1(_0598_),
    .B2(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1726_ (.A1(_0577_),
    .A2(_0803_),
    .A3(_0765_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1727_ (.A1(_0686_),
    .A2(_0804_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1728_ (.A1(_0799_),
    .A2(_0805_),
    .B(_0530_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1729_ (.A1(_0799_),
    .A2(_0805_),
    .B(_0806_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1730_ (.I(_0607_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1731_ (.I(_0563_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1732_ (.I(_0621_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1733_ (.A1(_0615_),
    .A2(_0666_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1734_ (.A1(_0652_),
    .A2(_0590_),
    .A3(_0501_),
    .B(_0629_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1735_ (.A1(_0809_),
    .A2(_0810_),
    .B1(_0811_),
    .B2(_0571_),
    .C(_0812_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1736_ (.A1(_0612_),
    .A2(_0813_),
    .B1(_0729_),
    .B2(_0732_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1737_ (.A1(_0606_),
    .A2(_0649_),
    .A3(_0659_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1738_ (.A1(_0543_),
    .A2(_0706_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1739_ (.A1(_0549_),
    .A2(_0537_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1740_ (.A1(_0795_),
    .A2(_0816_),
    .A3(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1741_ (.A1(_0689_),
    .A2(_0628_),
    .A3(_0818_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1742_ (.A1(_0721_),
    .A2(_0663_),
    .A3(_0742_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1743_ (.A1(_0789_),
    .A2(_0592_),
    .B(_0699_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1744_ (.A1(_0820_),
    .A2(_0821_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1745_ (.A1(_0790_),
    .A2(_0791_),
    .B1(_0779_),
    .B2(_0604_),
    .C(_0699_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1746_ (.A1(_0822_),
    .A2(_0823_),
    .B(_0703_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1747_ (.A1(_0819_),
    .A2(_0824_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1748_ (.A1(_0814_),
    .A2(_0815_),
    .B(_0825_),
    .C(_0641_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1749_ (.A1(_0819_),
    .A2(_0824_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1750_ (.A1(_0641_),
    .A2(_0814_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1751_ (.A1(_0735_),
    .A2(_0827_),
    .A3(_0828_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1752_ (.A1(_0506_),
    .A2(_0717_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1753_ (.A1(_0826_),
    .A2(_0829_),
    .B(_0830_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1754_ (.I(_0831_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1755_ (.I(_0718_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1756_ (.I(_0833_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1757_ (.I(_0735_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1758_ (.A1(_0835_),
    .A2(_0828_),
    .B(_0827_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1759_ (.A1(_0835_),
    .A2(_0827_),
    .A3(_0828_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1760_ (.A1(_0834_),
    .A2(_0836_),
    .A3(_0837_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1761_ (.I(\p_shaping_Q.p_shaping_I.bit_in ),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1762_ (.A1(_0746_),
    .A2(_0747_),
    .B(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1763_ (.A1(_0650_),
    .A2(_0739_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1764_ (.A1(_0793_),
    .A2(_0673_),
    .B1(_0691_),
    .B2(_0692_),
    .C(_0758_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1765_ (.A1(_0789_),
    .A2(_0592_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1766_ (.A1(_0820_),
    .A2(_0843_),
    .A3(_0628_),
    .A4(_0681_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1767_ (.A1(_0663_),
    .A2(_0777_),
    .A3(_0666_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1768_ (.A1(_0706_),
    .A2(_0810_),
    .B(_0699_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1769_ (.A1(_0845_),
    .A2(_0846_),
    .B(_0658_),
    .C(_0722_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1770_ (.A1(_0841_),
    .A2(_0842_),
    .B(_0844_),
    .C(_0847_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1771_ (.A1(_0840_),
    .A2(_0848_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1772_ (.A1(_0808_),
    .A2(_0832_),
    .A3(_0838_),
    .A4(_0849_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1773_ (.I(_0831_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1774_ (.A1(_0808_),
    .A2(_0851_),
    .A3(_0838_),
    .B(_0849_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1775_ (.A1(_0850_),
    .A2(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1776_ (.A1(_0776_),
    .A2(_0807_),
    .A3(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1777_ (.A1(_0772_),
    .A2(_0854_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1778_ (.I(_0855_),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1779_ (.A1(_0577_),
    .A2(_0803_),
    .A3(_0765_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1780_ (.I(_0751_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1781_ (.A1(_0799_),
    .A2(_0856_),
    .B(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1782_ (.I(_0612_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1783_ (.I(_0721_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1784_ (.A1(_0860_),
    .A2(_0742_),
    .B(_0674_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1785_ (.A1(_0700_),
    .A2(_0731_),
    .A3(_0861_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1786_ (.I(_0547_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1787_ (.A1(_0761_),
    .A2(_0863_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1788_ (.A1(_0795_),
    .A2(_0742_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1789_ (.I(_0573_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1790_ (.A1(_0694_),
    .A2(_0864_),
    .B(_0865_),
    .C(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1791_ (.A1(_0664_),
    .A2(_0333_),
    .B(_0572_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1792_ (.A1(_0783_),
    .A2(_0619_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1793_ (.A1(_0868_),
    .A2(_0869_),
    .B(_0631_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1794_ (.A1(_0859_),
    .A2(_0862_),
    .A3(_0867_),
    .B1(_0870_),
    .B2(_0723_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1795_ (.A1(_0858_),
    .A2(_0871_),
    .B(_0531_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1796_ (.A1(_0858_),
    .A2(_0871_),
    .B(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1797_ (.A1(_0814_),
    .A2(_0819_),
    .A3(_0824_),
    .B(_0520_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1798_ (.I(_0874_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1799_ (.I(_0859_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1800_ (.I(_0817_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1801_ (.I(_0673_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1802_ (.A1(_0694_),
    .A2(_0785_),
    .B1(_0877_),
    .B2(_0878_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1803_ (.I0(_0688_),
    .I1(_0879_),
    .S(_0700_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1804_ (.A1(_0761_),
    .A2(_0860_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1805_ (.A1(_0860_),
    .A2(_0603_),
    .B(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1806_ (.I(_0809_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1807_ (.I(_0789_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1808_ (.I(_0884_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1809_ (.I(_0599_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1810_ (.I(_0794_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1811_ (.A1(_0809_),
    .A2(_0887_),
    .B(_0884_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1812_ (.A1(_0883_),
    .A2(_0885_),
    .B1(_0886_),
    .B2(_0888_),
    .C(_0728_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1813_ (.A1(_0876_),
    .A2(_0880_),
    .B1(_0882_),
    .B2(_0759_),
    .C(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1814_ (.A1(_0835_),
    .A2(_0875_),
    .B(_0890_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1815_ (.A1(_0835_),
    .A2(_0874_),
    .A3(_0890_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1816_ (.A1(_0833_),
    .A2(_0891_),
    .A3(_0892_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1817_ (.A1(_0634_),
    .A2(_0683_),
    .A3(_0746_),
    .A4(_0848_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1818_ (.A1(_0523_),
    .A2(_0894_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1819_ (.I(_0753_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1820_ (.A1(_0756_),
    .A2(_0817_),
    .B(_0884_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1821_ (.A1(_0676_),
    .A2(_0543_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1822_ (.A1(_0898_),
    .A2(_0743_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1823_ (.A1(_0690_),
    .A2(_0868_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1824_ (.A1(_0886_),
    .A2(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1825_ (.A1(_0720_),
    .A2(_0593_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1826_ (.A1(_0821_),
    .A2(_0901_),
    .B1(_0902_),
    .B2(_0809_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1827_ (.A1(_0896_),
    .A2(_0897_),
    .A3(_0899_),
    .B1(_0903_),
    .B2(_0859_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1828_ (.A1(_0895_),
    .A2(_0904_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1829_ (.A1(_0607_),
    .A2(_0832_),
    .A3(_0893_),
    .A4(_0905_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1830_ (.I(_0607_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1831_ (.A1(_0907_),
    .A2(_0851_),
    .A3(_0893_),
    .B(_0905_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1832_ (.A1(_0873_),
    .A2(_0906_),
    .A3(_0908_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1833_ (.I(_0906_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1834_ (.A1(_0910_),
    .A2(_0908_),
    .B(_0873_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1835_ (.A1(_0907_),
    .A2(_0851_),
    .A3(_0838_),
    .A4(_0849_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1836_ (.A1(_0807_),
    .A2(_0852_),
    .B(_0912_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1837_ (.A1(_0909_),
    .A2(_0911_),
    .A3(_0913_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1838_ (.A1(_0909_),
    .A2(_0911_),
    .B(_0913_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1839_ (.A1(_0914_),
    .A2(_0915_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1840_ (.A1(_0807_),
    .A2(_0853_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1841_ (.A1(_0776_),
    .A2(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1842_ (.A1(_0772_),
    .A2(_0854_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1843_ (.A1(_0918_),
    .A2(_0919_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1844_ (.A1(_0916_),
    .A2(_0920_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1845_ (.I(_0921_),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1846_ (.A1(_0873_),
    .A2(_0910_),
    .A3(_0908_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1847_ (.A1(_0836_),
    .A2(_0837_),
    .B(_0833_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1848_ (.A1(_0793_),
    .A2(_0603_),
    .B1(_0697_),
    .B2(_0739_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1849_ (.I(_0581_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1850_ (.A1(_0676_),
    .A2(_0925_),
    .B(_0568_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1851_ (.A1(_0705_),
    .A2(_0612_),
    .A3(_0924_),
    .A4(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1852_ (.A1(_0810_),
    .A2(_0654_),
    .B(_0896_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1853_ (.I(_0680_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1854_ (.A1(_0929_),
    .A2(_0926_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1855_ (.A1(_0927_),
    .A2(_0928_),
    .A3(_0930_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1856_ (.I0(_0521_),
    .I1(_0874_),
    .S(_0931_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1857_ (.A1(_0830_),
    .A2(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1858_ (.A1(_0609_),
    .A2(_0923_),
    .A3(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1859_ (.I(_0739_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1860_ (.A1(_0935_),
    .A2(_0613_),
    .B(_0865_),
    .C(_0705_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1861_ (.I(_0755_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1862_ (.A1(_0866_),
    .A2(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1863_ (.A1(_0884_),
    .A2(_0592_),
    .B(_0644_),
    .C(_0937_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1864_ (.A1(_0859_),
    .A2(_0936_),
    .A3(_0938_),
    .B1(_0598_),
    .B2(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1865_ (.A1(_0894_),
    .A2(_0904_),
    .B(_0522_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1866_ (.A1(_0940_),
    .A2(_0941_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1867_ (.I(_0896_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1868_ (.I(_0440_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1869_ (.A1(_0694_),
    .A2(_0756_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1870_ (.A1(_0944_),
    .A2(_0945_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1871_ (.A1(_0943_),
    .A2(_0946_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1872_ (.I(_0704_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1873_ (.A1(_0613_),
    .A2(_0588_),
    .B(_0866_),
    .C(_0935_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1874_ (.A1(_0925_),
    .A2(_0784_),
    .B1(_0594_),
    .B2(_0878_),
    .C(_0700_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1875_ (.A1(_0948_),
    .A2(_0949_),
    .A3(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1876_ (.A1(_0947_),
    .A2(_0951_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1877_ (.A1(_0782_),
    .A2(_0788_),
    .A3(_0798_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1878_ (.A1(_0953_),
    .A2(_0804_),
    .A3(_0871_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1879_ (.A1(_0751_),
    .A2(_0952_),
    .A3(_0954_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1880_ (.A1(_0857_),
    .A2(_0954_),
    .B(_0952_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1881_ (.A1(_0530_),
    .A2(_0955_),
    .A3(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _1882_ (.A1(_0934_),
    .A2(_0942_),
    .A3(_0957_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1883_ (.A1(_0910_),
    .A2(_0922_),
    .B(_0958_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1884_ (.A1(_0910_),
    .A2(_0922_),
    .A3(_0958_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1885_ (.A1(_0959_),
    .A2(_0960_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1886_ (.A1(_0909_),
    .A2(_0911_),
    .A3(_0913_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1887_ (.A1(_0915_),
    .A2(_0920_),
    .B(_0962_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1888_ (.A1(_0961_),
    .A2(_0963_),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1889_ (.I(_0964_),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1890_ (.A1(_0927_),
    .A2(_0928_),
    .A3(_0930_),
    .B(_0641_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1891_ (.A1(_0793_),
    .A2(_0795_),
    .A3(_0794_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1892_ (.A1(_0866_),
    .A2(_0693_),
    .A3(_0817_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1893_ (.A1(_0966_),
    .A2(_0967_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1894_ (.A1(_0863_),
    .A2(_0604_),
    .B(_0896_),
    .C(_0626_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1895_ (.A1(_0863_),
    .A2(_0674_),
    .B(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1896_ (.A1(_0935_),
    .A2(_0816_),
    .A3(_0929_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1897_ (.A1(_0876_),
    .A2(_0968_),
    .B(_0970_),
    .C(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1898_ (.A1(_0875_),
    .A2(_0965_),
    .B(_0972_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1899_ (.A1(_0875_),
    .A2(_0965_),
    .A3(_0972_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1900_ (.A1(_0833_),
    .A2(_0973_),
    .A3(_0974_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1901_ (.A1(_0894_),
    .A2(_0904_),
    .A3(_0940_),
    .B(_0522_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1902_ (.I(_0976_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1903_ (.A1(_0674_),
    .A2(_0779_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1904_ (.A1(_0701_),
    .A2(_0593_),
    .A3(_0978_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1905_ (.A1(_0948_),
    .A2(_0484_),
    .A3(_0979_),
    .B1(_0924_),
    .B2(_0943_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1906_ (.I0(_0977_),
    .I1(_0523_),
    .S(_0980_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1907_ (.A1(_0808_),
    .A2(_0832_),
    .A3(_0975_),
    .A4(_0981_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1908_ (.A1(_0808_),
    .A2(_0832_),
    .A3(_0975_),
    .B(_0981_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1909_ (.I(_0720_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1910_ (.I(_0984_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1911_ (.A1(_0883_),
    .A2(_0985_),
    .A3(_0691_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1912_ (.A1(_0743_),
    .A2(_0645_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1913_ (.A1(_0860_),
    .A2(_0878_),
    .B(_0877_),
    .C(_0984_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1914_ (.A1(_0987_),
    .A2(_0988_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1915_ (.A1(_0948_),
    .A2(_0986_),
    .A3(_0989_),
    .B1(_0944_),
    .B2(_0943_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1916_ (.A1(_0704_),
    .A2(_0949_),
    .A3(_0950_),
    .B1(_0943_),
    .B2(_0946_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1917_ (.A1(_0953_),
    .A2(_0804_),
    .A3(_0871_),
    .A4(_0991_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1918_ (.A1(_0751_),
    .A2(_0992_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1919_ (.A1(_0990_),
    .A2(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1920_ (.A1(_0531_),
    .A2(_0982_),
    .A3(_0983_),
    .A4(_0994_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1921_ (.A1(_0982_),
    .A2(_0983_),
    .B1(_0994_),
    .B2(_0532_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1922_ (.A1(_0995_),
    .A2(_0996_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1923_ (.A1(_0907_),
    .A2(_0851_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1924_ (.A1(_0998_),
    .A2(_0933_),
    .B(_0942_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1925_ (.A1(_0998_),
    .A2(_0933_),
    .A3(_0942_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1926_ (.A1(_0999_),
    .A2(_0957_),
    .B(_1000_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1927_ (.A1(_0997_),
    .A2(_1001_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1928_ (.A1(_0918_),
    .A2(_0919_),
    .B(_0916_),
    .C(_0961_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1929_ (.A1(_0962_),
    .A2(_0959_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1930_ (.A1(_0960_),
    .A2(_1004_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1931_ (.A1(_1003_),
    .A2(_1005_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1932_ (.A1(_1002_),
    .A2(_1006_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1933_ (.I(_1007_),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1934_ (.A1(_0609_),
    .A2(_0923_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1935_ (.I(_1008_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1936_ (.A1(_1009_),
    .A2(_0975_),
    .A3(_0981_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1937_ (.A1(_0874_),
    .A2(_0965_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1938_ (.A1(_0816_),
    .A2(_0698_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1939_ (.A1(_0885_),
    .A2(_0791_),
    .B(_1012_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1940_ (.I(_0900_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1941_ (.A1(_0811_),
    .A2(_1014_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1942_ (.A1(_0761_),
    .A2(_0935_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1943_ (.A1(_0704_),
    .A2(_0812_),
    .A3(_1016_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1944_ (.A1(_0759_),
    .A2(_1013_),
    .B1(_1015_),
    .B2(_0787_),
    .C(_1017_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1945_ (.I0(\p_shaping_Q.p_shaping_I.bit_in_1 ),
    .I1(_1011_),
    .S(_1018_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1946_ (.A1(_0734_),
    .A2(_0735_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1947_ (.A1(_0718_),
    .A2(_1020_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1948_ (.A1(_0834_),
    .A2(_1019_),
    .B(_1021_),
    .C(_0640_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1949_ (.A1(_0878_),
    .A2(_0898_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1950_ (.A1(_0944_),
    .A2(_1023_),
    .B1(_0886_),
    .B2(_0885_),
    .C(_0812_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1951_ (.A1(_0876_),
    .A2(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1952_ (.A1(_0719_),
    .A2(_0502_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1953_ (.A1(_0948_),
    .A2(_0877_),
    .B(_1025_),
    .C(_1026_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1954_ (.A1(_0976_),
    .A2(_1027_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1955_ (.I(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1956_ (.I(_0993_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1957_ (.I(_0719_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1958_ (.I(_0985_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1959_ (.A1(_0985_),
    .A2(_0886_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _1960_ (.A1(_1032_),
    .A2(_0476_),
    .A3(_0731_),
    .B1(_0869_),
    .B2(_1014_),
    .B3(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1961_ (.A1(_1031_),
    .A2(_1034_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1962_ (.A1(_0857_),
    .A2(_0992_),
    .A3(_1035_),
    .B(_0530_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1963_ (.A1(_1030_),
    .A2(_1035_),
    .B(_1036_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1964_ (.A1(_1022_),
    .A2(_1029_),
    .A3(_1037_),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1965_ (.A1(_1010_),
    .A2(_0995_),
    .B(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1966_ (.A1(_1010_),
    .A2(_0995_),
    .A3(_1038_),
    .Z(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1967_ (.A1(_1039_),
    .A2(_1040_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1968_ (.I(_0997_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1969_ (.A1(_1042_),
    .A2(_1001_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1970_ (.A1(_1002_),
    .A2(_1006_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1971_ (.A1(_1043_),
    .A2(_1044_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1972_ (.A1(_1041_),
    .A2(_1045_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1973_ (.I(_1046_),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1974_ (.A1(_0703_),
    .A2(_0925_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1975_ (.A1(_0695_),
    .A2(_0677_),
    .B(_0843_),
    .C(_1047_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1976_ (.A1(_0728_),
    .A2(_1048_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1977_ (.A1(_0883_),
    .A2(_0887_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1978_ (.A1(_0810_),
    .A2(_0791_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1979_ (.A1(_1050_),
    .A2(_0698_),
    .B(_1051_),
    .C(_0984_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1980_ (.A1(_0984_),
    .A2(_0688_),
    .B1(_0816_),
    .B2(_0698_),
    .C(_1051_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1981_ (.A1(_1049_),
    .A2(_1052_),
    .B1(_1053_),
    .B2(_0719_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1982_ (.A1(_1011_),
    .A2(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1983_ (.A1(_0521_),
    .A2(_1054_),
    .B(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1984_ (.A1(_0834_),
    .A2(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1985_ (.A1(_1008_),
    .A2(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1986_ (.A1(_0756_),
    .A2(_0877_),
    .B(_0695_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1987_ (.A1(_0985_),
    .A2(_0553_),
    .A3(_1059_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1988_ (.A1(_0839_),
    .A2(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1989_ (.A1(_0504_),
    .A2(_1061_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1990_ (.A1(_0523_),
    .A2(_0504_),
    .B1(_0977_),
    .B2(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1991_ (.A1(_1058_),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1992_ (.I(_0857_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1993_ (.A1(_0695_),
    .A2(_0627_),
    .B(_0938_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1994_ (.A1(_0568_),
    .A2(_1014_),
    .B(_1032_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1995_ (.A1(_1031_),
    .A2(_1066_),
    .A3(_1067_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1996_ (.A1(_1065_),
    .A2(_0880_),
    .B(_1030_),
    .C(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1997_ (.A1(_1065_),
    .A2(_1068_),
    .B(_1069_),
    .C(_0532_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1998_ (.A1(_1064_),
    .A2(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1999_ (.A1(_1022_),
    .A2(_1029_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2000_ (.A1(_1022_),
    .A2(_1029_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2001_ (.A1(_1072_),
    .A2(_1037_),
    .B(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2002_ (.A1(_1071_),
    .A2(_1074_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2003_ (.A1(_1002_),
    .A2(_1041_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2004_ (.A1(_1003_),
    .A2(_1005_),
    .B(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2005_ (.I(_1039_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2006_ (.A1(_1043_),
    .A2(_1040_),
    .B(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2007_ (.A1(_1077_),
    .A2(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2008_ (.A1(_1075_),
    .A2(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2009_ (.I(_1081_),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2010_ (.A1(_1058_),
    .A2(_1063_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2011_ (.A1(_1064_),
    .A2(_1070_),
    .B(_1082_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2012_ (.I(_0876_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2013_ (.A1(_0783_),
    .A2(_0784_),
    .B(_0925_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2014_ (.A1(_1032_),
    .A2(_0588_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2015_ (.A1(_1085_),
    .A2(_1086_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2016_ (.A1(_1031_),
    .A2(_0569_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2017_ (.A1(_1084_),
    .A2(_1060_),
    .B1(_1087_),
    .B2(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2018_ (.A1(_0875_),
    .A2(_0965_),
    .B(_1089_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2019_ (.A1(\p_shaping_Q.p_shaping_I.bit_in_1 ),
    .A2(_1089_),
    .B(_1090_),
    .C(_0834_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2020_ (.A1(_1009_),
    .A2(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2021_ (.A1(_1084_),
    .A2(_0944_),
    .A3(_0691_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2022_ (.A1(_1026_),
    .A2(_0633_),
    .A3(_1093_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2023_ (.A1(_0977_),
    .A2(_1094_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2024_ (.A1(_0839_),
    .A2(_1094_),
    .B(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2025_ (.A1(_1092_),
    .A2(_1096_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2026_ (.I(_0532_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2027_ (.I(_1032_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2028_ (.A1(_1099_),
    .A2(_1014_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2029_ (.A1(_1031_),
    .A2(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2030_ (.A1(_0887_),
    .A2(_0692_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2031_ (.A1(_0588_),
    .A2(_1102_),
    .B(_0937_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2032_ (.A1(_1099_),
    .A2(_1103_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2033_ (.A1(_1101_),
    .A2(_1104_),
    .B(_1030_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2034_ (.A1(_1065_),
    .A2(_1101_),
    .A3(_1104_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2035_ (.A1(_1098_),
    .A2(_1105_),
    .A3(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2036_ (.A1(_1097_),
    .A2(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2037_ (.A1(_1071_),
    .A2(_1074_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2038_ (.A1(_1077_),
    .A2(_1079_),
    .B(_1075_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2039_ (.A1(_1109_),
    .A2(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2040_ (.A1(_1083_),
    .A2(_1108_),
    .A3(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2041_ (.I(_1112_),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2042_ (.A1(_0830_),
    .A2(_1011_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2043_ (.A1(_1021_),
    .A2(_1113_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2044_ (.A1(_0937_),
    .A2(_1023_),
    .B(_0701_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2045_ (.A1(_0929_),
    .A2(_0946_),
    .B1(_1115_),
    .B2(_1084_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2046_ (.A1(_1114_),
    .A2(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2047_ (.A1(_0640_),
    .A2(_1117_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2048_ (.A1(_0503_),
    .A2(_0977_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2049_ (.A1(_0839_),
    .A2(_0503_),
    .B(_0633_),
    .C(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2050_ (.A1(_1118_),
    .A2(_1120_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2051_ (.I(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2052_ (.A1(_1099_),
    .A2(_0688_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2053_ (.A1(_1101_),
    .A2(_1123_),
    .B(_1030_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2054_ (.A1(_1065_),
    .A2(_1101_),
    .A3(_1123_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2055_ (.A1(_1098_),
    .A2(_1124_),
    .A3(_1125_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2056_ (.I(_1126_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2057_ (.A1(_1122_),
    .A2(_1127_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2058_ (.A1(_1098_),
    .A2(_1097_),
    .A3(_1105_),
    .A4(_1106_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2059_ (.A1(_1009_),
    .A2(_1091_),
    .A3(_1096_),
    .B(_1129_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2060_ (.A1(_1128_),
    .A2(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2061_ (.A1(_1083_),
    .A2(_1108_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2062_ (.A1(_1071_),
    .A2(_1074_),
    .B(_1132_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2063_ (.A1(_1083_),
    .A2(_1108_),
    .B1(_1133_),
    .B2(_1110_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2064_ (.A1(_1131_),
    .A2(_1134_),
    .Z(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2065_ (.I(_1135_),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2066_ (.A1(_1118_),
    .A2(_1120_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2067_ (.A1(_1122_),
    .A2(_1127_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2068_ (.A1(_0929_),
    .A2(_0945_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2069_ (.A1(_0574_),
    .A2(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2070_ (.A1(_0521_),
    .A2(_1139_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2071_ (.A1(_1011_),
    .A2(_1139_),
    .B(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2072_ (.A1(_0830_),
    .A2(_1141_),
    .B(_1009_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2073_ (.A1(_1120_),
    .A2(_1126_),
    .A3(_1142_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2074_ (.A1(_1136_),
    .A2(_1137_),
    .B(_1143_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2075_ (.A1(_1136_),
    .A2(_1137_),
    .A3(_1143_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2076_ (.A1(_1144_),
    .A2(_1145_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2077_ (.A1(_1128_),
    .A2(_1130_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2078_ (.A1(_1131_),
    .A2(_1134_),
    .B(_1147_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2079_ (.A1(_1146_),
    .A2(_1148_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2080_ (.I(_1149_),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2081_ (.A1(_1131_),
    .A2(_1134_),
    .A3(_1146_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2082_ (.A1(_1136_),
    .A2(_1137_),
    .A3(_1143_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2083_ (.A1(_1147_),
    .A2(_1151_),
    .B(_1144_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2084_ (.A1(_1127_),
    .A2(_1142_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2085_ (.A1(_1127_),
    .A2(_1142_),
    .B(_1120_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2086_ (.A1(_1153_),
    .A2(_1154_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2087_ (.A1(_1150_),
    .A2(_1152_),
    .A3(_1155_),
    .B1(_1114_),
    .B2(_0907_),
    .ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2088_ (.A1(_0639_),
    .A2(_0712_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2089_ (.I(_1156_),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2090_ (.A1(net33),
    .A2(net32),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2091_ (.I(_1157_),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2092_ (.I(_1158_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2093_ (.I(_0226_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2094_ (.I(_1258_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2095_ (.I(_0140_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2096_ (.A1(_1161_),
    .A2(_1162_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2097_ (.A1(_1160_),
    .A2(_1163_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2098_ (.I(_0215_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2099_ (.I(_1258_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2100_ (.I(_1166_),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2101_ (.I(_1167_),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2102_ (.I(_1162_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2103_ (.A1(_1165_),
    .A2(_1168_),
    .B(_1169_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2104_ (.I(_1181_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2105_ (.I(_1172_),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2106_ (.I(_1173_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2107_ (.I(net32),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2108_ (.A1(_0129_),
    .A2(_1175_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2109_ (.I(_1176_),
    .Z(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2110_ (.I(_0096_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2111_ (.A1(_1174_),
    .A2(_1177_),
    .B(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2112_ (.I(_0107_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2113_ (.I(_1180_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2114_ (.A1(_1159_),
    .A2(_1164_),
    .B1(_1171_),
    .B2(_1179_),
    .C(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2115_ (.A1(_1175_),
    .A2(_1192_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2116_ (.A1(_0096_),
    .A2(_1184_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2117_ (.I(_1185_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2118_ (.I(_0226_),
    .Z(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2119_ (.I(_1187_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2120_ (.A1(_1236_),
    .A2(_1181_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2121_ (.I(_1189_),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2122_ (.A1(_0215_),
    .A2(_1161_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2123_ (.A1(_1188_),
    .A2(_1190_),
    .B(_1191_),
    .C(_1334_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2124_ (.A1(_0107_),
    .A2(_1323_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2125_ (.I(_1194_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2126_ (.A1(_1186_),
    .A2(_1193_),
    .B(_1195_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2127_ (.A1(_0054_),
    .A2(_1175_),
    .A3(_0140_),
    .Z(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2128_ (.A1(_0237_),
    .A2(_1197_),
    .B(_0065_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2129_ (.A1(_0043_),
    .A2(_1198_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2130_ (.I(_1199_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2131_ (.I(_1170_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2132_ (.I(_1201_),
    .Z(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2133_ (.A1(_0054_),
    .A2(_1279_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2134_ (.I(_0054_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2135_ (.I(_1205_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2136_ (.I(_1173_),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2137_ (.A1(_1206_),
    .A2(_1202_),
    .A3(_1207_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2138_ (.A1(_1202_),
    .A2(_1204_),
    .B(_1208_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2139_ (.A1(_1183_),
    .A2(_1196_),
    .B1(_1200_),
    .B2(_1209_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2140_ (.A1(\p_shaping_I.p_shaping_I.counter[1] ),
    .A2(\p_shaping_I.p_shaping_I.counter[0] ),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2141_ (.I(_1211_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2142_ (.A1(_1210_),
    .A2(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2143_ (.I(_0085_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2144_ (.I(_1192_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2145_ (.A1(_1216_),
    .A2(_1158_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2146_ (.I(_0226_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2147_ (.A1(_1173_),
    .A2(_1176_),
    .B(_1218_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2148_ (.I(_0129_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2149_ (.I(_1214_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2150_ (.A1(_1220_),
    .A2(_1221_),
    .A3(_1216_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2151_ (.A1(_1217_),
    .A2(_1219_),
    .B(_1180_),
    .C(_1222_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2152_ (.A1(_1215_),
    .A2(_1223_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2153_ (.I(_1221_),
    .Z(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2154_ (.A1(_1247_),
    .A2(_1268_),
    .B(_1192_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2155_ (.I(_1227_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2156_ (.I(_1180_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2157_ (.A1(_1226_),
    .A2(_1228_),
    .B(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2158_ (.I(_1175_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2159_ (.A1(_1220_),
    .A2(_1231_),
    .B(_1173_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2160_ (.I(_1166_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2161_ (.A1(_1233_),
    .A2(_1216_),
    .B(_1160_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2162_ (.I(_1189_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2163_ (.A1(_1233_),
    .A2(_1216_),
    .B(_1235_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2164_ (.A1(_0096_),
    .A2(_1176_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2165_ (.I(_0118_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2166_ (.A1(_1232_),
    .A2(_1234_),
    .B1(_1237_),
    .B2(_1238_),
    .C(_1239_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2167_ (.A1(_1230_),
    .A2(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2168_ (.A1(_1224_),
    .A2(_1241_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2169_ (.I(\p_shaping_I.p_shaping_I.counter[1] ),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2170_ (.I(_1160_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2171_ (.I(_1191_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2172_ (.A1(_1231_),
    .A2(_0237_),
    .A3(_1235_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2173_ (.A1(_1178_),
    .A2(_1227_),
    .B(_1246_),
    .C(_1180_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2174_ (.I(_1279_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2175_ (.A1(_1225_),
    .A2(_1249_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2176_ (.A1(_1218_),
    .A2(_1158_),
    .B(_0043_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2177_ (.I(_1162_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2178_ (.I(_0065_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2179_ (.A1(_1165_),
    .A2(_1250_),
    .B1(_1251_),
    .B2(_1252_),
    .C(_1253_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2180_ (.I(_1170_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2181_ (.A1(_1255_),
    .A2(_1253_),
    .B(_1239_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2182_ (.A1(_1244_),
    .A2(_1245_),
    .B1(_1248_),
    .B2(_1254_),
    .C(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2183_ (.I(_1257_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2184_ (.A1(_1243_),
    .A2(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2185_ (.A1(_1242_),
    .A2(_1260_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2186_ (.A1(_1213_),
    .A2(_1261_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2187_ (.I(_1262_),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2188_ (.A1(_1242_),
    .A2(_1260_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2189_ (.A1(_1213_),
    .A2(_1261_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2190_ (.I(_0074_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2191_ (.I(_1163_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2192_ (.I(_1221_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2193_ (.A1(_1206_),
    .A2(_1266_),
    .B(_1267_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2194_ (.A1(_1190_),
    .A2(_1266_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2195_ (.I(_1312_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2196_ (.A1(_1269_),
    .A2(_1270_),
    .B(_1271_),
    .C(_1217_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2197_ (.I(_1239_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2198_ (.A1(_1265_),
    .A2(_1272_),
    .B(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2199_ (.I(_1247_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2200_ (.I(_1172_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2201_ (.A1(_1275_),
    .A2(_1168_),
    .A3(_1276_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2202_ (.A1(_1161_),
    .A2(_0237_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2203_ (.A1(_1278_),
    .A2(_1204_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2204_ (.I(_1312_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2205_ (.A1(_1186_),
    .A2(_1277_),
    .B(_1280_),
    .C(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2206_ (.A1(_1275_),
    .A2(_1276_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2207_ (.A1(_1187_),
    .A2(_1290_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2208_ (.A1(_1267_),
    .A2(_1283_),
    .B(_1284_),
    .C(_1229_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2209_ (.A1(_1273_),
    .A2(_1282_),
    .A3(_1285_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2210_ (.A1(_1274_),
    .A2(_1286_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2211_ (.A1(_0511_),
    .A2(_1210_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2212_ (.A1(_1287_),
    .A2(_1288_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2213_ (.A1(_1211_),
    .A2(_1289_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2214_ (.I(\p_shaping_I.p_shaping_I.counter[1] ),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2215_ (.I(\p_shaping_I.p_shaping_I.bit_in_2 ),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2216_ (.A1(_0107_),
    .A2(_0118_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2217_ (.I(_1294_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2218_ (.A1(_1255_),
    .A2(_1159_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2219_ (.A1(_1205_),
    .A2(_1167_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2220_ (.A1(_1247_),
    .A2(_1161_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2221_ (.A1(_1203_),
    .A2(_1298_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2222_ (.A1(_1201_),
    .A2(_1169_),
    .A3(_1297_),
    .B(_1299_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2223_ (.A1(_1233_),
    .A2(_0248_),
    .B(_1235_),
    .C(_1187_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2224_ (.A1(_1221_),
    .A2(_0248_),
    .A3(_1158_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2225_ (.A1(_1302_),
    .A2(_1303_),
    .B(_1194_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2226_ (.A1(_1295_),
    .A2(_1296_),
    .B1(_1300_),
    .B2(_1199_),
    .C(_1304_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2227_ (.A1(_1293_),
    .A2(_1259_),
    .A3(_1305_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2228_ (.I(\p_shaping_I.p_shaping_I.bit_in_2 ),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2229_ (.A1(_1307_),
    .A2(_1259_),
    .B(_1305_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2230_ (.A1(_1292_),
    .A2(_1306_),
    .A3(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2231_ (.A1(_1225_),
    .A2(_1227_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2232_ (.A1(_1310_),
    .A2(_1302_),
    .A3(_1303_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2233_ (.A1(_1312_),
    .A2(_1323_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2234_ (.A1(_1167_),
    .A2(_1172_),
    .B(_0215_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2235_ (.A1(_1255_),
    .A2(_1313_),
    .A3(_1314_),
    .B(_0161_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2236_ (.A1(_1205_),
    .A2(_1233_),
    .B(_1187_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2237_ (.A1(_1195_),
    .A2(_1284_),
    .A3(_1316_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2238_ (.A1(_1345_),
    .A2(_1311_),
    .B(_1315_),
    .C(_1317_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2239_ (.A1(_1215_),
    .A2(_1223_),
    .B1(_1230_),
    .B2(_1240_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2240_ (.A1(\p_shaping_I.p_shaping_I.bit_in ),
    .A2(_1319_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2241_ (.A1(_1318_),
    .A2(_1320_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2242_ (.A1(_1291_),
    .A2(_1309_),
    .A3(_1321_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2243_ (.A1(_1263_),
    .A2(_1264_),
    .B(_1322_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2244_ (.A1(_1309_),
    .A2(_1321_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2245_ (.A1(_1309_),
    .A2(_1321_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2246_ (.A1(_1291_),
    .A2(_1325_),
    .B(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2247_ (.I(_1211_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2248_ (.I(_1328_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2249_ (.A1(_0508_),
    .A2(_0517_),
    .Z(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2250_ (.A1(_0280_),
    .A2(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2251_ (.I(_1195_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2252_ (.A1(_1236_),
    .A2(_1258_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2253_ (.A1(_1169_),
    .A2(_1333_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2254_ (.I(_1172_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2255_ (.A1(_0194_),
    .A2(_1336_),
    .B(_1218_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2256_ (.I(_1167_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2257_ (.A1(_1338_),
    .A2(_1174_),
    .B(_1178_),
    .C(_1165_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2258_ (.A1(_1335_),
    .A2(_1337_),
    .B(_1339_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2259_ (.I(_1268_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2260_ (.A1(_1341_),
    .A2(_1188_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2261_ (.A1(_1275_),
    .A2(_1249_),
    .B(_0194_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2262_ (.A1(_1226_),
    .A2(_1190_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2263_ (.A1(_1342_),
    .A2(_1343_),
    .B(_1295_),
    .C(_1344_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2264_ (.A1(_1255_),
    .A2(_1174_),
    .A3(_1333_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2265_ (.A1(_1341_),
    .A2(_0258_),
    .B(_1229_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2266_ (.I(_0043_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2267_ (.A1(_0023_),
    .A2(_0024_),
    .A3(_1339_),
    .B(_0025_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2268_ (.A1(_1332_),
    .A2(_1340_),
    .B(_0022_),
    .C(_0026_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2269_ (.A1(_1183_),
    .A2(_1196_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2270_ (.A1(_1200_),
    .A2(_1209_),
    .B1(_1274_),
    .B2(_1286_),
    .C(_0028_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2271_ (.A1(_0511_),
    .A2(_0029_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2272_ (.A1(_1331_),
    .A2(_0027_),
    .A3(_0030_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2273_ (.A1(_1329_),
    .A2(_0031_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2274_ (.I(_1334_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2275_ (.A1(_1226_),
    .A2(_1232_),
    .B(_1185_),
    .C(_1253_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2276_ (.A1(_1205_),
    .A2(_1231_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2277_ (.A1(_1249_),
    .A2(_0036_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2278_ (.A1(_1201_),
    .A2(_1336_),
    .A3(_1177_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2279_ (.A1(_1278_),
    .A2(_1294_),
    .A3(_0037_),
    .A4(_0038_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2280_ (.A1(_1220_),
    .A2(_1231_),
    .B(_0248_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2281_ (.A1(_0065_),
    .A2(_0118_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2282_ (.A1(_1164_),
    .A2(_0040_),
    .B1(_1238_),
    .B2(_1163_),
    .C(_0041_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2283_ (.A1(_0034_),
    .A2(_0035_),
    .B(_0039_),
    .C(_0042_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2284_ (.A1(_1259_),
    .A2(_1305_),
    .B(_1293_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2285_ (.A1(_0044_),
    .A2(_0045_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2286_ (.A1(_1319_),
    .A2(_1318_),
    .B(\p_shaping_I.p_shaping_I.bit_in ),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2287_ (.I(_1220_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2288_ (.A1(_0048_),
    .A2(_1184_),
    .B(_1218_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2289_ (.A1(_1336_),
    .A2(_1177_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2290_ (.A1(_0049_),
    .A2(_0050_),
    .B(_1284_),
    .C(_0025_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2291_ (.A1(_1341_),
    .A2(_1235_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2292_ (.A1(_1267_),
    .A2(_1297_),
    .B1(_0052_),
    .B2(_1278_),
    .C(_1334_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2293_ (.A1(_0051_),
    .A2(_0053_),
    .B(_1182_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2294_ (.I(_1333_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2295_ (.A1(_1174_),
    .A2(_0056_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2296_ (.A1(_1295_),
    .A2(_0057_),
    .A3(_1219_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2297_ (.A1(_0055_),
    .A2(_0058_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2298_ (.A1(_0047_),
    .A2(_0059_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2299_ (.A1(_1243_),
    .A2(_0046_),
    .A3(_0060_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2300_ (.I(_1243_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2301_ (.A1(_0062_),
    .A2(_0046_),
    .B(_0060_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2302_ (.A1(_0061_),
    .A2(_0063_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2303_ (.A1(_1327_),
    .A2(_0033_),
    .A3(_0064_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2304_ (.A1(_1324_),
    .A2(_0066_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2305_ (.I(_0067_),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2306_ (.A1(_1329_),
    .A2(_0031_),
    .A3(_0061_),
    .A4(_0063_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2307_ (.I(_1329_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2308_ (.A1(_0021_),
    .A2(_0031_),
    .B1(_0061_),
    .B2(_0063_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2309_ (.A1(_1327_),
    .A2(_0068_),
    .A3(_0069_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2310_ (.A1(_1324_),
    .A2(_0066_),
    .B(_0070_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2311_ (.A1(_0062_),
    .A2(_0046_),
    .A3(_0060_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2312_ (.A1(_0072_),
    .A2(_0068_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2313_ (.I(_0027_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2314_ (.A1(_1202_),
    .A2(_0057_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2315_ (.A1(_0076_),
    .A2(_1270_),
    .B(_1199_),
    .C(_1222_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2316_ (.A1(_1244_),
    .A2(_1266_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2317_ (.I(_1281_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2318_ (.A1(_1246_),
    .A2(_0078_),
    .B(_0079_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2319_ (.A1(_1206_),
    .A2(_1207_),
    .B(_1281_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2320_ (.I(_1335_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2321_ (.A1(_1222_),
    .A2(_0081_),
    .A3(_0082_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2322_ (.A1(_0034_),
    .A2(_0080_),
    .A3(_0083_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2323_ (.A1(_0077_),
    .A2(_0084_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2324_ (.I(\p_shaping_I.p_shaping_I.bit_in_1 ),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2325_ (.A1(_0075_),
    .A2(_0029_),
    .B(_0086_),
    .C(_0087_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2326_ (.I(_1169_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2327_ (.A1(_0089_),
    .A2(_1245_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2328_ (.A1(_1207_),
    .A2(_0056_),
    .B(_1271_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2329_ (.A1(_0049_),
    .A2(_0090_),
    .B(_0091_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2330_ (.A1(_0074_),
    .A2(_0092_),
    .B(_0034_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2331_ (.I(_0025_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2332_ (.A1(_0094_),
    .A2(_1282_),
    .A3(_1285_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2333_ (.A1(_0093_),
    .A2(_0095_),
    .B(_1210_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2334_ (.A1(_0077_),
    .A2(_0084_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2335_ (.A1(_0087_),
    .A2(_0075_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2336_ (.A1(_0512_),
    .A2(_0097_),
    .B(_0098_),
    .C(_0099_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2337_ (.A1(_0291_),
    .A2(_1330_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2338_ (.I(_0101_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2339_ (.A1(_0088_),
    .A2(_0100_),
    .B(_0102_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2340_ (.A1(_0101_),
    .A2(_0088_),
    .A3(_0100_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2341_ (.A1(_1329_),
    .A2(_0103_),
    .A3(_0104_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2342_ (.A1(_1257_),
    .A2(_1305_),
    .A3(_0044_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2343_ (.I(_0106_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2344_ (.I(_1345_),
    .Z(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2345_ (.A1(_1160_),
    .A2(_1314_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2346_ (.A1(_1162_),
    .A2(_1157_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2347_ (.A1(_1168_),
    .A2(_1249_),
    .B(_0111_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2348_ (.A1(_0110_),
    .A2(_0112_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2349_ (.A1(_1217_),
    .A2(_1219_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2350_ (.I(_1190_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2351_ (.A1(_0114_),
    .A2(_1237_),
    .B1(_1337_),
    .B2(_0115_),
    .C(_1195_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2352_ (.A1(_1341_),
    .A2(_1276_),
    .B(_1178_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2353_ (.A1(_0150_),
    .A2(_0117_),
    .B1(_1204_),
    .B2(_1164_),
    .C(_1294_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2354_ (.I(_0119_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2355_ (.A1(_0109_),
    .A2(_0113_),
    .B(_0116_),
    .C(_0120_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2356_ (.I(_0121_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2357_ (.A1(_1293_),
    .A2(_0108_),
    .B(_0122_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2358_ (.A1(\p_shaping_I.p_shaping_I.bit_in_2 ),
    .A2(_0121_),
    .A3(_0106_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2359_ (.A1(_1292_),
    .A2(_0123_),
    .A3(_0124_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2360_ (.I(_0269_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2361_ (.I(_1343_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2362_ (.A1(_1229_),
    .A2(_1239_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2363_ (.A1(_0040_),
    .A2(_1316_),
    .B1(_0127_),
    .B2(_1238_),
    .C(_0128_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2364_ (.A1(_0194_),
    .A2(_1276_),
    .B(_1201_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2365_ (.A1(_1245_),
    .A2(_0131_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2366_ (.A1(_1253_),
    .A2(_1197_),
    .A3(_1299_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2367_ (.A1(_1275_),
    .A2(_1168_),
    .B(_1336_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2368_ (.A1(_1226_),
    .A2(_0134_),
    .B(_1246_),
    .C(_1281_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2369_ (.A1(_0132_),
    .A2(_0133_),
    .B(_0025_),
    .C(_0135_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2370_ (.A1(_1273_),
    .A2(_0126_),
    .B(_0130_),
    .C(_0136_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2371_ (.A1(_1319_),
    .A2(_1318_),
    .A3(_0055_),
    .A4(_0058_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2372_ (.A1(_0509_),
    .A2(_0138_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2373_ (.A1(_0137_),
    .A2(_0139_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2374_ (.A1(_0125_),
    .A2(_0141_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2375_ (.A1(_0105_),
    .A2(_0142_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2376_ (.A1(_0073_),
    .A2(_0143_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2377_ (.A1(_0071_),
    .A2(_0144_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2378_ (.I(_0145_),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2379_ (.I(_0034_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2380_ (.A1(_0089_),
    .A2(_1298_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2381_ (.A1(_0081_),
    .A2(_0147_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2382_ (.A1(_0114_),
    .A2(_0148_),
    .B(_1198_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2383_ (.I(_1250_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2384_ (.A1(_0048_),
    .A2(_0151_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2385_ (.A1(_0048_),
    .A2(_0204_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2386_ (.I(_1295_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2387_ (.A1(_1278_),
    .A2(_1283_),
    .B(_0153_),
    .C(_0154_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2388_ (.A1(_0146_),
    .A2(_0149_),
    .B1(_0152_),
    .B2(_1332_),
    .C(_0155_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2389_ (.A1(_0075_),
    .A2(_0098_),
    .B(_0511_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2390_ (.A1(_0030_),
    .A2(_0157_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2391_ (.A1(_0156_),
    .A2(_0158_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2392_ (.A1(_1328_),
    .A2(_0103_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2393_ (.A1(_0102_),
    .A2(_0159_),
    .B(_0160_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2394_ (.A1(_0122_),
    .A2(_0108_),
    .B(_1293_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2395_ (.A1(_1267_),
    .A2(_0150_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2396_ (.I(_1337_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2397_ (.A1(_0164_),
    .A2(_0052_),
    .B1(_0082_),
    .B2(_0165_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2398_ (.A1(_1313_),
    .A2(_0166_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2399_ (.A1(_1165_),
    .A2(_1252_),
    .B(_1188_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2400_ (.A1(_1271_),
    .A2(_0168_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2401_ (.A1(_1273_),
    .A2(_1238_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2402_ (.A1(_1202_),
    .A2(_0057_),
    .A3(_0147_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2403_ (.I(_0128_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2404_ (.A1(_0173_),
    .A2(_0023_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2405_ (.A1(_0169_),
    .A2(_0170_),
    .B1(_0171_),
    .B2(_0174_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2406_ (.A1(_0167_),
    .A2(_0175_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2407_ (.A1(_0163_),
    .A2(_0176_),
    .B(_1243_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2408_ (.A1(_0163_),
    .A2(_0176_),
    .B(_0177_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2409_ (.A1(_0137_),
    .A2(_0138_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2410_ (.A1(_0508_),
    .A2(_0179_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2411_ (.I(_0094_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2412_ (.I(_1206_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2413_ (.A1(_0048_),
    .A2(_1252_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2414_ (.A1(_1188_),
    .A2(_1197_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2415_ (.A1(_0184_),
    .A2(_0185_),
    .B(_0078_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2416_ (.A1(_0182_),
    .A2(_0169_),
    .B1(_0186_),
    .B2(_0079_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2417_ (.A1(_1297_),
    .A2(_0117_),
    .B(_1299_),
    .C(_0050_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2418_ (.A1(_0109_),
    .A2(_0188_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2419_ (.A1(_0181_),
    .A2(_0187_),
    .B(_0189_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2420_ (.A1(_0180_),
    .A2(_0190_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2421_ (.A1(_0178_),
    .A2(_0191_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2422_ (.A1(_0162_),
    .A2(_0192_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2423_ (.A1(_0160_),
    .A2(_0104_),
    .A3(_0142_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2424_ (.A1(_0125_),
    .A2(_0141_),
    .B(_0195_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _2425_ (.A1(_0193_),
    .A2(_0196_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2426_ (.A1(_0073_),
    .A2(_0143_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2427_ (.A1(_0071_),
    .A2(_0144_),
    .B(_0198_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2428_ (.A1(_0197_),
    .A2(_0199_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2429_ (.I(_0200_),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2430_ (.A1(_0178_),
    .A2(_0191_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2431_ (.A1(_0162_),
    .A2(_0192_),
    .B(_0201_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2432_ (.I(_0102_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2433_ (.I(_1207_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2434_ (.A1(_0205_),
    .A2(_0153_),
    .B(_1316_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2435_ (.I(_1244_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2436_ (.A1(_0207_),
    .A2(_1343_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2437_ (.I(_1310_),
    .Z(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2438_ (.A1(_0131_),
    .A2(_0206_),
    .B1(_0208_),
    .B2(_0209_),
    .C(_1313_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2439_ (.A1(_1338_),
    .A2(_0151_),
    .B(_1280_),
    .C(_0173_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2440_ (.A1(_0041_),
    .A2(_0209_),
    .A3(_0208_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2441_ (.A1(_0210_),
    .A2(_0211_),
    .A3(_0212_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2442_ (.A1(_0157_),
    .A2(_0213_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2443_ (.A1(_0513_),
    .A2(_0213_),
    .B(_0214_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2444_ (.A1(_0203_),
    .A2(_0216_),
    .B(_0160_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2445_ (.I(_1292_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2446_ (.I(_1301_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2447_ (.I(_1225_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2448_ (.A1(_0220_),
    .A2(_1228_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2449_ (.A1(_0219_),
    .A2(_0221_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2450_ (.A1(_0173_),
    .A2(_0222_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2451_ (.A1(_1252_),
    .A2(_0036_),
    .B(_1244_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2452_ (.A1(_1232_),
    .A2(_0224_),
    .B(_0079_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2453_ (.A1(_0056_),
    .A2(_1186_),
    .B1(_1234_),
    .B2(_1204_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2454_ (.I(_1271_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2455_ (.A1(_0225_),
    .A2(_0131_),
    .B1(_0227_),
    .B2(_0228_),
    .C(_0094_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2456_ (.A1(_0223_),
    .A2(_0229_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2457_ (.I(_1307_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2458_ (.I(_0231_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2459_ (.A1(_0232_),
    .A2(_0176_),
    .B(_0163_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2460_ (.A1(_0230_),
    .A2(_0233_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2461_ (.A1(_0218_),
    .A2(_0234_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2462_ (.A1(_0179_),
    .A2(_0190_),
    .B(_0516_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2463_ (.A1(_0205_),
    .A2(_1159_),
    .B(_0117_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2464_ (.A1(_0151_),
    .A2(_0238_),
    .B(_1200_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2465_ (.A1(_1186_),
    .A2(_1277_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2466_ (.A1(_1344_),
    .A2(_0154_),
    .A3(_0240_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2467_ (.A1(_0041_),
    .A2(_0151_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2468_ (.A1(_0239_),
    .A2(_0241_),
    .A3(_0242_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2469_ (.A1(_0236_),
    .A2(_0243_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _2470_ (.A1(_0217_),
    .A2(_0235_),
    .A3(_0244_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2471_ (.A1(_0193_),
    .A2(_0196_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2472_ (.A1(_0197_),
    .A2(_0199_),
    .B(_0246_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2473_ (.A1(_0202_),
    .A2(_0245_),
    .A3(_0247_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2474_ (.I(_0249_),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2475_ (.I(_0181_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2476_ (.A1(_1338_),
    .A2(_0089_),
    .B(_0220_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2477_ (.I(_1342_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2478_ (.A1(_0079_),
    .A2(_0090_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2479_ (.I(_0089_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2480_ (.A1(_0254_),
    .A2(_0252_),
    .A3(_0253_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2481_ (.A1(_0252_),
    .A2(_0040_),
    .A3(_0253_),
    .B(_0255_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2482_ (.A1(_0251_),
    .A2(_0091_),
    .B(_0256_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2483_ (.A1(_0204_),
    .A2(_0115_),
    .B1(_1283_),
    .B2(_1284_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2484_ (.A1(_0220_),
    .A2(_0150_),
    .A3(_0052_),
    .B(_0109_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2485_ (.A1(_0250_),
    .A2(_0257_),
    .B1(_0259_),
    .B2(_0260_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2486_ (.A1(_0087_),
    .A2(_0213_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2487_ (.A1(_0157_),
    .A2(_0262_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2488_ (.A1(_0261_),
    .A2(_0263_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2489_ (.A1(_0102_),
    .A2(_0264_),
    .B(_0160_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2490_ (.I(_0182_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2491_ (.I(_0228_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2492_ (.I(_0207_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2493_ (.A1(_0268_),
    .A2(_0254_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2494_ (.A1(_0266_),
    .A2(_0267_),
    .A3(_0270_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2495_ (.I(_1197_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2496_ (.I(_0272_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2497_ (.A1(_0252_),
    .A2(_0258_),
    .A3(_0271_),
    .B1(_0253_),
    .B2(_0273_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2498_ (.A1(_0252_),
    .A2(_0258_),
    .A3(_0273_),
    .A4(_0253_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2499_ (.A1(_0250_),
    .A2(_0275_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2500_ (.A1(_0219_),
    .A2(_0109_),
    .B1(_0274_),
    .B2(_0276_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2501_ (.A1(_0167_),
    .A2(_0175_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2502_ (.A1(_0122_),
    .A2(_0108_),
    .A3(_0278_),
    .A4(_0230_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2503_ (.A1(_0231_),
    .A2(_0279_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2504_ (.I(_1307_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2505_ (.A1(_0122_),
    .A2(_0108_),
    .A3(_0278_),
    .A4(_0230_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2506_ (.A1(_0282_),
    .A2(_0277_),
    .A3(_0283_),
    .B(_0218_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2507_ (.A1(_0277_),
    .A2(_0281_),
    .B(_0284_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2508_ (.A1(_1182_),
    .A2(_0188_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2509_ (.I0(_0187_),
    .I1(_0286_),
    .S(_0094_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2510_ (.A1(_0137_),
    .A2(_0138_),
    .A3(_0287_),
    .A4(_0243_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2511_ (.A1(_0515_),
    .A2(_0288_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2512_ (.I(_0181_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2513_ (.I(_1182_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2514_ (.A1(_0164_),
    .A2(_0082_),
    .B(_0292_),
    .C(_0168_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2515_ (.A1(_0228_),
    .A2(_1203_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2516_ (.A1(_0131_),
    .A2(_0206_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2517_ (.I(_0295_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2518_ (.A1(_0290_),
    .A2(_0293_),
    .A3(_0294_),
    .B1(_0173_),
    .B2(_0296_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2519_ (.I0(_0289_),
    .I1(\p_shaping_I.p_shaping_I.bit_in ),
    .S(_0297_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2520_ (.A1(_0265_),
    .A2(_0285_),
    .A3(_0298_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2521_ (.A1(_0235_),
    .A2(_0244_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2522_ (.A1(_0235_),
    .A2(_0244_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2523_ (.A1(_0217_),
    .A2(_0300_),
    .B(_0301_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2524_ (.A1(_0299_),
    .A2(_0302_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2525_ (.A1(_0202_),
    .A2(_0245_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _2526_ (.A1(_0193_),
    .A2(_0196_),
    .B1(_0197_),
    .B2(_0199_),
    .C1(_0202_),
    .C2(_0245_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2527_ (.A1(_0304_),
    .A2(_0305_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2528_ (.A1(_0303_),
    .A2(_0306_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2529_ (.I(_0307_),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2530_ (.A1(_0285_),
    .A2(_0298_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2531_ (.A1(_0285_),
    .A2(_0298_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2532_ (.A1(_0265_),
    .A2(_0308_),
    .A3(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2533_ (.A1(_0075_),
    .A2(_0030_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2534_ (.A1(_1331_),
    .A2(_0312_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2535_ (.I(_0263_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2536_ (.A1(_0115_),
    .A2(_0165_),
    .B1(_0185_),
    .B2(_0111_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2537_ (.I(_0268_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2538_ (.A1(_0316_),
    .A2(_1266_),
    .A3(_0184_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2539_ (.A1(_0254_),
    .A2(_1159_),
    .B(_0268_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2540_ (.A1(_0057_),
    .A2(_0318_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2541_ (.A1(_0154_),
    .A2(_0317_),
    .A3(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2542_ (.I(_0267_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2543_ (.A1(_0182_),
    .A2(_0251_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2544_ (.A1(_0321_),
    .A2(_0323_),
    .B(_0269_),
    .C(_0250_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2545_ (.A1(_1332_),
    .A2(_0315_),
    .B(_0320_),
    .C(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2546_ (.A1(_0512_),
    .A2(_0325_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2547_ (.A1(_0314_),
    .A2(_0325_),
    .B(_0326_),
    .C(_0203_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2548_ (.A1(_1212_),
    .A2(_0313_),
    .A3(_0327_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2549_ (.A1(_0082_),
    .A2(_0165_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2550_ (.A1(_0329_),
    .A2(_0294_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2551_ (.A1(_0207_),
    .A2(_0272_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2552_ (.A1(_0267_),
    .A2(_0184_),
    .A3(_0050_),
    .A4(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2553_ (.A1(_0330_),
    .A2(_0332_),
    .B(_0250_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2554_ (.A1(_0232_),
    .A2(_0279_),
    .B(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2555_ (.I(_0334_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2556_ (.A1(_0282_),
    .A2(_0283_),
    .A3(_0336_),
    .B(_1292_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2557_ (.A1(_0335_),
    .A2(_0337_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2558_ (.A1(_0220_),
    .A2(_1290_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2559_ (.A1(_0182_),
    .A2(_0205_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2560_ (.A1(_0207_),
    .A2(_0340_),
    .B(_0024_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2561_ (.A1(_0339_),
    .A2(_1228_),
    .B(_0341_),
    .C(_0181_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2562_ (.A1(_0161_),
    .A2(_1270_),
    .B(_0342_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2563_ (.A1(_0289_),
    .A2(_0343_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2564_ (.A1(_0338_),
    .A2(_0345_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2565_ (.A1(_0328_),
    .A2(_0346_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2566_ (.A1(_0308_),
    .A2(_0310_),
    .B(_0347_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2567_ (.A1(_0308_),
    .A2(_0310_),
    .A3(_0347_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2568_ (.A1(_0348_),
    .A2(_0349_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2569_ (.I(_0299_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2570_ (.A1(_0351_),
    .A2(_0302_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2571_ (.A1(_0304_),
    .A2(_0303_),
    .A3(_0305_),
    .B(_0352_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2572_ (.A1(_0350_),
    .A2(_0353_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2573_ (.I(_0354_),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2574_ (.A1(_0021_),
    .A2(_0103_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2575_ (.A1(_1200_),
    .A2(_0319_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2576_ (.A1(_0316_),
    .A2(_0115_),
    .B1(_1245_),
    .B2(_0165_),
    .C(_0292_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2577_ (.A1(_0081_),
    .A2(_0318_),
    .B(_0358_),
    .C(_0290_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2578_ (.A1(_0154_),
    .A2(_1164_),
    .A3(_1343_),
    .B1(_0357_),
    .B2(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2579_ (.A1(_0513_),
    .A2(_0360_),
    .B(_1331_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2580_ (.A1(_0314_),
    .A2(_0360_),
    .B(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2581_ (.A1(_0356_),
    .A2(_0362_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2582_ (.A1(_0205_),
    .A2(_1177_),
    .B(_0268_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2583_ (.A1(_0266_),
    .A2(_0251_),
    .B1(_0364_),
    .B2(_0147_),
    .C(_0267_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2584_ (.A1(_0288_),
    .A2(_0366_),
    .B(_0183_),
    .C(_0515_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2585_ (.A1(_0183_),
    .A2(_0515_),
    .B(_0367_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2586_ (.A1(_0228_),
    .A2(_0146_),
    .A3(_0209_),
    .A4(_0331_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2587_ (.A1(_0146_),
    .A2(_0224_),
    .A3(_0091_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2588_ (.A1(_0242_),
    .A2(_0369_),
    .A3(_0370_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2589_ (.A1(_0282_),
    .A2(_0149_),
    .B(_0281_),
    .C(_0371_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2590_ (.A1(_1307_),
    .A2(_0371_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2591_ (.A1(_0218_),
    .A2(_0372_),
    .A3(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2592_ (.A1(_0368_),
    .A2(_0374_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2593_ (.A1(_0363_),
    .A2(_0375_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2594_ (.I(_0377_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2595_ (.A1(_0328_),
    .A2(_0346_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2596_ (.A1(_0335_),
    .A2(_0337_),
    .A3(_0345_),
    .B(_0379_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2597_ (.A1(_0378_),
    .A2(_0380_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2598_ (.I(_0349_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2599_ (.A1(_0352_),
    .A2(_0348_),
    .B(_0382_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2600_ (.A1(_0304_),
    .A2(_0303_),
    .A3(_0305_),
    .A4(_0350_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2601_ (.A1(_0383_),
    .A2(_0384_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2602_ (.A1(_0381_),
    .A2(_0385_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2603_ (.I(_0386_),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2604_ (.A1(_0368_),
    .A2(_0374_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2605_ (.A1(_0363_),
    .A2(_0375_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2606_ (.I(_0290_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2607_ (.I(_0316_),
    .Z(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2608_ (.A1(_0391_),
    .A2(_0340_),
    .B(_0224_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2609_ (.A1(_0321_),
    .A2(_0209_),
    .B1(_0091_),
    .B2(_0392_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2610_ (.I(_0290_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2611_ (.A1(_0394_),
    .A2(_0366_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2612_ (.A1(_0390_),
    .A2(_0393_),
    .B(_0395_),
    .C(_0314_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2613_ (.A1(_0390_),
    .A2(_0393_),
    .B(_0395_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2614_ (.A1(_0087_),
    .A2(_0398_),
    .B(_0203_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2615_ (.A1(_0396_),
    .A2(_0399_),
    .B(_0356_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2616_ (.A1(_0219_),
    .A2(_0272_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2617_ (.A1(_0292_),
    .A2(_0331_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2618_ (.A1(_0294_),
    .A2(_0401_),
    .B(_0402_),
    .C(_0394_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2619_ (.A1(_0232_),
    .A2(_0279_),
    .B(_0403_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2620_ (.A1(_0232_),
    .A2(_0403_),
    .B(_0404_),
    .C(_0062_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2621_ (.A1(_0146_),
    .A2(_1203_),
    .A3(_0219_),
    .B(_0172_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2622_ (.A1(_0289_),
    .A2(_0406_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2623_ (.A1(_0516_),
    .A2(_0406_),
    .B(_0407_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2624_ (.A1(_0400_),
    .A2(_0405_),
    .A3(_0409_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2625_ (.A1(_0388_),
    .A2(_0389_),
    .B(_0410_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2626_ (.A1(_0388_),
    .A2(_0389_),
    .A3(_0410_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2627_ (.A1(_0411_),
    .A2(_0412_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2628_ (.A1(_0378_),
    .A2(_0380_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2629_ (.A1(_0383_),
    .A2(_0384_),
    .B(_0381_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2630_ (.A1(_0414_),
    .A2(_0415_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2631_ (.A1(_0413_),
    .A2(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2632_ (.I(_0417_),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2633_ (.A1(_0316_),
    .A2(_0321_),
    .A3(_0272_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2634_ (.A1(_0394_),
    .A2(_0402_),
    .A3(_0419_),
    .B(_0281_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2635_ (.A1(_0394_),
    .A2(_0282_),
    .A3(_0402_),
    .A4(_0419_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2636_ (.A1(_0062_),
    .A2(_0421_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2637_ (.A1(_0172_),
    .A2(_0289_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2638_ (.A1(_0172_),
    .A2(_0516_),
    .B(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2639_ (.A1(_0420_),
    .A2(_0422_),
    .A3(_0424_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2640_ (.I(_0425_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2641_ (.A1(_0420_),
    .A2(_0422_),
    .B(_0424_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2642_ (.A1(_0426_),
    .A2(_0427_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2643_ (.A1(_1331_),
    .A2(_0263_),
    .B(_0313_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2644_ (.A1(_0391_),
    .A2(_1228_),
    .B(_0294_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2645_ (.A1(_0041_),
    .A2(_0222_),
    .B1(_0431_),
    .B2(_0390_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2646_ (.A1(_0430_),
    .A2(_0432_),
    .Z(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2647_ (.A1(_1212_),
    .A2(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2648_ (.A1(_0428_),
    .A2(_0434_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2649_ (.A1(_0405_),
    .A2(_0409_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2650_ (.A1(_0405_),
    .A2(_0409_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2651_ (.A1(_0400_),
    .A2(_0436_),
    .B(_0437_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2652_ (.A1(_0435_),
    .A2(_0438_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2653_ (.A1(_0378_),
    .A2(_0380_),
    .B(_0411_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2654_ (.A1(_0415_),
    .A2(_0441_),
    .B(_0412_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2655_ (.A1(_0439_),
    .A2(_0442_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2656_ (.I(_0443_),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2657_ (.A1(_0426_),
    .A2(_0427_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2658_ (.A1(_0444_),
    .A2(_0434_),
    .B(_0426_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2659_ (.A1(_1332_),
    .A2(_0221_),
    .B(_1256_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2660_ (.A1(_0314_),
    .A2(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2661_ (.A1(_0513_),
    .A2(_0446_),
    .B(_0447_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2662_ (.A1(_0203_),
    .A2(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2663_ (.A1(_0356_),
    .A2(_0449_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2664_ (.A1(_0428_),
    .A2(_0451_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2665_ (.A1(_0435_),
    .A2(_0438_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2666_ (.A1(_0415_),
    .A2(_0441_),
    .B(_0439_),
    .C(_0412_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2667_ (.A1(_0453_),
    .A2(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2668_ (.A1(_0445_),
    .A2(_0452_),
    .A3(_0455_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2669_ (.I(_0456_),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2670_ (.A1(_0445_),
    .A2(_0452_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2671_ (.A1(_0453_),
    .A2(_0454_),
    .A3(_0457_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2672_ (.A1(_1212_),
    .A2(_0430_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2673_ (.A1(_0427_),
    .A2(_0451_),
    .B(_0425_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2674_ (.A1(_0445_),
    .A2(_0452_),
    .B1(_0459_),
    .B2(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2675_ (.A1(_0459_),
    .A2(_0461_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2676_ (.A1(_0458_),
    .A2(_0462_),
    .B(_0463_),
    .ZN(net9));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2677_ (.A1(_1263_),
    .A2(_1264_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2678_ (.A1(_1322_),
    .A2(_0464_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2679_ (.I(_0465_),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2680_ (.A1(\p_shaping_Q.p_shaping_I.counter[0] ),
    .A2(_1098_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2681_ (.A1(_0007_),
    .A2(_0466_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2682_ (.A1(net67),
    .A2(net3),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2683_ (.I(_0467_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2684_ (.I(_0469_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2685_ (.A1(_1338_),
    .A2(_0470_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2686_ (.I(_0471_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2687_ (.I(_0469_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2688_ (.A1(_0266_),
    .A2(_0472_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2689_ (.A1(net47),
    .A2(_0056_),
    .A3(_0472_),
    .B(_0473_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2690_ (.A1(_0266_),
    .A2(_0204_),
    .A3(net65),
    .A4(net3),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2691_ (.A1(_0254_),
    .A2(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2692_ (.A1(_0050_),
    .A2(_0472_),
    .B(_0475_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2693_ (.A1(_1290_),
    .A2(_0467_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2694_ (.A1(_0391_),
    .A2(_0477_),
    .Z(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2695_ (.I(_0478_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2696_ (.A1(_0183_),
    .A2(_0269_),
    .A3(_0469_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2697_ (.A1(_0391_),
    .A2(_0321_),
    .A3(_0477_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2698_ (.A1(_0270_),
    .A2(_0474_),
    .B(_0292_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2699_ (.A1(_0480_),
    .A2(_0481_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2700_ (.A1(_0479_),
    .A2(_0482_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2701_ (.A1(_0390_),
    .A2(_0480_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2702_ (.A1(_0479_),
    .A2(_0483_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2703_ (.A1(_0863_),
    .A2(_0469_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2704_ (.I(_0485_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2705_ (.A1(_0883_),
    .A2(_0470_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2706_ (.A1(net48),
    .A2(_0784_),
    .A3(_0472_),
    .B(_0486_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2707_ (.A1(_0783_),
    .A2(net63),
    .A3(net3),
    .A4(_0864_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2708_ (.A1(_0619_),
    .A2(_0470_),
    .B(_0887_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2709_ (.A1(_0487_),
    .A2(_0488_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2710_ (.I(_0489_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2711_ (.A1(_0885_),
    .A2(_0487_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2712_ (.I(_0490_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2713_ (.A1(_0505_),
    .A2(_0470_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2714_ (.A1(_0679_),
    .A2(_0467_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2715_ (.A1(_0701_),
    .A2(_0493_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2716_ (.A1(_0492_),
    .A2(_0494_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2717_ (.A1(_1099_),
    .A2(_0493_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2718_ (.A1(_1084_),
    .A2(_0495_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2719_ (.A1(_0492_),
    .A2(_0496_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2720_ (.A1(_0218_),
    .A2(\p_shaping_I.p_shaping_I.counter[0] ),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2721_ (.A1(_0021_),
    .A2(_0497_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2722_ (.D(_0006_),
    .RN(net56),
    .CLK(net49),
    .Q(\p_shaping_Q.p_shaping_I.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2723_ (.D(_0007_),
    .RN(net56),
    .CLK(net49),
    .Q(\p_shaping_Q.p_shaping_I.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2724_ (.D(\gen_sym.Reg_2M.data_in ),
    .RN(net52),
    .CLK(net45),
    .Q(\gen_sym.Reg_Sym.data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2725_ (.D(\gen_sym.Reg_2M.data_out ),
    .RN(net53),
    .CLK(net45),
    .Q(\gen_sym.Reg_Sym.data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2726_ (.D(\gen_sym.Reg_2M.data_in ),
    .RN(net52),
    .CLK(\gen_sym.Reg_2M.enable ),
    .Q(\gen_sym.Reg_2M.data_out ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2727_ (.D(\mapper.bit_Q[1] ),
    .RN(net53),
    .CLK(net48),
    .Q(\p_shaping_Q.p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2728_ (.D(\p_shaping_I.p_shaping_I.bit_in_1 ),
    .RN(net60),
    .CLK(net46),
    .Q(\p_shaping_I.p_shaping_I.bit_in_2 ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _2729_ (.D(_0000_),
    .Q(\p_shaping_I.p_shaping_I.ctl_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2730_ (.D(_0008_),
    .RN(net54),
    .CLK(net64),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2731_ (.D(_0009_),
    .RN(net56),
    .CLK(net65),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2732_ (.D(_0010_),
    .RN(net56),
    .CLK(net65),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2733_ (.D(_0011_),
    .RN(net59),
    .CLK(net67),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2734_ (.D(_0012_),
    .RN(net57),
    .CLK(net65),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2735_ (.D(_0013_),
    .RN(net57),
    .CLK(net66),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2736_ (.D(\p_shaping_I.p_shaping_I.bit_in ),
    .RN(net60),
    .CLK(net46),
    .Q(\p_shaping_I.p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2737_ (.D(\p_shaping_Q.p_shaping_I.bit_in_1 ),
    .RN(net59),
    .CLK(net48),
    .Q(\p_shaping_Q.p_shaping_I.bit_in_2 ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _2738_ (.D(_0002_),
    .Q(\p_shaping_Q.p_shaping_I.ctl_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _2739_ (.D(_0014_),
    .SETN(net55),
    .CLK(net63),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2740_ (.D(_0015_),
    .RN(net52),
    .CLK(net64),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2741_ (.D(_0016_),
    .RN(net55),
    .CLK(net63),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _2742_ (.D(_0017_),
    .SETN(net55),
    .CLK(net63),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _2743_ (.D(_0018_),
    .SETN(net52),
    .CLK(net64),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2744_ (.D(_0019_),
    .RN(net53),
    .CLK(net64),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2745_ (.D(net44),
    .RN(net59),
    .CLK(net49),
    .Q(\p_shaping_Q.p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2746_ (.D(_0020_),
    .RN(net60),
    .CLK(net46),
    .Q(\p_shaping_I.p_shaping_I.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2747_ (.D(_0021_),
    .RN(net60),
    .CLK(net46),
    .Q(\p_shaping_I.p_shaping_I.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(ACK),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input2 (.I(Bit_In),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input3 (.I(EN),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(REQ_SAMPLE),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(RST),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output6 (.I(net6),
    .Z(I[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output7 (.I(net7),
    .Z(I[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output8 (.I(net8),
    .Z(I[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output9 (.I(net9),
    .Z(I[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output10 (.I(net10),
    .Z(I[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output11 (.I(net11),
    .Z(I[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output12 (.I(net12),
    .Z(I[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output13 (.I(net13),
    .Z(I[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net14),
    .Z(I[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output15 (.I(net15),
    .Z(I[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(I[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(I[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(I[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(Q[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(Q[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(Q[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(Q[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(Q[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(Q[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(Q[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(Q[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(Q[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(Q[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(Q[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(Q[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(Q[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(addI[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(addI[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(addI[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(addI[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(addI[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(addI[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(addQ[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(addQ[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(addQ[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(addQ[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(addQ[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(addQ[5]));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout44 (.I(\p_shaping_Q.p_shaping_I.bit_in ),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout45 (.I(net47),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout46 (.I(_0004_),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout47 (.I(_0004_),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout48 (.I(_0005_),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout49 (.I(_0005_),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout50 (.I(net42),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout51 (.I(net40),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout52 (.I(net54),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout53 (.I(net54),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout54 (.I(net55),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout55 (.I(net62),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout56 (.I(net58),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout57 (.I(net58),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout58 (.I(net61),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout59 (.I(net61),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout60 (.I(net62),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout61 (.I(net62),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout62 (.I(net5),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout63 (.I(net68),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout64 (.I(net68),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout65 (.I(net66),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout66 (.I(net67),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout67 (.I(net68),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout68 (.I(net4),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(ACK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(Bit_In));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(EN));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(REQ_SAMPLE));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(RST));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__D (.I(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__D (.I(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__A1 (.I(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__A1 (.I(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__A1 (.I(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__A2 (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__A1 (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__B (.I(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__A2 (.I(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__B (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__I (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__C (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__B (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2313__I (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__A2 (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__A2 (.I(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A2 (.I(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__I (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__B (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A1 (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__A1 (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A2 (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__A1 (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A2 (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__A1 (.I(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__A1 (.I(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2440__A1 (.I(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__C (.I(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__I (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__B (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A1 (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1368__A1 (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A3 (.I(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2285__A1 (.I(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A2 (.I(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A2 (.I(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A2 (.I(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A1 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A1 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A1 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__A1 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2329__A1 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A1 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A1 (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A3 (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__C (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A2 (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A3 (.I(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A2 (.I(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__B1 (.I(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__A3 (.I(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2297__A1 (.I(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A2 (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A1 (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__A2 (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2295__A2 (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__A1 (.I(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A2 (.I(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__A2 (.I(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A2 (.I(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A3 (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__B (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A3 (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__A1 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__I (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__B (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1367__B (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A1 (.I(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__I (.I(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1368__A2 (.I(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__A2 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__A1 (.I(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__A1 (.I(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A2 (.I(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__A1 (.I(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A2 (.I(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__B1 (.I(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A3 (.I(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__I (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1376__A1 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A1 (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A1 (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A1 (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2325__C (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__I (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A2 (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A1 (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__A1 (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__B1 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A3 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__A2 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2329__B (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__A2 (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__S (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__C (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__I (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2332__A1 (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2164__A1 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__A1 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__I (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1375__A1 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__A2 (.I(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__A1 (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__I (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A2 (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__B (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__A1 (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A1 (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__B2 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__B (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__A1 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__A1 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A2 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A1 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A2 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__B2 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__B (.I(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__A2 (.I(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__A2 (.I(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__A2 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__I (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A1 (.I(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A1 (.I(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A2 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__I (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2108__A1 (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1380__I (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1374__A1 (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A1 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A2 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__A1 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A2 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__A2 (.I(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A1 (.I(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__A1 (.I(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__A1 (.I(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A2 (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__A2 (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__A2 (.I(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__A2 (.I(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2374__A2 (.I(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__B2 (.I(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A3 (.I(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__A2 (.I(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A2 (.I(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__A2 (.I(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A2 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A2 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__A1 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1375__A4 (.I(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2467__A2 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__A1 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A2 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A2 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__C (.I(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A1 (.I(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__B (.I(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1376__A2 (.I(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A2 (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A1 (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A1 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A1 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__B (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1377__A2 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__B1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__C (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__I (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A1 (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__I0 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__A2 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A2 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2418__A2 (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A2 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A2 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__A2 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A2 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__A2 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2471__A2 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A2 (.I(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__B2 (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__A2 (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__A2 (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__A2 (.I(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A1 (.I(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A2 (.I(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1385__A1 (.I(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__A1 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__A2 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__A1 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__A1 (.I(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__I (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A2 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__A2 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A2 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__B (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2122__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2098__I (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1384__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A3 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__B (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A2 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A2 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__A1 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2491__I (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__B2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2505__A4 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__A4 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A1 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A1 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A1 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__A2 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A4 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2469__A2 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A2 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A2 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__A3 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__B (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__A2 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A2 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1384__A3 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__I (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__B (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__C (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A1 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A1 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A2 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__A2 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A2 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1385__A2 (.I(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__B1 (.I(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A1 (.I(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__C (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__I (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A2 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__A2 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__B (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__I (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1386__A2 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2507__A1 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__A2 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A2 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__I (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2606__I (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__C (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2337__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1444__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1432__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1388__I (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__B (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__C (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__B (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__S (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A3 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__I (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__I (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A1 (.I(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1415__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__I (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__B (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2557__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__I (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2605__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A1 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2604__A2 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A2 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1409__A2 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1397__I (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2645__B2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__C (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1563__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1552__A3 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1415__A2 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A1 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1575__B (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__I (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1469__I (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1401__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A3 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__I (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1504__I (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1486__I (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__I (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1400__A3 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__A4 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__A3 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__A1 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__B (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__A3 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A2 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__I (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1407__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__I (.I(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__I (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1485__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1473__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1412__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1405__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__I (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__I (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1533__I (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1475__A2 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1460__I (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1405__A2 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2703__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__A3 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__I (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__I (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A2 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__A3 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2692__A2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A3 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A2 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__A3 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1406__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1407__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1544__A1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1501__A1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1481__I (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1411__A1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1413__A2 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1414__B (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__A1 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1415__A3 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2713__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1440__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1416__I (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1422__A1 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1419__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__A1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1428__I (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1420__I (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__B (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1425__I (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__A1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1433__A1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1446__I (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1439__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1431__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1430__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A1 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__B (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1431__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__A1 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A1 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__I0 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1441__A1 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__B (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__B (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__A1 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1437__I (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1990__A1 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1906__I1 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A1 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1439__A2 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__B (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1881__A1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__B (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1450__I (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1920__A1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__B (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__A1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1451__I (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2026__I (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__C (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__B2 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1497__A1 (.I(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1595__B (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__A1 (.I(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1612__I (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1494__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1463__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__B (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1523__B (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1459__A1 (.I(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__I (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__B (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1503__B (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__I (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__B (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1463__B (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1786__I (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1535__A1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1472__A1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1676__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1472__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1712__A1 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__A1 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1547__A1 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1472__C (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__A3 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1567__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1535__B (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__A2 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1648__A2 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__A2 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1476__I (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__B (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1552__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1488__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1584__I (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1570__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1515__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1482__I (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__I (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1647__I (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1487__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__A1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__I (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__I (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1487__B (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1850__B (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1488__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2016__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__B2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__B2 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__S (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1494__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__B (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__B (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1594__A1 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1493__A1 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__I (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A1 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1563__A1 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1493__A2 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__A1 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1494__B (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__A2 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1600__A2 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1578__I (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1499__I (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__I (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A3 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1626__I (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__A2 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1532__I (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__B1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__A2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1538__I (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1507__A2 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__B2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1570__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1536__I0 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1511__A1 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1514__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1904__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1513__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__B1 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1514__B (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1608__I (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1516__A2 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__B1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__B1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__B1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__I (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1524__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1591__I (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1545__A1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1536__I1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1522__A1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__A1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1546__A1 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1522__A3 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1579__B2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1524__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__A2 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__B2 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1524__A3 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__B2 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A1 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A1 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__A2 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1529__A1 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1830__I (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1730__I (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1527__I (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1934__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1529__A2 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__I0 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1733__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1585__A2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1547__A3 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1535__A2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A2 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1537__A2 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__A1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__B1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__A1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__A2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__A1 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1542__B2 (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1567__C (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1541__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__I (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1541__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1553__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1564__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1546__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__C (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1599__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1546__B (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1993__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__A3 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A1 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__B (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__B (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1641__I (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__B (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1550__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__B (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__C (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1553__B (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__B (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__A2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1553__C (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1557__I (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1633__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__C (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1634__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1582__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__B (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__B (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1567__B1 (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__A2 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A2 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__I1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1566__A2 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__A1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1596__I (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1592__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1579__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__A3 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A3 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__A2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__I (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__A1 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__A1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__A1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1585__A1 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__A3 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__A2 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__A2 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1592__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__I (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1659__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1594__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__B (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1850__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1613__A2 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__A2 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1678__B (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1662__A3 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1599__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__A1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__B (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__I (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__I (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__A4 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1685__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__C (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__A2 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__A2 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__A3 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1635__B (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A2 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__A2 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__I0 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1609__A2 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__A3 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1911__A3 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__B1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__A1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__B2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__A1 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__A2 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1685__A1 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__B1 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1615__I (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__B2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1979__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1768__B (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__C (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__B (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__I (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__C (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__S (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1621__I (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__B (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1904__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__B (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__B (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__I (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1916__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__I (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__C (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__B2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1768__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1738__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__A3 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__A3 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1981__B2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1957__I (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__I (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__I (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__B2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__B (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__A2 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__A2 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1659__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__C (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__B (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A3 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__B (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__A3 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__A2 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A3 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1657__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1859__I (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__B2 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A2 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__A1 (.I(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__B1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__A2 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__A2 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1742__A3 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__A2 (.I(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1822__A2 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__B (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1667__C (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__A3 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__A2 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__B1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__C (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__I (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__B2 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1720__B (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1681__C (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1942__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1804__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1683__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A3 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1726__A3 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__A2 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__A2 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1696__I (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A3 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1691__I (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1703__B2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__A1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__B1 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1703__B1 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__A4 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A2 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__A2 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__B2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1710__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1714__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__A3 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__B2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__A2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__A2 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__B (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__A3 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__A3 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1729__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__B2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1836__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A2 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__B2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A1 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__I (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__A1 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__A1 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__A1 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1768__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__B1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__C (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1943__A2 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__C (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__A2 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__A2 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__B1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1938__A1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__A2 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A2 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__A3 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A3 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1747__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1857__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__B (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__C (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1984__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1760__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__B (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__B (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__A2 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1769__A1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__A4 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A4 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__B (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1772__A4 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__I (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__I (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1962__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1880__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__B (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__A1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__B2 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1799__I (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A1 (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2703__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__A2 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__A4 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A2 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1823__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__B1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__A2 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__A3 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1878__A3 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1795__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1846__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__B (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__I (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A2 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1953__A2 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__B (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__B1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1996__A2 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__A2 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1911__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__A1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1820__B (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__B (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__A1 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__B2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1939__A1 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__B1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1812__B1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__B (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2030__A1 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1977__A2 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A2 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A3 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__B (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A2 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1894__B (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__B (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1827__A1 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1865__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1828__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1831__B (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1829__A4 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__B2 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1831__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__I (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__B1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__A3 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__B (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1850__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1890__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__A2 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2068__A1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__A3 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1854__A1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1942__A2 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__C (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__A1 (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2031__B (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__C (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__A2 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1864__B2 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__A3 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1925__A3 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__B (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__A2 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__B1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1916__A3 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__A3 (.I(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1878__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A2 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__A3 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__B (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__A3 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__B (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__A3 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1936__A3 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1908__B (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__A4 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__B1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1920__A4 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1933__I (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1994__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__B2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1941__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1945__S (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__A1 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__B (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__A3 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__I (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__A2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1991__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__I (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__B2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A2 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__B (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__A2 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2055__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2052__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2032__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2028__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__A2 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__A2 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__A2 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__B (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__A1 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2066__A2 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__A2 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__A2 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__A2 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__I (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__A3 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2092__I (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A2 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__B (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A1 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2177__I (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2102__I (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2096__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__B2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__I (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2097__A2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__B2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__C (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__A1 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2256__I (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__A2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2101__I (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__I (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2103__B (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__B (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__I (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2106__I (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2289__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__A3 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__B (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__B (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__A1 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2111__B (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__C (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__I (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__B (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__I (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__I (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2293__B (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__C (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__A1 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__A1 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A1 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__A2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2205__A1 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__A1 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A1 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__B (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__A2 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__A1 (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__I (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A2 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__A1 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__A2 (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2154__B (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__I (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1349__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__C (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2251__I (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A1 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__B (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__A2 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__I (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2414__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__B (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A2 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__B (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__B2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2130__I (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__B (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__B1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__B (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__A1 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__A1 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2132__I (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A2 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__A2 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1363__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__B2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__B1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A2 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2276__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__I (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__I (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__A1 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__I (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2213__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__I (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__A2 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2189__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2186__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A2 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__A2 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A3 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2145__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__B (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__B (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2176__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__B (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2349__A2 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A3 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__A2 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2287__I (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2150__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2321__A1 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__C (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2151__C (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__I (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A1 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A1 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1358__A1 (.I(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2275__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2231__A2 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__A2 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2155__I (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__A1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__B (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__C (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__B (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2275__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__A2 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__A1 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__B1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A2 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__B1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A2 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__B2 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__B1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__B2 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__A2 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2197__I (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__B (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__C (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__B (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2300__I (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__B (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__I (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__B1 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A1 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__A2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__A2 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__B (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__B (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2175__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2399__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__B2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2366__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2275__C (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2179__C (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__A1 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__A1 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2218__A1 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__A1 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__B (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2182__C (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2183__I (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2194__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__B (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__I (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__A1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__B (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__B (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2370__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2209__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__B (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2205__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__A1 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__B2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__A1 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A1 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2174__I (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2133__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1367__A3 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1357__A3 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2368__C (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__B (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__I (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2205__C (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__B1 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__B2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__B (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__B (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1358__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2556__B (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__I (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2359__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2230__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__C (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2279__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2217__I (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2386__I (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__B (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2292__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2222__A3 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A2 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2221__A2 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2226__B1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A1 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2342__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2284__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__B (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2227__A3 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A1 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__I (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__I (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2229__A1 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__I (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2232__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2438__C (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2398__A1 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__A2 (.I(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2345__A2 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__A3 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2434__B (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__A2 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__A3 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2304__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2309__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2643__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__B (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2272__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__B2 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__I (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__A3 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A2 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__I (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__B1 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2578__A3 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2361__I (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__I (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1363__B (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__D (.I(\p_shaping_I.p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__I1 (.I(\p_shaping_I.p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2286__B (.I(\p_shaping_I.p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2240__A1 (.I(\p_shaping_I.p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(\p_shaping_Q.p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__I (.I(\p_shaping_Q.p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__D (.I(\p_shaping_Q.p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A1 (.I(\p_shaping_Q.p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1945__I0 (.I(\p_shaping_Q.p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1434__I (.I(\p_shaping_Q.p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__I (.I(\p_shaping_Q.p_shaping_I.bit_in_2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__I (.I(\p_shaping_Q.p_shaping_I.bit_in_2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__B (.I(\p_shaping_Q.p_shaping_I.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1526__A2 (.I(\p_shaping_Q.p_shaping_I.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1449__I (.I(\p_shaping_Q.p_shaping_I.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1442__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__A3 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__A4 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1442__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout68_I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout62_I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output7_I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output9_I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output13_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2107__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1354__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__A1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1372__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1352__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1373__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1347__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1381__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1350__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1346__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1370__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1366__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1359__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1371__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1364__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1360__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1501__A2 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1389__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1454__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1410__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1392__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1403__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1393__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output43_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1458__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1408__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1604__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1436__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__D (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout45_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1444__A2 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__CLK (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1448__A2 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2723__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__CLK (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1412__A2 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1402__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__SETN (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__RN (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__RN (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__RN (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__RN (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__RN (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2725__RN (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1427__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2742__SETN (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__RN (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__SETN (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__RN (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__RN (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__RN (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1438__A1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout59_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout60_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout61_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__CLK (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__CLK (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__A3 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout66_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__CLK (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout67_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout63_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout64_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_508 ();
endmodule

