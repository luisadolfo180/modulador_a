magic
tech gf180mcuC
magscale 1 10
timestamp 1670198983
<< metal1 >>
rect 6738 56590 6750 56642
rect 6802 56639 6814 56642
rect 7634 56639 7646 56642
rect 6802 56593 7646 56639
rect 6802 56590 6814 56593
rect 7634 56590 7646 56593
rect 7698 56590 7710 56642
rect 40338 56590 40350 56642
rect 40402 56639 40414 56642
rect 41122 56639 41134 56642
rect 40402 56593 41134 56639
rect 40402 56590 40414 56593
rect 41122 56590 41134 56593
rect 41186 56590 41198 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 4622 56306 4674 56318
rect 4622 56242 4674 56254
rect 16382 56306 16434 56318
rect 16382 56242 16434 56254
rect 27470 56306 27522 56318
rect 27470 56242 27522 56254
rect 31278 56306 31330 56318
rect 31278 56242 31330 56254
rect 33630 56306 33682 56318
rect 33630 56242 33682 56254
rect 38334 56306 38386 56318
rect 38334 56242 38386 56254
rect 38782 56306 38834 56318
rect 38782 56242 38834 56254
rect 39454 56306 39506 56318
rect 39454 56242 39506 56254
rect 42814 56306 42866 56318
rect 42814 56242 42866 56254
rect 14142 56194 14194 56206
rect 2258 56142 2270 56194
rect 2322 56142 2334 56194
rect 14142 56130 14194 56142
rect 22654 56194 22706 56206
rect 22654 56130 22706 56142
rect 26126 56194 26178 56206
rect 26126 56130 26178 56142
rect 26574 56194 26626 56206
rect 43598 56194 43650 56206
rect 30258 56142 30270 56194
rect 30322 56142 30334 56194
rect 35186 56142 35198 56194
rect 35250 56142 35262 56194
rect 41122 56142 41134 56194
rect 41186 56142 41198 56194
rect 55794 56142 55806 56194
rect 55858 56142 55870 56194
rect 26574 56130 26626 56142
rect 43598 56130 43650 56142
rect 17502 56082 17554 56094
rect 22542 56082 22594 56094
rect 25678 56082 25730 56094
rect 28254 56082 28306 56094
rect 7186 56030 7198 56082
rect 7250 56030 7262 56082
rect 12786 56030 12798 56082
rect 12850 56030 12862 56082
rect 18498 56030 18510 56082
rect 18562 56030 18574 56082
rect 24434 56030 24446 56082
rect 24498 56030 24510 56082
rect 27906 56030 27918 56082
rect 27970 56030 27982 56082
rect 17502 56018 17554 56030
rect 22542 56018 22594 56030
rect 25678 56018 25730 56030
rect 28254 56018 28306 56030
rect 28478 56082 28530 56094
rect 28478 56018 28530 56030
rect 34414 56082 34466 56094
rect 39790 56082 39842 56094
rect 36082 56030 36094 56082
rect 36146 56030 36158 56082
rect 42242 56030 42254 56082
rect 42306 56030 42318 56082
rect 46610 56030 46622 56082
rect 46674 56030 46686 56082
rect 52770 56030 52782 56082
rect 52834 56030 52846 56082
rect 54674 56030 54686 56082
rect 54738 56030 54750 56082
rect 34414 56018 34466 56030
rect 39790 56018 39842 56030
rect 4174 55970 4226 55982
rect 3042 55918 3054 55970
rect 3106 55918 3118 55970
rect 4174 55906 4226 55918
rect 5070 55970 5122 55982
rect 5070 55906 5122 55918
rect 6078 55970 6130 55982
rect 6078 55906 6130 55918
rect 6526 55970 6578 55982
rect 8990 55970 9042 55982
rect 7634 55918 7646 55970
rect 7698 55918 7710 55970
rect 6526 55906 6578 55918
rect 8990 55906 9042 55918
rect 9774 55970 9826 55982
rect 9774 55906 9826 55918
rect 10222 55970 10274 55982
rect 10222 55906 10274 55918
rect 10670 55970 10722 55982
rect 10670 55906 10722 55918
rect 11118 55970 11170 55982
rect 13694 55970 13746 55982
rect 12114 55918 12126 55970
rect 12178 55918 12190 55970
rect 11118 55906 11170 55918
rect 13694 55906 13746 55918
rect 14590 55970 14642 55982
rect 14590 55906 14642 55918
rect 15038 55970 15090 55982
rect 15038 55906 15090 55918
rect 15486 55970 15538 55982
rect 15486 55906 15538 55918
rect 15934 55970 15986 55982
rect 15934 55906 15986 55918
rect 16830 55970 16882 55982
rect 16830 55906 16882 55918
rect 17950 55970 18002 55982
rect 20190 55970 20242 55982
rect 19058 55918 19070 55970
rect 19122 55918 19134 55970
rect 17950 55906 18002 55918
rect 20190 55906 20242 55918
rect 20750 55970 20802 55982
rect 20750 55906 20802 55918
rect 21310 55970 21362 55982
rect 21310 55906 21362 55918
rect 22094 55970 22146 55982
rect 25342 55970 25394 55982
rect 23538 55918 23550 55970
rect 23602 55918 23614 55970
rect 22094 55906 22146 55918
rect 25342 55906 25394 55918
rect 28366 55970 28418 55982
rect 31614 55970 31666 55982
rect 29250 55918 29262 55970
rect 29314 55918 29326 55970
rect 28366 55906 28418 55918
rect 31614 55906 31666 55918
rect 32174 55970 32226 55982
rect 32174 55906 32226 55918
rect 33182 55970 33234 55982
rect 33182 55906 33234 55918
rect 33966 55970 34018 55982
rect 33966 55906 34018 55918
rect 36990 55970 37042 55982
rect 36990 55906 37042 55918
rect 37550 55970 37602 55982
rect 37550 55906 37602 55918
rect 37998 55970 38050 55982
rect 37998 55906 38050 55918
rect 40238 55970 40290 55982
rect 40238 55906 40290 55918
rect 43150 55970 43202 55982
rect 43150 55906 43202 55918
rect 46174 55970 46226 55982
rect 47282 55918 47294 55970
rect 47346 55918 47358 55970
rect 53442 55918 53454 55970
rect 53506 55918 53518 55970
rect 46174 55906 46226 55918
rect 22654 55858 22706 55870
rect 14354 55806 14366 55858
rect 14418 55855 14430 55858
rect 15026 55855 15038 55858
rect 14418 55809 15038 55855
rect 14418 55806 14430 55809
rect 15026 55806 15038 55809
rect 15090 55806 15102 55858
rect 15810 55806 15822 55858
rect 15874 55855 15886 55858
rect 16370 55855 16382 55858
rect 15874 55809 16382 55855
rect 15874 55806 15886 55809
rect 16370 55806 16382 55809
rect 16434 55806 16446 55858
rect 20178 55806 20190 55858
rect 20242 55855 20254 55858
rect 20850 55855 20862 55858
rect 20242 55809 20862 55855
rect 20242 55806 20254 55809
rect 20850 55806 20862 55809
rect 20914 55806 20926 55858
rect 30930 55806 30942 55858
rect 30994 55855 31006 55858
rect 31602 55855 31614 55858
rect 30994 55809 31614 55855
rect 30994 55806 31006 55809
rect 31602 55806 31614 55809
rect 31666 55806 31678 55858
rect 22654 55794 22706 55806
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 20290 55470 20302 55522
rect 20354 55519 20366 55522
rect 21074 55519 21086 55522
rect 20354 55473 21086 55519
rect 20354 55470 20366 55473
rect 21074 55470 21086 55473
rect 21138 55470 21150 55522
rect 30370 55470 30382 55522
rect 30434 55519 30446 55522
rect 30930 55519 30942 55522
rect 30434 55473 30942 55519
rect 30434 55470 30446 55473
rect 30930 55470 30942 55473
rect 30994 55470 31006 55522
rect 53890 55470 53902 55522
rect 53954 55519 53966 55522
rect 54674 55519 54686 55522
rect 53954 55473 54686 55519
rect 53954 55470 53966 55473
rect 54674 55470 54686 55473
rect 54738 55470 54750 55522
rect 5854 55410 5906 55422
rect 1922 55358 1934 55410
rect 1986 55358 1998 55410
rect 5854 55346 5906 55358
rect 12910 55410 12962 55422
rect 12910 55346 12962 55358
rect 19854 55410 19906 55422
rect 19854 55346 19906 55358
rect 20302 55410 20354 55422
rect 20302 55346 20354 55358
rect 25790 55410 25842 55422
rect 25790 55346 25842 55358
rect 28478 55410 28530 55422
rect 28478 55346 28530 55358
rect 30606 55410 30658 55422
rect 30606 55346 30658 55358
rect 32958 55410 33010 55422
rect 32958 55346 33010 55358
rect 36542 55410 36594 55422
rect 36542 55346 36594 55358
rect 37886 55410 37938 55422
rect 44606 55410 44658 55422
rect 38882 55358 38894 55410
rect 38946 55358 38958 55410
rect 45826 55358 45838 55410
rect 45890 55358 45902 55410
rect 56018 55358 56030 55410
rect 56082 55358 56094 55410
rect 37886 55346 37938 55358
rect 44606 55346 44658 55358
rect 7534 55298 7586 55310
rect 2818 55246 2830 55298
rect 2882 55246 2894 55298
rect 7534 55234 7586 55246
rect 15038 55298 15090 55310
rect 15038 55234 15090 55246
rect 15150 55298 15202 55310
rect 24894 55298 24946 55310
rect 15250 55246 15262 55298
rect 15314 55246 15326 55298
rect 19170 55246 19182 55298
rect 19234 55246 19246 55298
rect 22082 55246 22094 55298
rect 22146 55246 22158 55298
rect 24210 55246 24222 55298
rect 24274 55246 24286 55298
rect 15150 55234 15202 55246
rect 24894 55234 24946 55246
rect 25230 55298 25282 55310
rect 25230 55234 25282 55246
rect 28030 55298 28082 55310
rect 28030 55234 28082 55246
rect 28254 55298 28306 55310
rect 28254 55234 28306 55246
rect 29934 55298 29986 55310
rect 29934 55234 29986 55246
rect 34302 55298 34354 55310
rect 34302 55234 34354 55246
rect 39342 55298 39394 55310
rect 39342 55234 39394 55246
rect 40014 55298 40066 55310
rect 43374 55298 43426 55310
rect 43138 55246 43150 55298
rect 43202 55246 43214 55298
rect 40014 55234 40066 55246
rect 43374 55234 43426 55246
rect 44046 55298 44098 55310
rect 44046 55234 44098 55246
rect 44494 55298 44546 55310
rect 45714 55246 45726 55298
rect 45778 55246 45790 55298
rect 54898 55246 54910 55298
rect 54962 55246 54974 55298
rect 44494 55234 44546 55246
rect 5070 55186 5122 55198
rect 5070 55122 5122 55134
rect 7198 55186 7250 55198
rect 7198 55122 7250 55134
rect 9438 55186 9490 55198
rect 9438 55122 9490 55134
rect 12126 55186 12178 55198
rect 12126 55122 12178 55134
rect 12574 55186 12626 55198
rect 12574 55122 12626 55134
rect 14702 55186 14754 55198
rect 14702 55122 14754 55134
rect 16270 55186 16322 55198
rect 16270 55122 16322 55134
rect 16606 55186 16658 55198
rect 16606 55122 16658 55134
rect 17166 55186 17218 55198
rect 17166 55122 17218 55134
rect 17278 55186 17330 55198
rect 17278 55122 17330 55134
rect 18174 55186 18226 55198
rect 18174 55122 18226 55134
rect 23102 55186 23154 55198
rect 23102 55122 23154 55134
rect 26238 55186 26290 55198
rect 26238 55122 26290 55134
rect 30158 55186 30210 55198
rect 30158 55122 30210 55134
rect 31166 55186 31218 55198
rect 31166 55122 31218 55134
rect 35758 55186 35810 55198
rect 35758 55122 35810 55134
rect 36094 55186 36146 55198
rect 36094 55122 36146 55134
rect 38558 55186 38610 55198
rect 38558 55122 38610 55134
rect 41134 55186 41186 55198
rect 41134 55122 41186 55134
rect 42478 55186 42530 55198
rect 42478 55122 42530 55134
rect 46622 55186 46674 55198
rect 46622 55122 46674 55134
rect 47182 55186 47234 55198
rect 47182 55122 47234 55134
rect 47518 55186 47570 55198
rect 47518 55122 47570 55134
rect 3726 55074 3778 55086
rect 3726 55010 3778 55022
rect 4174 55074 4226 55086
rect 4174 55010 4226 55022
rect 4622 55074 4674 55086
rect 4622 55010 4674 55022
rect 6302 55074 6354 55086
rect 6302 55010 6354 55022
rect 6750 55074 6802 55086
rect 6750 55010 6802 55022
rect 8094 55074 8146 55086
rect 8094 55010 8146 55022
rect 8542 55074 8594 55086
rect 8542 55010 8594 55022
rect 8878 55074 8930 55086
rect 10670 55074 10722 55086
rect 11678 55074 11730 55086
rect 9762 55022 9774 55074
rect 9826 55022 9838 55074
rect 10994 55022 11006 55074
rect 11058 55022 11070 55074
rect 8878 55010 8930 55022
rect 10670 55010 10722 55022
rect 11678 55010 11730 55022
rect 13694 55074 13746 55086
rect 13694 55010 13746 55022
rect 14142 55074 14194 55086
rect 17502 55074 17554 55086
rect 15138 55022 15150 55074
rect 15202 55022 15214 55074
rect 14142 55010 14194 55022
rect 17502 55010 17554 55022
rect 18286 55074 18338 55086
rect 18286 55010 18338 55022
rect 18398 55074 18450 55086
rect 18398 55010 18450 55022
rect 19406 55074 19458 55086
rect 19406 55010 19458 55022
rect 20862 55074 20914 55086
rect 20862 55010 20914 55022
rect 22318 55074 22370 55086
rect 22318 55010 22370 55022
rect 23214 55074 23266 55086
rect 23214 55010 23266 55022
rect 23326 55074 23378 55086
rect 23326 55010 23378 55022
rect 23998 55074 24050 55086
rect 23998 55010 24050 55022
rect 25006 55074 25058 55086
rect 25006 55010 25058 55022
rect 25678 55074 25730 55086
rect 25678 55010 25730 55022
rect 26686 55074 26738 55086
rect 26686 55010 26738 55022
rect 27134 55074 27186 55086
rect 27134 55010 27186 55022
rect 28926 55074 28978 55086
rect 28926 55010 28978 55022
rect 29710 55074 29762 55086
rect 29710 55010 29762 55022
rect 30046 55074 30098 55086
rect 30046 55010 30098 55022
rect 31390 55074 31442 55086
rect 31390 55010 31442 55022
rect 31614 55074 31666 55086
rect 31614 55010 31666 55022
rect 31726 55074 31778 55086
rect 31726 55010 31778 55022
rect 32174 55074 32226 55086
rect 32174 55010 32226 55022
rect 32622 55074 32674 55086
rect 32622 55010 32674 55022
rect 33406 55074 33458 55086
rect 33406 55010 33458 55022
rect 33966 55074 34018 55086
rect 33966 55010 34018 55022
rect 34862 55074 34914 55086
rect 37438 55074 37490 55086
rect 35186 55022 35198 55074
rect 35250 55022 35262 55074
rect 34862 55010 34914 55022
rect 37438 55010 37490 55022
rect 38782 55074 38834 55086
rect 38782 55010 38834 55022
rect 39790 55074 39842 55086
rect 39790 55010 39842 55022
rect 39902 55074 39954 55086
rect 39902 55010 39954 55022
rect 40462 55074 40514 55086
rect 40462 55010 40514 55022
rect 41246 55074 41298 55086
rect 41246 55010 41298 55022
rect 41470 55074 41522 55086
rect 41470 55010 41522 55022
rect 41918 55074 41970 55086
rect 41918 55010 41970 55022
rect 44718 55074 44770 55086
rect 44718 55010 44770 55022
rect 53902 55074 53954 55086
rect 53902 55010 53954 55022
rect 54350 55074 54402 55086
rect 54350 55010 54402 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 5182 54738 5234 54750
rect 5182 54674 5234 54686
rect 7422 54738 7474 54750
rect 7422 54674 7474 54686
rect 8654 54738 8706 54750
rect 8654 54674 8706 54686
rect 13918 54738 13970 54750
rect 13918 54674 13970 54686
rect 19070 54738 19122 54750
rect 19070 54674 19122 54686
rect 20414 54738 20466 54750
rect 20414 54674 20466 54686
rect 20526 54738 20578 54750
rect 20526 54674 20578 54686
rect 22094 54738 22146 54750
rect 22094 54674 22146 54686
rect 23550 54738 23602 54750
rect 23550 54674 23602 54686
rect 23662 54738 23714 54750
rect 23662 54674 23714 54686
rect 25790 54738 25842 54750
rect 25790 54674 25842 54686
rect 26350 54738 26402 54750
rect 26350 54674 26402 54686
rect 30718 54738 30770 54750
rect 30718 54674 30770 54686
rect 30942 54738 30994 54750
rect 36990 54738 37042 54750
rect 36194 54686 36206 54738
rect 36258 54686 36270 54738
rect 30942 54674 30994 54686
rect 36990 54674 37042 54686
rect 40798 54738 40850 54750
rect 40798 54674 40850 54686
rect 45838 54738 45890 54750
rect 45838 54674 45890 54686
rect 9886 54626 9938 54638
rect 9886 54562 9938 54574
rect 10334 54626 10386 54638
rect 10334 54562 10386 54574
rect 10446 54626 10498 54638
rect 24446 54626 24498 54638
rect 12450 54574 12462 54626
rect 12514 54574 12526 54626
rect 12786 54574 12798 54626
rect 12850 54574 12862 54626
rect 14802 54574 14814 54626
rect 14866 54574 14878 54626
rect 10446 54562 10498 54574
rect 24446 54562 24498 54574
rect 24558 54626 24610 54638
rect 24558 54562 24610 54574
rect 26574 54626 26626 54638
rect 27694 54626 27746 54638
rect 37774 54626 37826 54638
rect 26898 54574 26910 54626
rect 26962 54574 26974 54626
rect 27906 54574 27918 54626
rect 27970 54574 27982 54626
rect 34402 54574 34414 54626
rect 34466 54574 34478 54626
rect 26574 54562 26626 54574
rect 27694 54562 27746 54574
rect 37774 54562 37826 54574
rect 42926 54626 42978 54638
rect 42926 54562 42978 54574
rect 43598 54626 43650 54638
rect 43598 54562 43650 54574
rect 43710 54626 43762 54638
rect 43710 54562 43762 54574
rect 44158 54626 44210 54638
rect 44158 54562 44210 54574
rect 8430 54514 8482 54526
rect 8430 54450 8482 54462
rect 9102 54514 9154 54526
rect 9102 54450 9154 54462
rect 10222 54514 10274 54526
rect 15598 54514 15650 54526
rect 16158 54514 16210 54526
rect 10994 54462 11006 54514
rect 11058 54462 11070 54514
rect 12226 54462 12238 54514
rect 12290 54462 12302 54514
rect 13122 54462 13134 54514
rect 13186 54462 13198 54514
rect 14914 54462 14926 54514
rect 14978 54462 14990 54514
rect 15922 54462 15934 54514
rect 15986 54462 15998 54514
rect 10222 54450 10274 54462
rect 15598 54450 15650 54462
rect 16158 54450 16210 54462
rect 16494 54514 16546 54526
rect 16494 54450 16546 54462
rect 16606 54514 16658 54526
rect 16606 54450 16658 54462
rect 17726 54514 17778 54526
rect 17726 54450 17778 54462
rect 18174 54514 18226 54526
rect 18174 54450 18226 54462
rect 20638 54514 20690 54526
rect 21086 54514 21138 54526
rect 20738 54462 20750 54514
rect 20802 54462 20814 54514
rect 20638 54450 20690 54462
rect 21086 54450 21138 54462
rect 21646 54514 21698 54526
rect 21646 54450 21698 54462
rect 21870 54514 21922 54526
rect 21870 54450 21922 54462
rect 24782 54514 24834 54526
rect 28702 54514 28754 54526
rect 30606 54514 30658 54526
rect 26786 54462 26798 54514
rect 26850 54462 26862 54514
rect 28018 54462 28030 54514
rect 28082 54462 28094 54514
rect 29138 54462 29150 54514
rect 29202 54462 29214 54514
rect 24782 54450 24834 54462
rect 28702 54450 28754 54462
rect 30606 54450 30658 54462
rect 31166 54514 31218 54526
rect 36878 54514 36930 54526
rect 32610 54462 32622 54514
rect 32674 54462 32686 54514
rect 35634 54462 35646 54514
rect 35698 54462 35710 54514
rect 31166 54450 31218 54462
rect 36878 54450 36930 54462
rect 38446 54514 38498 54526
rect 39342 54514 39394 54526
rect 38770 54462 38782 54514
rect 38834 54462 38846 54514
rect 38446 54450 38498 54462
rect 39342 54450 39394 54462
rect 40126 54514 40178 54526
rect 40126 54450 40178 54462
rect 40350 54514 40402 54526
rect 46174 54514 46226 54526
rect 42018 54462 42030 54514
rect 42082 54462 42094 54514
rect 40350 54450 40402 54462
rect 46174 54450 46226 54462
rect 2046 54402 2098 54414
rect 2046 54338 2098 54350
rect 2494 54402 2546 54414
rect 2494 54338 2546 54350
rect 2942 54402 2994 54414
rect 2942 54338 2994 54350
rect 3390 54402 3442 54414
rect 3390 54338 3442 54350
rect 3838 54402 3890 54414
rect 3838 54338 3890 54350
rect 4174 54402 4226 54414
rect 4174 54338 4226 54350
rect 4734 54402 4786 54414
rect 4734 54338 4786 54350
rect 5630 54402 5682 54414
rect 5630 54338 5682 54350
rect 6078 54402 6130 54414
rect 6078 54338 6130 54350
rect 6526 54402 6578 54414
rect 6526 54338 6578 54350
rect 6974 54402 7026 54414
rect 6974 54338 7026 54350
rect 7982 54402 8034 54414
rect 7982 54338 8034 54350
rect 8542 54402 8594 54414
rect 16382 54402 16434 54414
rect 12674 54350 12686 54402
rect 12738 54350 12750 54402
rect 8542 54338 8594 54350
rect 16382 54338 16434 54350
rect 19742 54402 19794 54414
rect 19742 54338 19794 54350
rect 21758 54402 21810 54414
rect 21758 54338 21810 54350
rect 22766 54402 22818 54414
rect 29934 54402 29986 54414
rect 26674 54350 26686 54402
rect 26738 54350 26750 54402
rect 22766 54338 22818 54350
rect 29934 54338 29986 54350
rect 31278 54402 31330 54414
rect 31278 54338 31330 54350
rect 31838 54402 31890 54414
rect 33518 54402 33570 54414
rect 37662 54402 37714 54414
rect 31938 54350 31950 54402
rect 32002 54350 32014 54402
rect 34178 54350 34190 54402
rect 34242 54350 34254 54402
rect 31838 54338 31890 54350
rect 33518 54338 33570 54350
rect 37662 54338 37714 54350
rect 39902 54402 39954 54414
rect 42130 54350 42142 54402
rect 42194 54350 42206 54402
rect 39902 54338 39954 54350
rect 14254 54290 14306 54302
rect 4050 54238 4062 54290
rect 4114 54287 4126 54290
rect 4610 54287 4622 54290
rect 4114 54241 4622 54287
rect 4114 54238 4126 54241
rect 4610 54238 4622 54241
rect 4674 54238 4686 54290
rect 14254 54226 14306 54238
rect 17950 54290 18002 54302
rect 17950 54226 18002 54238
rect 18398 54290 18450 54302
rect 18398 54226 18450 54238
rect 18622 54290 18674 54302
rect 18622 54226 18674 54238
rect 18846 54290 18898 54302
rect 18846 54226 18898 54238
rect 23438 54290 23490 54302
rect 23438 54226 23490 54238
rect 36990 54290 37042 54302
rect 36990 54226 37042 54238
rect 43598 54290 43650 54302
rect 43598 54226 43650 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 9438 53954 9490 53966
rect 22206 53954 22258 53966
rect 20514 53902 20526 53954
rect 20578 53902 20590 53954
rect 9438 53890 9490 53902
rect 22206 53890 22258 53902
rect 28254 53954 28306 53966
rect 28254 53890 28306 53902
rect 28478 53954 28530 53966
rect 28478 53890 28530 53902
rect 28926 53954 28978 53966
rect 28926 53890 28978 53902
rect 30494 53954 30546 53966
rect 30494 53890 30546 53902
rect 34190 53954 34242 53966
rect 34190 53890 34242 53902
rect 39454 53954 39506 53966
rect 39454 53890 39506 53902
rect 39566 53954 39618 53966
rect 39566 53890 39618 53902
rect 42702 53954 42754 53966
rect 42702 53890 42754 53902
rect 42926 53954 42978 53966
rect 42926 53890 42978 53902
rect 5070 53842 5122 53854
rect 5070 53778 5122 53790
rect 9102 53842 9154 53854
rect 9102 53778 9154 53790
rect 25454 53842 25506 53854
rect 25454 53778 25506 53790
rect 28030 53842 28082 53854
rect 28030 53778 28082 53790
rect 30830 53842 30882 53854
rect 33406 53842 33458 53854
rect 37550 53842 37602 53854
rect 32050 53790 32062 53842
rect 32114 53790 32126 53842
rect 33954 53790 33966 53842
rect 34018 53790 34030 53842
rect 30830 53778 30882 53790
rect 33406 53778 33458 53790
rect 37550 53778 37602 53790
rect 39790 53842 39842 53854
rect 39790 53778 39842 53790
rect 5742 53730 5794 53742
rect 9886 53730 9938 53742
rect 6962 53678 6974 53730
rect 7026 53678 7038 53730
rect 5742 53666 5794 53678
rect 9886 53666 9938 53678
rect 10670 53730 10722 53742
rect 10670 53666 10722 53678
rect 14702 53730 14754 53742
rect 14702 53666 14754 53678
rect 15038 53730 15090 53742
rect 15038 53666 15090 53678
rect 15598 53730 15650 53742
rect 15598 53666 15650 53678
rect 16046 53730 16098 53742
rect 16046 53666 16098 53678
rect 16942 53730 16994 53742
rect 16942 53666 16994 53678
rect 17614 53730 17666 53742
rect 17614 53666 17666 53678
rect 17838 53730 17890 53742
rect 17838 53666 17890 53678
rect 18062 53730 18114 53742
rect 18062 53666 18114 53678
rect 18174 53730 18226 53742
rect 18174 53666 18226 53678
rect 19966 53730 20018 53742
rect 19966 53666 20018 53678
rect 20190 53730 20242 53742
rect 29822 53730 29874 53742
rect 33630 53730 33682 53742
rect 21634 53678 21646 53730
rect 21698 53678 21710 53730
rect 22642 53678 22654 53730
rect 22706 53678 22718 53730
rect 24098 53678 24110 53730
rect 24162 53678 24174 53730
rect 30146 53678 30158 53730
rect 30210 53678 30222 53730
rect 31826 53678 31838 53730
rect 31890 53678 31902 53730
rect 20190 53666 20242 53678
rect 29822 53666 29874 53678
rect 33630 53666 33682 53678
rect 34638 53730 34690 53742
rect 34638 53666 34690 53678
rect 35870 53730 35922 53742
rect 35870 53666 35922 53678
rect 37662 53730 37714 53742
rect 41134 53730 41186 53742
rect 43598 53730 43650 53742
rect 37986 53678 37998 53730
rect 38050 53678 38062 53730
rect 43138 53678 43150 53730
rect 43202 53678 43214 53730
rect 37662 53666 37714 53678
rect 41134 53666 41186 53678
rect 43598 53666 43650 53678
rect 1822 53618 1874 53630
rect 1822 53554 1874 53566
rect 6750 53618 6802 53630
rect 6750 53554 6802 53566
rect 7646 53618 7698 53630
rect 7646 53554 7698 53566
rect 7758 53618 7810 53630
rect 7758 53554 7810 53566
rect 9326 53618 9378 53630
rect 9326 53554 9378 53566
rect 10110 53618 10162 53630
rect 10110 53554 10162 53566
rect 10222 53618 10274 53630
rect 10222 53554 10274 53566
rect 13806 53618 13858 53630
rect 13806 53554 13858 53566
rect 16606 53618 16658 53630
rect 16606 53554 16658 53566
rect 18846 53618 18898 53630
rect 25006 53618 25058 53630
rect 23986 53566 23998 53618
rect 24050 53566 24062 53618
rect 18846 53554 18898 53566
rect 25006 53554 25058 53566
rect 26574 53618 26626 53630
rect 26574 53554 26626 53566
rect 27022 53618 27074 53630
rect 27022 53554 27074 53566
rect 27358 53618 27410 53630
rect 27358 53554 27410 53566
rect 30382 53618 30434 53630
rect 30382 53554 30434 53566
rect 32734 53618 32786 53630
rect 32734 53554 32786 53566
rect 33966 53618 34018 53630
rect 33966 53554 34018 53566
rect 39902 53618 39954 53630
rect 39902 53554 39954 53566
rect 40910 53618 40962 53630
rect 40910 53554 40962 53566
rect 41358 53618 41410 53630
rect 41358 53554 41410 53566
rect 42590 53618 42642 53630
rect 42590 53554 42642 53566
rect 45838 53618 45890 53630
rect 45838 53554 45890 53566
rect 2270 53506 2322 53518
rect 2270 53442 2322 53454
rect 2718 53506 2770 53518
rect 2718 53442 2770 53454
rect 3166 53506 3218 53518
rect 3166 53442 3218 53454
rect 3614 53506 3666 53518
rect 3614 53442 3666 53454
rect 4062 53506 4114 53518
rect 4062 53442 4114 53454
rect 4510 53506 4562 53518
rect 4510 53442 4562 53454
rect 6302 53506 6354 53518
rect 6302 53442 6354 53454
rect 7982 53506 8034 53518
rect 7982 53442 8034 53454
rect 8654 53506 8706 53518
rect 8654 53442 8706 53454
rect 11118 53506 11170 53518
rect 11118 53442 11170 53454
rect 11230 53506 11282 53518
rect 11230 53442 11282 53454
rect 11342 53506 11394 53518
rect 11342 53442 11394 53454
rect 11902 53506 11954 53518
rect 11902 53442 11954 53454
rect 12574 53506 12626 53518
rect 12574 53442 12626 53454
rect 13022 53506 13074 53518
rect 13022 53442 13074 53454
rect 14142 53506 14194 53518
rect 14142 53442 14194 53454
rect 14814 53506 14866 53518
rect 14814 53442 14866 53454
rect 16718 53506 16770 53518
rect 16718 53442 16770 53454
rect 18958 53506 19010 53518
rect 18958 53442 19010 53454
rect 19182 53506 19234 53518
rect 19182 53442 19234 53454
rect 21870 53506 21922 53518
rect 21870 53442 21922 53454
rect 22094 53506 22146 53518
rect 24558 53506 24610 53518
rect 22754 53454 22766 53506
rect 22818 53454 22830 53506
rect 22978 53454 22990 53506
rect 23042 53454 23054 53506
rect 22094 53442 22146 53454
rect 24558 53442 24610 53454
rect 26126 53506 26178 53518
rect 26126 53442 26178 53454
rect 35086 53506 35138 53518
rect 35086 53442 35138 53454
rect 35646 53506 35698 53518
rect 35646 53442 35698 53454
rect 35758 53506 35810 53518
rect 35758 53442 35810 53454
rect 36094 53506 36146 53518
rect 36094 53442 36146 53454
rect 36766 53506 36818 53518
rect 36766 53442 36818 53454
rect 40350 53506 40402 53518
rect 40350 53442 40402 53454
rect 41022 53506 41074 53518
rect 41022 53442 41074 53454
rect 41918 53506 41970 53518
rect 41918 53442 41970 53454
rect 44046 53506 44098 53518
rect 44046 53442 44098 53454
rect 45950 53506 46002 53518
rect 45950 53442 46002 53454
rect 46062 53506 46114 53518
rect 46062 53442 46114 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 3502 53170 3554 53182
rect 3502 53106 3554 53118
rect 4286 53170 4338 53182
rect 4286 53106 4338 53118
rect 5630 53170 5682 53182
rect 5630 53106 5682 53118
rect 6190 53170 6242 53182
rect 6190 53106 6242 53118
rect 6526 53170 6578 53182
rect 6526 53106 6578 53118
rect 9774 53170 9826 53182
rect 9774 53106 9826 53118
rect 10670 53170 10722 53182
rect 10670 53106 10722 53118
rect 10894 53170 10946 53182
rect 10894 53106 10946 53118
rect 17614 53170 17666 53182
rect 17614 53106 17666 53118
rect 18398 53170 18450 53182
rect 18398 53106 18450 53118
rect 20526 53170 20578 53182
rect 23550 53170 23602 53182
rect 22530 53118 22542 53170
rect 22594 53118 22606 53170
rect 20526 53106 20578 53118
rect 23550 53106 23602 53118
rect 26798 53170 26850 53182
rect 26798 53106 26850 53118
rect 31166 53170 31218 53182
rect 31166 53106 31218 53118
rect 33742 53170 33794 53182
rect 33742 53106 33794 53118
rect 36766 53170 36818 53182
rect 36766 53106 36818 53118
rect 37550 53170 37602 53182
rect 37550 53106 37602 53118
rect 39118 53170 39170 53182
rect 39118 53106 39170 53118
rect 39566 53170 39618 53182
rect 39566 53106 39618 53118
rect 40014 53170 40066 53182
rect 40014 53106 40066 53118
rect 43038 53170 43090 53182
rect 43038 53106 43090 53118
rect 7310 53058 7362 53070
rect 26014 53058 26066 53070
rect 12674 53006 12686 53058
rect 12738 53006 12750 53058
rect 13682 53006 13694 53058
rect 13746 53006 13758 53058
rect 21410 53006 21422 53058
rect 21474 53006 21486 53058
rect 7310 52994 7362 53006
rect 26014 52994 26066 53006
rect 26126 53058 26178 53070
rect 26126 52994 26178 53006
rect 27918 53058 27970 53070
rect 27918 52994 27970 53006
rect 35646 53058 35698 53070
rect 35646 52994 35698 53006
rect 35758 53058 35810 53070
rect 35758 52994 35810 53006
rect 36542 53058 36594 53070
rect 36542 52994 36594 53006
rect 38222 53058 38274 53070
rect 38222 52994 38274 53006
rect 40798 53058 40850 53070
rect 40798 52994 40850 53006
rect 42478 53058 42530 53070
rect 42478 52994 42530 53006
rect 43598 53058 43650 53070
rect 43598 52994 43650 53006
rect 43710 53058 43762 53070
rect 43710 52994 43762 53006
rect 7198 52946 7250 52958
rect 7198 52882 7250 52894
rect 8094 52946 8146 52958
rect 8094 52882 8146 52894
rect 11006 52946 11058 52958
rect 13134 52946 13186 52958
rect 14702 52946 14754 52958
rect 21982 52946 22034 52958
rect 11890 52894 11902 52946
rect 11954 52894 11966 52946
rect 12562 52894 12574 52946
rect 12626 52894 12638 52946
rect 13346 52894 13358 52946
rect 13410 52894 13422 52946
rect 21186 52894 21198 52946
rect 21250 52894 21262 52946
rect 11006 52882 11058 52894
rect 13134 52882 13186 52894
rect 14702 52882 14754 52894
rect 21982 52882 22034 52894
rect 22206 52946 22258 52958
rect 22206 52882 22258 52894
rect 26686 52946 26738 52958
rect 26686 52882 26738 52894
rect 26910 52946 26962 52958
rect 26910 52882 26962 52894
rect 27358 52946 27410 52958
rect 27358 52882 27410 52894
rect 27806 52946 27858 52958
rect 35982 52946 36034 52958
rect 30930 52894 30942 52946
rect 30994 52894 31006 52946
rect 33954 52894 33966 52946
rect 34018 52894 34030 52946
rect 27806 52882 27858 52894
rect 35982 52882 36034 52894
rect 36430 52946 36482 52958
rect 36430 52882 36482 52894
rect 37438 52946 37490 52958
rect 41582 52946 41634 52958
rect 37762 52894 37774 52946
rect 37826 52894 37838 52946
rect 37438 52882 37490 52894
rect 41582 52882 41634 52894
rect 41806 52946 41858 52958
rect 42254 52946 42306 52958
rect 42130 52894 42142 52946
rect 42194 52894 42206 52946
rect 41806 52882 41858 52894
rect 42254 52882 42306 52894
rect 43934 52946 43986 52958
rect 44818 52894 44830 52946
rect 44882 52894 44894 52946
rect 45938 52894 45950 52946
rect 46002 52894 46014 52946
rect 43934 52882 43986 52894
rect 2158 52834 2210 52846
rect 2158 52770 2210 52782
rect 2606 52834 2658 52846
rect 2606 52770 2658 52782
rect 2942 52834 2994 52846
rect 2942 52770 2994 52782
rect 3950 52834 4002 52846
rect 3950 52770 4002 52782
rect 4846 52834 4898 52846
rect 4846 52770 4898 52782
rect 5294 52834 5346 52846
rect 5294 52770 5346 52782
rect 8654 52834 8706 52846
rect 8654 52770 8706 52782
rect 9102 52834 9154 52846
rect 9102 52770 9154 52782
rect 10334 52834 10386 52846
rect 10334 52770 10386 52782
rect 14366 52834 14418 52846
rect 14366 52770 14418 52782
rect 15262 52834 15314 52846
rect 15262 52770 15314 52782
rect 15598 52834 15650 52846
rect 15598 52770 15650 52782
rect 16158 52834 16210 52846
rect 16158 52770 16210 52782
rect 16494 52834 16546 52846
rect 16494 52770 16546 52782
rect 16942 52834 16994 52846
rect 16942 52770 16994 52782
rect 18958 52834 19010 52846
rect 18958 52770 19010 52782
rect 19406 52834 19458 52846
rect 19406 52770 19458 52782
rect 20190 52834 20242 52846
rect 20190 52770 20242 52782
rect 23102 52834 23154 52846
rect 23102 52770 23154 52782
rect 24446 52834 24498 52846
rect 24446 52770 24498 52782
rect 24782 52834 24834 52846
rect 24782 52770 24834 52782
rect 28478 52834 28530 52846
rect 28478 52770 28530 52782
rect 28926 52834 28978 52846
rect 28926 52770 28978 52782
rect 29374 52834 29426 52846
rect 29374 52770 29426 52782
rect 29822 52834 29874 52846
rect 29822 52770 29874 52782
rect 30270 52834 30322 52846
rect 30270 52770 30322 52782
rect 31614 52834 31666 52846
rect 31614 52770 31666 52782
rect 32062 52834 32114 52846
rect 32062 52770 32114 52782
rect 32622 52834 32674 52846
rect 32622 52770 32674 52782
rect 34526 52834 34578 52846
rect 34526 52770 34578 52782
rect 35198 52834 35250 52846
rect 35198 52770 35250 52782
rect 38670 52834 38722 52846
rect 42354 52782 42366 52834
rect 42418 52782 42430 52834
rect 44482 52782 44494 52834
rect 44546 52782 44558 52834
rect 38670 52770 38722 52782
rect 7310 52722 7362 52734
rect 26014 52722 26066 52734
rect 2034 52670 2046 52722
rect 2098 52719 2110 52722
rect 3714 52719 3726 52722
rect 2098 52673 3726 52719
rect 2098 52670 2110 52673
rect 3714 52670 3726 52673
rect 3778 52719 3790 52722
rect 4162 52719 4174 52722
rect 3778 52673 4174 52719
rect 3778 52670 3790 52673
rect 4162 52670 4174 52673
rect 4226 52670 4238 52722
rect 18274 52670 18286 52722
rect 18338 52719 18350 52722
rect 19170 52719 19182 52722
rect 18338 52673 19182 52719
rect 18338 52670 18350 52673
rect 19170 52670 19182 52673
rect 19234 52670 19246 52722
rect 7310 52658 7362 52670
rect 26014 52658 26066 52670
rect 27918 52722 27970 52734
rect 33630 52722 33682 52734
rect 28690 52670 28702 52722
rect 28754 52719 28766 52722
rect 29138 52719 29150 52722
rect 28754 52673 29150 52719
rect 28754 52670 28766 52673
rect 29138 52670 29150 52673
rect 29202 52719 29214 52722
rect 29810 52719 29822 52722
rect 29202 52673 29822 52719
rect 29202 52670 29214 52673
rect 29810 52670 29822 52673
rect 29874 52670 29886 52722
rect 46162 52670 46174 52722
rect 46226 52670 46238 52722
rect 27918 52658 27970 52670
rect 33630 52658 33682 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 12014 52386 12066 52398
rect 12014 52322 12066 52334
rect 18286 52386 18338 52398
rect 18286 52322 18338 52334
rect 18510 52386 18562 52398
rect 18510 52322 18562 52334
rect 19406 52386 19458 52398
rect 19406 52322 19458 52334
rect 20078 52386 20130 52398
rect 20078 52322 20130 52334
rect 25230 52386 25282 52398
rect 33070 52386 33122 52398
rect 27458 52334 27470 52386
rect 27522 52334 27534 52386
rect 25230 52322 25282 52334
rect 33070 52322 33122 52334
rect 44718 52386 44770 52398
rect 44718 52322 44770 52334
rect 4510 52274 4562 52286
rect 4510 52210 4562 52222
rect 5854 52274 5906 52286
rect 17502 52274 17554 52286
rect 12898 52222 12910 52274
rect 12962 52222 12974 52274
rect 5854 52210 5906 52222
rect 17502 52210 17554 52222
rect 19182 52274 19234 52286
rect 34414 52274 34466 52286
rect 37550 52274 37602 52286
rect 23538 52222 23550 52274
rect 23602 52222 23614 52274
rect 27122 52222 27134 52274
rect 27186 52222 27198 52274
rect 29810 52222 29822 52274
rect 29874 52222 29886 52274
rect 35522 52222 35534 52274
rect 35586 52222 35598 52274
rect 19182 52210 19234 52222
rect 34414 52210 34466 52222
rect 37550 52210 37602 52222
rect 40014 52274 40066 52286
rect 40014 52210 40066 52222
rect 40910 52274 40962 52286
rect 40910 52210 40962 52222
rect 41582 52274 41634 52286
rect 42466 52222 42478 52274
rect 42530 52222 42542 52274
rect 41582 52210 41634 52222
rect 3278 52162 3330 52174
rect 3278 52098 3330 52110
rect 5070 52162 5122 52174
rect 11454 52162 11506 52174
rect 6962 52110 6974 52162
rect 7026 52110 7038 52162
rect 7186 52110 7198 52162
rect 7250 52110 7262 52162
rect 8194 52110 8206 52162
rect 8258 52110 8270 52162
rect 8866 52110 8878 52162
rect 8930 52110 8942 52162
rect 9986 52110 9998 52162
rect 10050 52110 10062 52162
rect 5070 52098 5122 52110
rect 11454 52098 11506 52110
rect 11902 52162 11954 52174
rect 11902 52098 11954 52110
rect 12798 52162 12850 52174
rect 18174 52162 18226 52174
rect 14466 52110 14478 52162
rect 14530 52110 14542 52162
rect 12798 52098 12850 52110
rect 18174 52098 18226 52110
rect 19630 52162 19682 52174
rect 19630 52098 19682 52110
rect 20526 52162 20578 52174
rect 20526 52098 20578 52110
rect 20862 52162 20914 52174
rect 32510 52162 32562 52174
rect 36318 52162 36370 52174
rect 22530 52110 22542 52162
rect 22594 52110 22606 52162
rect 24098 52110 24110 52162
rect 24162 52110 24174 52162
rect 26338 52110 26350 52162
rect 26402 52110 26414 52162
rect 27234 52110 27246 52162
rect 27298 52110 27310 52162
rect 30034 52110 30046 52162
rect 30098 52110 30110 52162
rect 35858 52110 35870 52162
rect 35922 52110 35934 52162
rect 20862 52098 20914 52110
rect 32510 52098 32562 52110
rect 36318 52098 36370 52110
rect 36766 52162 36818 52174
rect 36766 52098 36818 52110
rect 40462 52162 40514 52174
rect 44382 52162 44434 52174
rect 42802 52110 42814 52162
rect 42866 52110 42878 52162
rect 40462 52098 40514 52110
rect 44382 52098 44434 52110
rect 45390 52162 45442 52174
rect 56030 52162 56082 52174
rect 54898 52110 54910 52162
rect 54962 52110 54974 52162
rect 45390 52098 45442 52110
rect 56030 52098 56082 52110
rect 7422 52050 7474 52062
rect 11118 52050 11170 52062
rect 14030 52050 14082 52062
rect 8306 51998 8318 52050
rect 8370 51998 8382 52050
rect 8754 51998 8766 52050
rect 8818 51998 8830 52050
rect 12562 51998 12574 52050
rect 12626 51998 12638 52050
rect 7422 51986 7474 51998
rect 11118 51986 11170 51998
rect 14030 51986 14082 51998
rect 15038 52050 15090 52062
rect 16270 52050 16322 52062
rect 15362 51998 15374 52050
rect 15426 51998 15438 52050
rect 15038 51986 15090 51998
rect 16270 51986 16322 51998
rect 16494 52050 16546 52062
rect 16494 51986 16546 51998
rect 20638 52050 20690 52062
rect 20638 51986 20690 51998
rect 22318 52050 22370 52062
rect 22318 51986 22370 51998
rect 22878 52050 22930 52062
rect 22878 51986 22930 51998
rect 23662 52050 23714 52062
rect 23662 51986 23714 51998
rect 24670 52050 24722 52062
rect 24670 51986 24722 51998
rect 24894 52050 24946 52062
rect 24894 51986 24946 51998
rect 25566 52050 25618 52062
rect 25566 51986 25618 51998
rect 26126 52050 26178 52062
rect 30718 52050 30770 52062
rect 28466 51998 28478 52050
rect 28530 51998 28542 52050
rect 26126 51986 26178 51998
rect 30718 51986 30770 51998
rect 31838 52050 31890 52062
rect 31838 51986 31890 51998
rect 32062 52050 32114 52062
rect 32062 51986 32114 51998
rect 32958 52050 33010 52062
rect 32958 51986 33010 51998
rect 33742 52050 33794 52062
rect 33742 51986 33794 51998
rect 38446 52050 38498 52062
rect 38446 51986 38498 51998
rect 43262 52050 43314 52062
rect 43262 51986 43314 51998
rect 1934 51938 1986 51950
rect 1934 51874 1986 51886
rect 2382 51938 2434 51950
rect 2382 51874 2434 51886
rect 2830 51938 2882 51950
rect 2830 51874 2882 51886
rect 3726 51938 3778 51950
rect 3726 51874 3778 51886
rect 4174 51938 4226 51950
rect 11230 51938 11282 51950
rect 9090 51886 9102 51938
rect 9154 51886 9166 51938
rect 4174 51874 4226 51886
rect 11230 51874 11282 51886
rect 12350 51938 12402 51950
rect 12350 51874 12402 51886
rect 13694 51938 13746 51950
rect 13694 51874 13746 51886
rect 13806 51938 13858 51950
rect 13806 51874 13858 51886
rect 13918 51938 13970 51950
rect 13918 51874 13970 51886
rect 16382 51938 16434 51950
rect 16382 51874 16434 51886
rect 16718 51938 16770 51950
rect 16718 51874 16770 51886
rect 18174 51938 18226 51950
rect 18174 51874 18226 51886
rect 21758 51938 21810 51950
rect 21758 51874 21810 51886
rect 22766 51938 22818 51950
rect 22766 51874 22818 51886
rect 23326 51938 23378 51950
rect 23326 51874 23378 51886
rect 23550 51938 23602 51950
rect 23550 51874 23602 51886
rect 25118 51938 25170 51950
rect 25118 51874 25170 51886
rect 28814 51938 28866 51950
rect 28814 51874 28866 51886
rect 31278 51938 31330 51950
rect 31278 51874 31330 51886
rect 31950 51938 32002 51950
rect 31950 51874 32002 51886
rect 33070 51938 33122 51950
rect 33070 51874 33122 51886
rect 33854 51938 33906 51950
rect 33854 51874 33906 51886
rect 34078 51938 34130 51950
rect 34078 51874 34130 51886
rect 37662 51938 37714 51950
rect 37662 51874 37714 51886
rect 38558 51938 38610 51950
rect 38558 51874 38610 51886
rect 38782 51938 38834 51950
rect 38782 51874 38834 51886
rect 39230 51938 39282 51950
rect 39230 51874 39282 51886
rect 39566 51938 39618 51950
rect 39566 51874 39618 51886
rect 44606 51938 44658 51950
rect 44606 51874 44658 51886
rect 45838 51938 45890 51950
rect 45838 51874 45890 51886
rect 45950 51938 46002 51950
rect 45950 51874 46002 51886
rect 46062 51938 46114 51950
rect 46062 51874 46114 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 1822 51602 1874 51614
rect 1822 51538 1874 51550
rect 2718 51602 2770 51614
rect 2718 51538 2770 51550
rect 5742 51602 5794 51614
rect 6862 51602 6914 51614
rect 8990 51602 9042 51614
rect 6514 51550 6526 51602
rect 6578 51550 6590 51602
rect 8530 51550 8542 51602
rect 8594 51550 8606 51602
rect 5742 51538 5794 51550
rect 6862 51538 6914 51550
rect 8990 51538 9042 51550
rect 9886 51602 9938 51614
rect 9886 51538 9938 51550
rect 14926 51602 14978 51614
rect 14926 51538 14978 51550
rect 17726 51602 17778 51614
rect 17726 51538 17778 51550
rect 17950 51602 18002 51614
rect 17950 51538 18002 51550
rect 19294 51602 19346 51614
rect 20526 51602 20578 51614
rect 20178 51550 20190 51602
rect 20242 51550 20254 51602
rect 19294 51538 19346 51550
rect 20526 51538 20578 51550
rect 21310 51602 21362 51614
rect 21310 51538 21362 51550
rect 22542 51602 22594 51614
rect 22542 51538 22594 51550
rect 23774 51602 23826 51614
rect 23774 51538 23826 51550
rect 24558 51602 24610 51614
rect 24558 51538 24610 51550
rect 31054 51602 31106 51614
rect 40350 51602 40402 51614
rect 34738 51550 34750 51602
rect 34802 51550 34814 51602
rect 35970 51550 35982 51602
rect 36034 51550 36046 51602
rect 39778 51550 39790 51602
rect 39842 51550 39854 51602
rect 31054 51538 31106 51550
rect 40350 51538 40402 51550
rect 41694 51602 41746 51614
rect 41694 51538 41746 51550
rect 48750 51602 48802 51614
rect 48750 51538 48802 51550
rect 5406 51490 5458 51502
rect 4834 51438 4846 51490
rect 4898 51438 4910 51490
rect 5406 51426 5458 51438
rect 7870 51490 7922 51502
rect 7870 51426 7922 51438
rect 7982 51490 8034 51502
rect 7982 51426 8034 51438
rect 8094 51490 8146 51502
rect 8094 51426 8146 51438
rect 12238 51490 12290 51502
rect 12238 51426 12290 51438
rect 16382 51490 16434 51502
rect 16382 51426 16434 51438
rect 16494 51490 16546 51502
rect 16494 51426 16546 51438
rect 23438 51490 23490 51502
rect 23438 51426 23490 51438
rect 23662 51490 23714 51502
rect 23662 51426 23714 51438
rect 24782 51490 24834 51502
rect 24782 51426 24834 51438
rect 25566 51490 25618 51502
rect 25566 51426 25618 51438
rect 26238 51490 26290 51502
rect 30382 51490 30434 51502
rect 36766 51490 36818 51502
rect 28466 51438 28478 51490
rect 28530 51438 28542 51490
rect 31714 51438 31726 51490
rect 31778 51438 31790 51490
rect 33842 51438 33854 51490
rect 33906 51438 33918 51490
rect 26238 51426 26290 51438
rect 30382 51426 30434 51438
rect 36766 51426 36818 51438
rect 38110 51490 38162 51502
rect 38882 51438 38894 51490
rect 38946 51438 38958 51490
rect 43586 51438 43598 51490
rect 43650 51438 43662 51490
rect 44930 51438 44942 51490
rect 44994 51438 45006 51490
rect 38110 51426 38162 51438
rect 9998 51378 10050 51390
rect 4610 51326 4622 51378
rect 4674 51326 4686 51378
rect 9998 51314 10050 51326
rect 10222 51378 10274 51390
rect 11006 51378 11058 51390
rect 10434 51326 10446 51378
rect 10498 51326 10510 51378
rect 10222 51314 10274 51326
rect 11006 51314 11058 51326
rect 11342 51378 11394 51390
rect 11342 51314 11394 51326
rect 11678 51378 11730 51390
rect 11678 51314 11730 51326
rect 12126 51378 12178 51390
rect 12126 51314 12178 51326
rect 12462 51378 12514 51390
rect 12462 51314 12514 51326
rect 12798 51378 12850 51390
rect 16158 51378 16210 51390
rect 17614 51378 17666 51390
rect 18958 51378 19010 51390
rect 13682 51326 13694 51378
rect 13746 51326 13758 51378
rect 15138 51326 15150 51378
rect 15202 51326 15214 51378
rect 16930 51326 16942 51378
rect 16994 51326 17006 51378
rect 18162 51326 18174 51378
rect 18226 51326 18238 51378
rect 12798 51314 12850 51326
rect 16158 51314 16210 51326
rect 17614 51314 17666 51326
rect 18958 51314 19010 51326
rect 19406 51378 19458 51390
rect 19406 51314 19458 51326
rect 19518 51378 19570 51390
rect 19518 51314 19570 51326
rect 22094 51378 22146 51390
rect 22766 51378 22818 51390
rect 22418 51326 22430 51378
rect 22482 51326 22494 51378
rect 22094 51314 22146 51326
rect 22766 51314 22818 51326
rect 23886 51378 23938 51390
rect 23886 51314 23938 51326
rect 23998 51378 24050 51390
rect 23998 51314 24050 51326
rect 24894 51378 24946 51390
rect 30046 51378 30098 51390
rect 35646 51378 35698 51390
rect 44494 51378 44546 51390
rect 48414 51378 48466 51390
rect 26562 51326 26574 51378
rect 26626 51326 26638 51378
rect 27906 51326 27918 51378
rect 27970 51326 27982 51378
rect 28354 51326 28366 51378
rect 28418 51326 28430 51378
rect 31602 51326 31614 51378
rect 31666 51326 31678 51378
rect 33730 51326 33742 51378
rect 33794 51326 33806 51378
rect 34850 51326 34862 51378
rect 34914 51326 34926 51378
rect 38770 51326 38782 51378
rect 38834 51326 38846 51378
rect 39666 51326 39678 51378
rect 39730 51326 39742 51378
rect 42130 51326 42142 51378
rect 42194 51326 42206 51378
rect 42914 51326 42926 51378
rect 42978 51326 42990 51378
rect 44818 51326 44830 51378
rect 44882 51326 44894 51378
rect 45938 51326 45950 51378
rect 46002 51326 46014 51378
rect 24894 51314 24946 51326
rect 30046 51314 30098 51326
rect 35646 51314 35698 51326
rect 44494 51314 44546 51326
rect 48414 51314 48466 51326
rect 2270 51266 2322 51278
rect 2270 51202 2322 51214
rect 3166 51266 3218 51278
rect 3166 51202 3218 51214
rect 3614 51266 3666 51278
rect 3614 51202 3666 51214
rect 4062 51266 4114 51278
rect 4062 51202 4114 51214
rect 10110 51266 10162 51278
rect 11454 51266 11506 51278
rect 14366 51266 14418 51278
rect 21870 51266 21922 51278
rect 27022 51266 27074 51278
rect 29374 51266 29426 51278
rect 10658 51214 10670 51266
rect 10722 51263 10734 51266
rect 10882 51263 10894 51266
rect 10722 51217 10894 51263
rect 10722 51214 10734 51217
rect 10882 51214 10894 51217
rect 10946 51214 10958 51266
rect 13906 51214 13918 51266
rect 13970 51214 13982 51266
rect 16482 51214 16494 51266
rect 16546 51214 16558 51266
rect 22642 51214 22654 51266
rect 22706 51214 22718 51266
rect 28242 51214 28254 51266
rect 28306 51214 28318 51266
rect 10110 51202 10162 51214
rect 11454 51202 11506 51214
rect 14366 51202 14418 51214
rect 21870 51202 21922 51214
rect 27022 51202 27074 51214
rect 29374 51202 29426 51214
rect 35422 51266 35474 51278
rect 35422 51202 35474 51214
rect 37326 51266 37378 51278
rect 40798 51266 40850 51278
rect 47854 51266 47906 51278
rect 38210 51214 38222 51266
rect 38274 51214 38286 51266
rect 42802 51214 42814 51266
rect 42866 51214 42878 51266
rect 45714 51214 45726 51266
rect 45778 51214 45790 51266
rect 37326 51202 37378 51214
rect 40798 51202 40850 51214
rect 47854 51202 47906 51214
rect 26574 51154 26626 51166
rect 3490 51102 3502 51154
rect 3554 51151 3566 51154
rect 4050 51151 4062 51154
rect 3554 51105 4062 51151
rect 3554 51102 3566 51105
rect 4050 51102 4062 51105
rect 4114 51102 4126 51154
rect 26574 51090 26626 51102
rect 32398 51154 32450 51166
rect 32398 51090 32450 51102
rect 32734 51154 32786 51166
rect 32734 51090 32786 51102
rect 36542 51154 36594 51166
rect 36542 51090 36594 51102
rect 36878 51154 36930 51166
rect 36878 51090 36930 51102
rect 37886 51154 37938 51166
rect 37886 51090 37938 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 5854 50818 5906 50830
rect 5854 50754 5906 50766
rect 9662 50818 9714 50830
rect 9662 50754 9714 50766
rect 9998 50818 10050 50830
rect 26574 50818 26626 50830
rect 12450 50766 12462 50818
rect 12514 50766 12526 50818
rect 9998 50754 10050 50766
rect 26574 50754 26626 50766
rect 27246 50818 27298 50830
rect 27246 50754 27298 50766
rect 27918 50818 27970 50830
rect 27918 50754 27970 50766
rect 34190 50818 34242 50830
rect 34190 50754 34242 50766
rect 34526 50818 34578 50830
rect 34526 50754 34578 50766
rect 8206 50706 8258 50718
rect 15710 50706 15762 50718
rect 24446 50706 24498 50718
rect 37438 50706 37490 50718
rect 44158 50706 44210 50718
rect 46510 50706 46562 50718
rect 6626 50654 6638 50706
rect 6690 50654 6702 50706
rect 10994 50654 11006 50706
rect 11058 50654 11070 50706
rect 14242 50654 14254 50706
rect 14306 50654 14318 50706
rect 16034 50654 16046 50706
rect 16098 50654 16110 50706
rect 29922 50654 29934 50706
rect 29986 50654 29998 50706
rect 36082 50654 36094 50706
rect 36146 50654 36158 50706
rect 38098 50654 38110 50706
rect 38162 50654 38174 50706
rect 46050 50654 46062 50706
rect 46114 50654 46126 50706
rect 8206 50642 8258 50654
rect 15710 50642 15762 50654
rect 24446 50642 24498 50654
rect 37438 50642 37490 50654
rect 44158 50642 44210 50654
rect 46510 50642 46562 50654
rect 4622 50594 4674 50606
rect 3042 50542 3054 50594
rect 3106 50542 3118 50594
rect 4386 50542 4398 50594
rect 4450 50542 4462 50594
rect 4622 50530 4674 50542
rect 4846 50594 4898 50606
rect 12014 50594 12066 50606
rect 13918 50594 13970 50606
rect 17726 50594 17778 50606
rect 9986 50542 9998 50594
rect 10050 50542 10062 50594
rect 11330 50542 11342 50594
rect 11394 50542 11406 50594
rect 11554 50542 11566 50594
rect 11618 50542 11630 50594
rect 12226 50542 12238 50594
rect 12290 50542 12302 50594
rect 13682 50542 13694 50594
rect 13746 50542 13758 50594
rect 16146 50542 16158 50594
rect 16210 50542 16222 50594
rect 4846 50530 4898 50542
rect 12014 50530 12066 50542
rect 13918 50530 13970 50542
rect 17726 50530 17778 50542
rect 19182 50594 19234 50606
rect 19182 50530 19234 50542
rect 20078 50594 20130 50606
rect 20078 50530 20130 50542
rect 22318 50594 22370 50606
rect 22318 50530 22370 50542
rect 25790 50594 25842 50606
rect 27470 50594 27522 50606
rect 32398 50594 32450 50606
rect 26226 50542 26238 50594
rect 26290 50542 26302 50594
rect 29810 50542 29822 50594
rect 29874 50542 29886 50594
rect 25790 50530 25842 50542
rect 27470 50530 27522 50542
rect 32398 50530 32450 50542
rect 32734 50594 32786 50606
rect 42254 50594 42306 50606
rect 34514 50542 34526 50594
rect 34578 50542 34590 50594
rect 35522 50542 35534 50594
rect 35586 50542 35598 50594
rect 36194 50542 36206 50594
rect 36258 50542 36270 50594
rect 39554 50542 39566 50594
rect 39618 50542 39630 50594
rect 41570 50542 41582 50594
rect 41634 50542 41646 50594
rect 32734 50530 32786 50542
rect 42254 50530 42306 50542
rect 42478 50594 42530 50606
rect 45826 50542 45838 50594
rect 45890 50542 45902 50594
rect 42478 50530 42530 50542
rect 5966 50482 6018 50494
rect 1922 50430 1934 50482
rect 1986 50430 1998 50482
rect 5966 50418 6018 50430
rect 9102 50482 9154 50494
rect 9102 50418 9154 50430
rect 14142 50482 14194 50494
rect 14142 50418 14194 50430
rect 14254 50482 14306 50494
rect 14254 50418 14306 50430
rect 15262 50482 15314 50494
rect 15262 50418 15314 50430
rect 17390 50482 17442 50494
rect 17390 50418 17442 50430
rect 18286 50482 18338 50494
rect 18286 50418 18338 50430
rect 22878 50482 22930 50494
rect 22878 50418 22930 50430
rect 23774 50482 23826 50494
rect 23774 50418 23826 50430
rect 23886 50482 23938 50494
rect 23886 50418 23938 50430
rect 24894 50482 24946 50494
rect 24894 50418 24946 50430
rect 27806 50482 27858 50494
rect 27806 50418 27858 50430
rect 28030 50482 28082 50494
rect 28030 50418 28082 50430
rect 28478 50482 28530 50494
rect 28478 50418 28530 50430
rect 30718 50482 30770 50494
rect 30718 50418 30770 50430
rect 31166 50482 31218 50494
rect 31166 50418 31218 50430
rect 32062 50482 32114 50494
rect 32062 50418 32114 50430
rect 33406 50482 33458 50494
rect 33406 50418 33458 50430
rect 35086 50482 35138 50494
rect 40238 50482 40290 50494
rect 36530 50430 36542 50482
rect 36594 50430 36606 50482
rect 38322 50430 38334 50482
rect 38386 50430 38398 50482
rect 35086 50418 35138 50430
rect 40238 50418 40290 50430
rect 3950 50370 4002 50382
rect 3950 50306 4002 50318
rect 4510 50370 4562 50382
rect 4510 50306 4562 50318
rect 5854 50370 5906 50382
rect 5854 50306 5906 50318
rect 7086 50370 7138 50382
rect 7086 50306 7138 50318
rect 7870 50370 7922 50382
rect 7870 50306 7922 50318
rect 8654 50370 8706 50382
rect 8654 50306 8706 50318
rect 18622 50370 18674 50382
rect 18622 50306 18674 50318
rect 19518 50370 19570 50382
rect 19518 50306 19570 50318
rect 20190 50370 20242 50382
rect 20190 50306 20242 50318
rect 20414 50370 20466 50382
rect 20414 50306 20466 50318
rect 20862 50370 20914 50382
rect 20862 50306 20914 50318
rect 21982 50370 22034 50382
rect 21982 50306 22034 50318
rect 23214 50370 23266 50382
rect 23214 50306 23266 50318
rect 24110 50370 24162 50382
rect 24110 50306 24162 50318
rect 26462 50370 26514 50382
rect 26462 50306 26514 50318
rect 32510 50370 32562 50382
rect 32510 50306 32562 50318
rect 40798 50370 40850 50382
rect 40798 50306 40850 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 1934 50034 1986 50046
rect 1934 49970 1986 49982
rect 2382 50034 2434 50046
rect 2382 49970 2434 49982
rect 4062 50034 4114 50046
rect 4062 49970 4114 49982
rect 5854 50034 5906 50046
rect 12350 50034 12402 50046
rect 16046 50034 16098 50046
rect 10994 49982 11006 50034
rect 11058 49982 11070 50034
rect 13234 49982 13246 50034
rect 13298 49982 13310 50034
rect 5854 49970 5906 49982
rect 12350 49970 12402 49982
rect 16046 49970 16098 49982
rect 16718 50034 16770 50046
rect 16718 49970 16770 49982
rect 19854 50034 19906 50046
rect 19854 49970 19906 49982
rect 19966 50034 20018 50046
rect 19966 49970 20018 49982
rect 21758 50034 21810 50046
rect 21758 49970 21810 49982
rect 22318 50034 22370 50046
rect 22318 49970 22370 49982
rect 23326 50034 23378 50046
rect 23326 49970 23378 49982
rect 26014 50034 26066 50046
rect 28030 50034 28082 50046
rect 27234 49982 27246 50034
rect 27298 49982 27310 50034
rect 26014 49970 26066 49982
rect 28030 49970 28082 49982
rect 28366 50034 28418 50046
rect 28366 49970 28418 49982
rect 29374 50034 29426 50046
rect 29374 49970 29426 49982
rect 31278 50034 31330 50046
rect 31278 49970 31330 49982
rect 31950 50034 32002 50046
rect 31950 49970 32002 49982
rect 32622 50034 32674 50046
rect 37886 50034 37938 50046
rect 36530 49982 36542 50034
rect 36594 49982 36606 50034
rect 32622 49970 32674 49982
rect 37886 49970 37938 49982
rect 39118 50034 39170 50046
rect 39118 49970 39170 49982
rect 39566 50034 39618 50046
rect 39566 49970 39618 49982
rect 40574 50034 40626 50046
rect 40574 49970 40626 49982
rect 41918 50034 41970 50046
rect 41918 49970 41970 49982
rect 42142 50034 42194 50046
rect 42142 49970 42194 49982
rect 45054 50034 45106 50046
rect 45054 49970 45106 49982
rect 15934 49922 15986 49934
rect 3154 49870 3166 49922
rect 3218 49870 3230 49922
rect 11890 49870 11902 49922
rect 11954 49870 11966 49922
rect 15934 49858 15986 49870
rect 16942 49922 16994 49934
rect 16942 49858 16994 49870
rect 23214 49922 23266 49934
rect 23214 49858 23266 49870
rect 24222 49922 24274 49934
rect 24222 49858 24274 49870
rect 24334 49922 24386 49934
rect 24334 49858 24386 49870
rect 24894 49922 24946 49934
rect 24894 49858 24946 49870
rect 27806 49922 27858 49934
rect 27806 49858 27858 49870
rect 32062 49922 32114 49934
rect 32062 49858 32114 49870
rect 41806 49922 41858 49934
rect 41806 49858 41858 49870
rect 42478 49922 42530 49934
rect 42478 49858 42530 49870
rect 2830 49810 2882 49822
rect 2830 49746 2882 49758
rect 3726 49810 3778 49822
rect 3726 49746 3778 49758
rect 4062 49810 4114 49822
rect 4062 49746 4114 49758
rect 4286 49810 4338 49822
rect 7086 49810 7138 49822
rect 8654 49810 8706 49822
rect 6850 49758 6862 49810
rect 6914 49758 6926 49810
rect 7522 49758 7534 49810
rect 7586 49758 7598 49810
rect 8082 49758 8094 49810
rect 8146 49758 8158 49810
rect 4286 49746 4338 49758
rect 7086 49746 7138 49758
rect 8654 49746 8706 49758
rect 11566 49810 11618 49822
rect 11566 49746 11618 49758
rect 12910 49810 12962 49822
rect 16382 49810 16434 49822
rect 15474 49758 15486 49810
rect 15538 49758 15550 49810
rect 15698 49758 15710 49810
rect 15762 49758 15774 49810
rect 12910 49746 12962 49758
rect 16382 49746 16434 49758
rect 20078 49810 20130 49822
rect 22654 49810 22706 49822
rect 21522 49758 21534 49810
rect 21586 49758 21598 49810
rect 20078 49746 20130 49758
rect 22654 49746 22706 49758
rect 24558 49810 24610 49822
rect 24558 49746 24610 49758
rect 28254 49810 28306 49822
rect 40126 49810 40178 49822
rect 36754 49758 36766 49810
rect 36818 49758 36830 49810
rect 28254 49746 28306 49758
rect 40126 49746 40178 49758
rect 40350 49810 40402 49822
rect 40350 49746 40402 49758
rect 44718 49810 44770 49822
rect 44718 49746 44770 49758
rect 45166 49810 45218 49822
rect 45166 49746 45218 49758
rect 45390 49810 45442 49822
rect 45390 49746 45442 49758
rect 5070 49698 5122 49710
rect 5070 49634 5122 49646
rect 5406 49698 5458 49710
rect 5406 49634 5458 49646
rect 9998 49698 10050 49710
rect 9998 49634 10050 49646
rect 10446 49698 10498 49710
rect 10446 49634 10498 49646
rect 10670 49698 10722 49710
rect 10670 49634 10722 49646
rect 14030 49698 14082 49710
rect 14030 49634 14082 49646
rect 14478 49698 14530 49710
rect 14478 49634 14530 49646
rect 14926 49698 14978 49710
rect 14926 49634 14978 49646
rect 17614 49698 17666 49710
rect 17614 49634 17666 49646
rect 18398 49698 18450 49710
rect 18398 49634 18450 49646
rect 18846 49698 18898 49710
rect 18846 49634 18898 49646
rect 19630 49698 19682 49710
rect 19630 49634 19682 49646
rect 20862 49698 20914 49710
rect 20862 49634 20914 49646
rect 25566 49698 25618 49710
rect 25566 49634 25618 49646
rect 26686 49698 26738 49710
rect 28926 49698 28978 49710
rect 28354 49646 28366 49698
rect 28418 49646 28430 49698
rect 26686 49634 26738 49646
rect 28926 49634 28978 49646
rect 29822 49698 29874 49710
rect 29822 49634 29874 49646
rect 30270 49698 30322 49710
rect 30270 49634 30322 49646
rect 30718 49698 30770 49710
rect 30718 49634 30770 49646
rect 31838 49698 31890 49710
rect 31838 49634 31890 49646
rect 33518 49698 33570 49710
rect 33518 49634 33570 49646
rect 33966 49698 34018 49710
rect 33966 49634 34018 49646
rect 34750 49698 34802 49710
rect 34750 49634 34802 49646
rect 35198 49698 35250 49710
rect 35198 49634 35250 49646
rect 35646 49698 35698 49710
rect 35646 49634 35698 49646
rect 37326 49698 37378 49710
rect 37326 49634 37378 49646
rect 38222 49698 38274 49710
rect 38222 49634 38274 49646
rect 38670 49698 38722 49710
rect 38670 49634 38722 49646
rect 40238 49698 40290 49710
rect 40238 49634 40290 49646
rect 43486 49698 43538 49710
rect 43486 49634 43538 49646
rect 17054 49586 17106 49598
rect 6962 49534 6974 49586
rect 7026 49534 7038 49586
rect 14578 49534 14590 49586
rect 14642 49583 14654 49586
rect 14914 49583 14926 49586
rect 14642 49537 14926 49583
rect 14642 49534 14654 49537
rect 14914 49534 14926 49537
rect 14978 49534 14990 49586
rect 17054 49522 17106 49534
rect 19406 49586 19458 49598
rect 19406 49522 19458 49534
rect 23326 49586 23378 49598
rect 23326 49522 23378 49534
rect 26910 49586 26962 49598
rect 43598 49586 43650 49598
rect 30258 49534 30270 49586
rect 30322 49583 30334 49586
rect 31042 49583 31054 49586
rect 30322 49537 31054 49583
rect 30322 49534 30334 49537
rect 31042 49534 31054 49537
rect 31106 49534 31118 49586
rect 26910 49522 26962 49534
rect 43598 49522 43650 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 4846 49250 4898 49262
rect 4846 49186 4898 49198
rect 11566 49250 11618 49262
rect 11566 49186 11618 49198
rect 13918 49250 13970 49262
rect 13918 49186 13970 49198
rect 14254 49250 14306 49262
rect 23214 49250 23266 49262
rect 32398 49250 32450 49262
rect 21410 49198 21422 49250
rect 21474 49247 21486 49250
rect 22194 49247 22206 49250
rect 21474 49201 22206 49247
rect 21474 49198 21486 49201
rect 22194 49198 22206 49201
rect 22258 49198 22270 49250
rect 25330 49198 25342 49250
rect 25394 49247 25406 49250
rect 25890 49247 25902 49250
rect 25394 49201 25902 49247
rect 25394 49198 25406 49201
rect 25890 49198 25902 49201
rect 25954 49198 25966 49250
rect 14254 49186 14306 49198
rect 23214 49186 23266 49198
rect 32398 49186 32450 49198
rect 40686 49250 40738 49262
rect 40686 49186 40738 49198
rect 3726 49138 3778 49150
rect 3726 49074 3778 49086
rect 5966 49138 6018 49150
rect 8990 49138 9042 49150
rect 7970 49086 7982 49138
rect 8034 49086 8046 49138
rect 5966 49074 6018 49086
rect 8990 49074 9042 49086
rect 12910 49138 12962 49150
rect 12910 49074 12962 49086
rect 16942 49138 16994 49150
rect 16942 49074 16994 49086
rect 18622 49138 18674 49150
rect 18622 49074 18674 49086
rect 19854 49138 19906 49150
rect 19854 49074 19906 49086
rect 24110 49138 24162 49150
rect 24110 49074 24162 49086
rect 24558 49138 24610 49150
rect 24558 49074 24610 49086
rect 25118 49138 25170 49150
rect 25118 49074 25170 49086
rect 25902 49138 25954 49150
rect 25902 49074 25954 49086
rect 27694 49138 27746 49150
rect 27694 49074 27746 49086
rect 28254 49138 28306 49150
rect 33854 49138 33906 49150
rect 33618 49086 33630 49138
rect 33682 49086 33694 49138
rect 28254 49074 28306 49086
rect 33854 49074 33906 49086
rect 36318 49138 36370 49150
rect 46610 49086 46622 49138
rect 46674 49086 46686 49138
rect 36318 49074 36370 49086
rect 2718 49026 2770 49038
rect 2718 48962 2770 48974
rect 6526 49026 6578 49038
rect 9438 49026 9490 49038
rect 6962 48974 6974 49026
rect 7026 48974 7038 49026
rect 7634 48974 7646 49026
rect 7698 48974 7710 49026
rect 6526 48962 6578 48974
rect 9438 48962 9490 48974
rect 13806 49026 13858 49038
rect 13806 48962 13858 48974
rect 14142 49026 14194 49038
rect 19070 49026 19122 49038
rect 16146 48974 16158 49026
rect 16210 48974 16222 49026
rect 17378 48974 17390 49026
rect 17442 48974 17454 49026
rect 18274 48974 18286 49026
rect 18338 48974 18350 49026
rect 18834 48974 18846 49026
rect 18898 48974 18910 49026
rect 14142 48962 14194 48974
rect 19070 48962 19122 48974
rect 19742 49026 19794 49038
rect 19742 48962 19794 48974
rect 23326 49026 23378 49038
rect 23326 48962 23378 48974
rect 23550 49026 23602 49038
rect 30606 49026 30658 49038
rect 37774 49026 37826 49038
rect 40238 49026 40290 49038
rect 30146 48974 30158 49026
rect 30210 48974 30222 49026
rect 33058 48974 33070 49026
rect 33122 48974 33134 49026
rect 34178 48974 34190 49026
rect 34242 48974 34254 49026
rect 38210 48974 38222 49026
rect 38274 48974 38286 49026
rect 23550 48962 23602 48974
rect 30606 48962 30658 48974
rect 37774 48962 37826 48974
rect 40238 48962 40290 48974
rect 40462 49026 40514 49038
rect 40462 48962 40514 48974
rect 43710 49026 43762 49038
rect 43710 48962 43762 48974
rect 43934 49026 43986 49038
rect 46498 48974 46510 49026
rect 46562 48974 46574 49026
rect 43934 48962 43986 48974
rect 1822 48914 1874 48926
rect 1822 48850 1874 48862
rect 4062 48914 4114 48926
rect 4062 48850 4114 48862
rect 4734 48914 4786 48926
rect 4734 48850 4786 48862
rect 4846 48914 4898 48926
rect 10558 48914 10610 48926
rect 11566 48914 11618 48926
rect 7970 48862 7982 48914
rect 8034 48862 8046 48914
rect 9762 48862 9774 48914
rect 9826 48862 9838 48914
rect 10882 48862 10894 48914
rect 10946 48862 10958 48914
rect 4846 48850 4898 48862
rect 10558 48850 10610 48862
rect 11566 48850 11618 48862
rect 11678 48914 11730 48926
rect 19966 48914 20018 48926
rect 16258 48862 16270 48914
rect 16322 48862 16334 48914
rect 16930 48862 16942 48914
rect 16994 48862 17006 48914
rect 11678 48850 11730 48862
rect 19966 48850 20018 48862
rect 26910 48914 26962 48926
rect 26910 48850 26962 48862
rect 27246 48914 27298 48926
rect 31502 48914 31554 48926
rect 29810 48862 29822 48914
rect 29874 48862 29886 48914
rect 27246 48850 27298 48862
rect 31502 48850 31554 48862
rect 32286 48914 32338 48926
rect 37550 48914 37602 48926
rect 33170 48862 33182 48914
rect 33234 48862 33246 48914
rect 32286 48850 32338 48862
rect 37550 48850 37602 48862
rect 41134 48914 41186 48926
rect 41134 48850 41186 48862
rect 41694 48914 41746 48926
rect 41694 48850 41746 48862
rect 42702 48914 42754 48926
rect 42702 48850 42754 48862
rect 42814 48914 42866 48926
rect 42814 48850 42866 48862
rect 43486 48914 43538 48926
rect 43486 48850 43538 48862
rect 45502 48914 45554 48926
rect 45502 48850 45554 48862
rect 45614 48914 45666 48926
rect 45614 48850 45666 48862
rect 47406 48914 47458 48926
rect 47406 48850 47458 48862
rect 3054 48802 3106 48814
rect 2146 48750 2158 48802
rect 2210 48750 2222 48802
rect 3054 48738 3106 48750
rect 3614 48802 3666 48814
rect 3614 48738 3666 48750
rect 3838 48802 3890 48814
rect 3838 48738 3890 48750
rect 12238 48802 12290 48814
rect 12238 48738 12290 48750
rect 15150 48802 15202 48814
rect 15150 48738 15202 48750
rect 15486 48802 15538 48814
rect 20190 48802 20242 48814
rect 18610 48750 18622 48802
rect 18674 48750 18686 48802
rect 15486 48738 15538 48750
rect 20190 48738 20242 48750
rect 20750 48802 20802 48814
rect 20750 48738 20802 48750
rect 21646 48802 21698 48814
rect 21646 48738 21698 48750
rect 22094 48802 22146 48814
rect 22094 48738 22146 48750
rect 22542 48802 22594 48814
rect 22542 48738 22594 48750
rect 23214 48802 23266 48814
rect 23214 48738 23266 48750
rect 25454 48802 25506 48814
rect 25454 48738 25506 48750
rect 26350 48802 26402 48814
rect 26350 48738 26402 48750
rect 28814 48802 28866 48814
rect 28814 48738 28866 48750
rect 30942 48802 30994 48814
rect 30942 48738 30994 48750
rect 32398 48802 32450 48814
rect 32398 48738 32450 48750
rect 35086 48802 35138 48814
rect 35086 48738 35138 48750
rect 35534 48802 35586 48814
rect 35534 48738 35586 48750
rect 36878 48802 36930 48814
rect 36878 48738 36930 48750
rect 37886 48802 37938 48814
rect 37886 48738 37938 48750
rect 37998 48802 38050 48814
rect 37998 48738 38050 48750
rect 38670 48802 38722 48814
rect 38670 48738 38722 48750
rect 41582 48802 41634 48814
rect 41582 48738 41634 48750
rect 43038 48802 43090 48814
rect 43038 48738 43090 48750
rect 43710 48802 43762 48814
rect 43710 48738 43762 48750
rect 45838 48802 45890 48814
rect 45838 48738 45890 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 4846 48466 4898 48478
rect 4846 48402 4898 48414
rect 7758 48466 7810 48478
rect 7758 48402 7810 48414
rect 11678 48466 11730 48478
rect 25566 48466 25618 48478
rect 15250 48414 15262 48466
rect 15314 48414 15326 48466
rect 11678 48402 11730 48414
rect 25566 48402 25618 48414
rect 27134 48466 27186 48478
rect 27134 48402 27186 48414
rect 29038 48466 29090 48478
rect 29038 48402 29090 48414
rect 31838 48466 31890 48478
rect 31838 48402 31890 48414
rect 32734 48466 32786 48478
rect 32734 48402 32786 48414
rect 34862 48466 34914 48478
rect 34862 48402 34914 48414
rect 35870 48466 35922 48478
rect 35870 48402 35922 48414
rect 38894 48466 38946 48478
rect 42130 48414 42142 48466
rect 42194 48414 42206 48466
rect 38894 48402 38946 48414
rect 3166 48354 3218 48366
rect 3166 48290 3218 48302
rect 4174 48354 4226 48366
rect 4174 48290 4226 48302
rect 6414 48354 6466 48366
rect 6414 48290 6466 48302
rect 6862 48354 6914 48366
rect 6862 48290 6914 48302
rect 7422 48354 7474 48366
rect 7422 48290 7474 48302
rect 8654 48354 8706 48366
rect 8654 48290 8706 48302
rect 9998 48354 10050 48366
rect 9998 48290 10050 48302
rect 10334 48354 10386 48366
rect 10334 48290 10386 48302
rect 12910 48354 12962 48366
rect 12910 48290 12962 48302
rect 13246 48354 13298 48366
rect 16606 48354 16658 48366
rect 14914 48302 14926 48354
rect 14978 48302 14990 48354
rect 15922 48302 15934 48354
rect 15986 48302 15998 48354
rect 13246 48290 13298 48302
rect 16606 48290 16658 48302
rect 16830 48354 16882 48366
rect 19854 48354 19906 48366
rect 18162 48302 18174 48354
rect 18226 48302 18238 48354
rect 16830 48290 16882 48302
rect 19854 48290 19906 48302
rect 20078 48354 20130 48366
rect 20078 48290 20130 48302
rect 23662 48354 23714 48366
rect 23662 48290 23714 48302
rect 24782 48354 24834 48366
rect 24782 48290 24834 48302
rect 32286 48354 32338 48366
rect 32286 48290 32338 48302
rect 32846 48354 32898 48366
rect 32846 48290 32898 48302
rect 33854 48354 33906 48366
rect 33854 48290 33906 48302
rect 33966 48354 34018 48366
rect 33966 48290 34018 48302
rect 36990 48354 37042 48366
rect 36990 48290 37042 48302
rect 37774 48354 37826 48366
rect 37774 48290 37826 48302
rect 38558 48354 38610 48366
rect 38558 48290 38610 48302
rect 39790 48354 39842 48366
rect 39790 48290 39842 48302
rect 44270 48354 44322 48366
rect 44270 48290 44322 48302
rect 44494 48354 44546 48366
rect 44494 48290 44546 48302
rect 45390 48354 45442 48366
rect 45390 48290 45442 48302
rect 2830 48242 2882 48254
rect 2830 48178 2882 48190
rect 5070 48242 5122 48254
rect 6302 48242 6354 48254
rect 5394 48190 5406 48242
rect 5458 48190 5470 48242
rect 5070 48178 5122 48190
rect 6302 48178 6354 48190
rect 6638 48242 6690 48254
rect 6638 48178 6690 48190
rect 8990 48242 9042 48254
rect 8990 48178 9042 48190
rect 10894 48242 10946 48254
rect 12686 48242 12738 48254
rect 18398 48242 18450 48254
rect 22990 48242 23042 48254
rect 11106 48190 11118 48242
rect 11170 48190 11182 48242
rect 11666 48190 11678 48242
rect 11730 48190 11742 48242
rect 13794 48190 13806 48242
rect 13858 48190 13870 48242
rect 14802 48190 14814 48242
rect 14866 48190 14878 48242
rect 15810 48190 15822 48242
rect 15874 48190 15886 48242
rect 17714 48190 17726 48242
rect 17778 48190 17790 48242
rect 18834 48190 18846 48242
rect 18898 48190 18910 48242
rect 19282 48190 19294 48242
rect 19346 48190 19358 48242
rect 10894 48178 10946 48190
rect 12686 48178 12738 48190
rect 18398 48178 18450 48190
rect 22990 48178 23042 48190
rect 23214 48242 23266 48254
rect 23886 48242 23938 48254
rect 23538 48190 23550 48242
rect 23602 48190 23614 48242
rect 23214 48178 23266 48190
rect 23886 48178 23938 48190
rect 26686 48242 26738 48254
rect 26686 48178 26738 48190
rect 27358 48242 27410 48254
rect 27358 48178 27410 48190
rect 29710 48242 29762 48254
rect 29710 48178 29762 48190
rect 29934 48242 29986 48254
rect 29934 48178 29986 48190
rect 30382 48242 30434 48254
rect 30382 48178 30434 48190
rect 32622 48242 32674 48254
rect 36878 48242 36930 48254
rect 33618 48190 33630 48242
rect 33682 48190 33694 48242
rect 36418 48190 36430 48242
rect 36482 48190 36494 48242
rect 32622 48178 32674 48190
rect 36878 48178 36930 48190
rect 37886 48242 37938 48254
rect 40014 48242 40066 48254
rect 38098 48190 38110 48242
rect 38162 48190 38174 48242
rect 37886 48178 37938 48190
rect 40014 48178 40066 48190
rect 41582 48242 41634 48254
rect 43362 48190 43374 48242
rect 43426 48190 43438 48242
rect 41582 48178 41634 48190
rect 1934 48130 1986 48142
rect 1934 48066 1986 48078
rect 2382 48130 2434 48142
rect 4958 48130 5010 48142
rect 4274 48078 4286 48130
rect 4338 48078 4350 48130
rect 2382 48066 2434 48078
rect 4958 48066 5010 48078
rect 12126 48130 12178 48142
rect 12126 48066 12178 48078
rect 13134 48130 13186 48142
rect 20638 48130 20690 48142
rect 16930 48078 16942 48130
rect 16994 48078 17006 48130
rect 20178 48078 20190 48130
rect 20242 48078 20254 48130
rect 13134 48066 13186 48078
rect 20638 48066 20690 48078
rect 21310 48130 21362 48142
rect 21310 48066 21362 48078
rect 21870 48130 21922 48142
rect 21870 48066 21922 48078
rect 22318 48130 22370 48142
rect 24558 48130 24610 48142
rect 26014 48130 26066 48142
rect 23762 48078 23774 48130
rect 23826 48078 23838 48130
rect 24882 48078 24894 48130
rect 24946 48078 24958 48130
rect 22318 48066 22370 48078
rect 24558 48066 24610 48078
rect 26014 48066 26066 48078
rect 27246 48130 27298 48142
rect 27246 48066 27298 48078
rect 27918 48130 27970 48142
rect 27918 48066 27970 48078
rect 28590 48130 28642 48142
rect 28590 48066 28642 48078
rect 29822 48130 29874 48142
rect 29822 48066 29874 48078
rect 30718 48130 30770 48142
rect 30718 48066 30770 48078
rect 31166 48130 31218 48142
rect 31166 48066 31218 48078
rect 35310 48130 35362 48142
rect 35310 48066 35362 48078
rect 37550 48130 37602 48142
rect 37550 48066 37602 48078
rect 40350 48130 40402 48142
rect 43710 48130 43762 48142
rect 43474 48078 43486 48130
rect 43538 48078 43550 48130
rect 40350 48066 40402 48078
rect 43710 48066 43762 48078
rect 45278 48130 45330 48142
rect 45278 48066 45330 48078
rect 3950 48018 4002 48030
rect 3950 47954 4002 47966
rect 11342 48018 11394 48030
rect 36654 48018 36706 48030
rect 28690 47966 28702 48018
rect 28754 48015 28766 48018
rect 29474 48015 29486 48018
rect 28754 47969 29486 48015
rect 28754 47966 28766 47969
rect 29474 47966 29486 47969
rect 29538 47966 29550 48018
rect 34402 47966 34414 48018
rect 34466 47966 34478 48018
rect 35410 47966 35422 48018
rect 35474 48015 35486 48018
rect 36194 48015 36206 48018
rect 35474 47969 36206 48015
rect 35474 47966 35486 47969
rect 36194 47966 36206 47969
rect 36258 47966 36270 48018
rect 11342 47954 11394 47966
rect 36654 47954 36706 47966
rect 41806 48018 41858 48030
rect 41806 47954 41858 47966
rect 44606 48018 44658 48030
rect 44606 47954 44658 47966
rect 45166 48018 45218 48030
rect 45166 47954 45218 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 14030 47682 14082 47694
rect 5730 47630 5742 47682
rect 5794 47679 5806 47682
rect 6290 47679 6302 47682
rect 5794 47633 6302 47679
rect 5794 47630 5806 47633
rect 6290 47630 6302 47633
rect 6354 47630 6366 47682
rect 14030 47618 14082 47630
rect 14142 47682 14194 47694
rect 14142 47618 14194 47630
rect 14366 47682 14418 47694
rect 20302 47682 20354 47694
rect 17602 47630 17614 47682
rect 17666 47630 17678 47682
rect 14366 47618 14418 47630
rect 20302 47618 20354 47630
rect 20526 47682 20578 47694
rect 20526 47618 20578 47630
rect 22542 47682 22594 47694
rect 22542 47618 22594 47630
rect 24446 47682 24498 47694
rect 37438 47682 37490 47694
rect 30930 47630 30942 47682
rect 30994 47630 31006 47682
rect 24446 47618 24498 47630
rect 37438 47618 37490 47630
rect 4510 47570 4562 47582
rect 3042 47518 3054 47570
rect 3106 47518 3118 47570
rect 4510 47506 4562 47518
rect 5630 47570 5682 47582
rect 5630 47506 5682 47518
rect 6190 47570 6242 47582
rect 6190 47506 6242 47518
rect 8318 47570 8370 47582
rect 8318 47506 8370 47518
rect 9214 47570 9266 47582
rect 9214 47506 9266 47518
rect 9998 47570 10050 47582
rect 9998 47506 10050 47518
rect 12014 47570 12066 47582
rect 18958 47570 19010 47582
rect 25454 47570 25506 47582
rect 31950 47570 32002 47582
rect 12786 47518 12798 47570
rect 12850 47518 12862 47570
rect 16258 47518 16270 47570
rect 16322 47518 16334 47570
rect 23314 47518 23326 47570
rect 23378 47518 23390 47570
rect 27122 47518 27134 47570
rect 27186 47518 27198 47570
rect 28466 47518 28478 47570
rect 28530 47518 28542 47570
rect 30258 47518 30270 47570
rect 30322 47518 30334 47570
rect 12014 47506 12066 47518
rect 18958 47506 19010 47518
rect 25454 47506 25506 47518
rect 31950 47506 32002 47518
rect 37886 47570 37938 47582
rect 37886 47506 37938 47518
rect 39006 47570 39058 47582
rect 39006 47506 39058 47518
rect 45614 47570 45666 47582
rect 45614 47506 45666 47518
rect 2046 47458 2098 47470
rect 8766 47458 8818 47470
rect 3154 47406 3166 47458
rect 3218 47406 3230 47458
rect 2046 47394 2098 47406
rect 8766 47394 8818 47406
rect 9438 47458 9490 47470
rect 14478 47458 14530 47470
rect 11106 47406 11118 47458
rect 11170 47406 11182 47458
rect 9438 47394 9490 47406
rect 14478 47394 14530 47406
rect 15262 47458 15314 47470
rect 17054 47458 17106 47470
rect 19630 47458 19682 47470
rect 16482 47406 16494 47458
rect 16546 47406 16558 47458
rect 17154 47406 17166 47458
rect 17218 47406 17230 47458
rect 17490 47406 17502 47458
rect 17554 47406 17566 47458
rect 15262 47394 15314 47406
rect 17054 47394 17106 47406
rect 19630 47394 19682 47406
rect 19854 47458 19906 47470
rect 21982 47458 22034 47470
rect 19954 47406 19966 47458
rect 20018 47406 20030 47458
rect 19854 47394 19906 47406
rect 21982 47394 22034 47406
rect 22766 47458 22818 47470
rect 23438 47458 23490 47470
rect 23090 47406 23102 47458
rect 23154 47406 23166 47458
rect 22766 47394 22818 47406
rect 23438 47394 23490 47406
rect 24110 47458 24162 47470
rect 28142 47458 28194 47470
rect 32846 47458 32898 47470
rect 24434 47406 24446 47458
rect 24498 47406 24510 47458
rect 26562 47406 26574 47458
rect 26626 47406 26638 47458
rect 27010 47406 27022 47458
rect 27074 47406 27086 47458
rect 30146 47406 30158 47458
rect 30210 47406 30222 47458
rect 24110 47394 24162 47406
rect 28142 47394 28194 47406
rect 32846 47394 32898 47406
rect 33742 47458 33794 47470
rect 33742 47394 33794 47406
rect 33854 47458 33906 47470
rect 33854 47394 33906 47406
rect 34302 47458 34354 47470
rect 35198 47458 35250 47470
rect 34962 47406 34974 47458
rect 35026 47406 35038 47458
rect 34302 47394 34354 47406
rect 35198 47394 35250 47406
rect 35422 47458 35474 47470
rect 35422 47394 35474 47406
rect 35534 47458 35586 47470
rect 35534 47394 35586 47406
rect 38110 47458 38162 47470
rect 38110 47394 38162 47406
rect 38334 47458 38386 47470
rect 38334 47394 38386 47406
rect 41022 47458 41074 47470
rect 43486 47458 43538 47470
rect 41458 47406 41470 47458
rect 41522 47406 41534 47458
rect 43922 47406 43934 47458
rect 43986 47406 43998 47458
rect 46050 47406 46062 47458
rect 46114 47406 46126 47458
rect 41022 47394 41074 47406
rect 43486 47394 43538 47406
rect 8990 47346 9042 47358
rect 6962 47294 6974 47346
rect 7026 47294 7038 47346
rect 8990 47282 9042 47294
rect 10334 47346 10386 47358
rect 10334 47282 10386 47294
rect 10894 47346 10946 47358
rect 10894 47282 10946 47294
rect 12574 47346 12626 47358
rect 28702 47346 28754 47358
rect 21634 47294 21646 47346
rect 21698 47294 21710 47346
rect 26002 47294 26014 47346
rect 26066 47294 26078 47346
rect 27570 47294 27582 47346
rect 27634 47294 27646 47346
rect 12574 47282 12626 47294
rect 28702 47282 28754 47294
rect 33182 47346 33234 47358
rect 33182 47282 33234 47294
rect 34078 47346 34130 47358
rect 34078 47282 34130 47294
rect 38558 47346 38610 47358
rect 38558 47282 38610 47294
rect 39678 47346 39730 47358
rect 39678 47282 39730 47294
rect 41918 47346 41970 47358
rect 41918 47282 41970 47294
rect 43374 47346 43426 47358
rect 43374 47282 43426 47294
rect 2382 47234 2434 47246
rect 2382 47170 2434 47182
rect 3054 47234 3106 47246
rect 3054 47170 3106 47182
rect 5070 47234 5122 47246
rect 5070 47170 5122 47182
rect 6638 47234 6690 47246
rect 6638 47170 6690 47182
rect 7870 47234 7922 47246
rect 7870 47170 7922 47182
rect 12798 47234 12850 47246
rect 12798 47170 12850 47182
rect 14926 47234 14978 47246
rect 14926 47170 14978 47182
rect 15150 47234 15202 47246
rect 15150 47170 15202 47182
rect 19742 47234 19794 47246
rect 19742 47170 19794 47182
rect 23214 47234 23266 47246
rect 23214 47170 23266 47182
rect 25118 47234 25170 47246
rect 25118 47170 25170 47182
rect 28478 47234 28530 47246
rect 28478 47170 28530 47182
rect 31502 47234 31554 47246
rect 31502 47170 31554 47182
rect 36094 47234 36146 47246
rect 45502 47234 45554 47246
rect 36418 47182 36430 47234
rect 36482 47182 36494 47234
rect 36094 47170 36146 47182
rect 45502 47170 45554 47182
rect 45726 47234 45778 47246
rect 45726 47170 45778 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 1934 46898 1986 46910
rect 1934 46834 1986 46846
rect 2830 46898 2882 46910
rect 5406 46898 5458 46910
rect 3154 46846 3166 46898
rect 3218 46846 3230 46898
rect 2830 46834 2882 46846
rect 5406 46834 5458 46846
rect 8094 46898 8146 46910
rect 8094 46834 8146 46846
rect 8878 46898 8930 46910
rect 8878 46834 8930 46846
rect 9662 46898 9714 46910
rect 9662 46834 9714 46846
rect 9774 46898 9826 46910
rect 9774 46834 9826 46846
rect 10670 46898 10722 46910
rect 10670 46834 10722 46846
rect 13918 46898 13970 46910
rect 13918 46834 13970 46846
rect 16382 46898 16434 46910
rect 16382 46834 16434 46846
rect 16494 46898 16546 46910
rect 16494 46834 16546 46846
rect 18510 46898 18562 46910
rect 18510 46834 18562 46846
rect 19070 46898 19122 46910
rect 19070 46834 19122 46846
rect 19854 46898 19906 46910
rect 19854 46834 19906 46846
rect 21086 46898 21138 46910
rect 21086 46834 21138 46846
rect 22542 46898 22594 46910
rect 26126 46898 26178 46910
rect 23090 46846 23102 46898
rect 23154 46846 23166 46898
rect 22542 46834 22594 46846
rect 26126 46834 26178 46846
rect 27582 46898 27634 46910
rect 27582 46834 27634 46846
rect 30718 46898 30770 46910
rect 30718 46834 30770 46846
rect 32510 46898 32562 46910
rect 32510 46834 32562 46846
rect 33630 46898 33682 46910
rect 33630 46834 33682 46846
rect 34414 46898 34466 46910
rect 34414 46834 34466 46846
rect 36542 46898 36594 46910
rect 36542 46834 36594 46846
rect 39230 46898 39282 46910
rect 39230 46834 39282 46846
rect 40462 46898 40514 46910
rect 40462 46834 40514 46846
rect 4286 46786 4338 46798
rect 4286 46722 4338 46734
rect 6526 46786 6578 46798
rect 6526 46722 6578 46734
rect 7982 46786 8034 46798
rect 7982 46722 8034 46734
rect 8766 46786 8818 46798
rect 8766 46722 8818 46734
rect 10222 46786 10274 46798
rect 10222 46722 10274 46734
rect 28030 46786 28082 46798
rect 28030 46722 28082 46734
rect 29934 46786 29986 46798
rect 29934 46722 29986 46734
rect 30270 46786 30322 46798
rect 30270 46722 30322 46734
rect 37662 46786 37714 46798
rect 37662 46722 37714 46734
rect 37998 46786 38050 46798
rect 37998 46722 38050 46734
rect 43710 46786 43762 46798
rect 43710 46722 43762 46734
rect 2270 46674 2322 46686
rect 2270 46610 2322 46622
rect 3838 46674 3890 46686
rect 3838 46610 3890 46622
rect 3950 46674 4002 46686
rect 3950 46610 4002 46622
rect 6414 46674 6466 46686
rect 6414 46610 6466 46622
rect 9102 46674 9154 46686
rect 11230 46674 11282 46686
rect 9986 46622 9998 46674
rect 10050 46622 10062 46674
rect 9102 46610 9154 46622
rect 11230 46610 11282 46622
rect 12126 46674 12178 46686
rect 16606 46674 16658 46686
rect 18398 46674 18450 46686
rect 13458 46622 13470 46674
rect 13522 46622 13534 46674
rect 13682 46622 13694 46674
rect 13746 46622 13758 46674
rect 16930 46622 16942 46674
rect 16994 46622 17006 46674
rect 18050 46622 18062 46674
rect 18114 46622 18126 46674
rect 12126 46610 12178 46622
rect 16606 46610 16658 46622
rect 18398 46610 18450 46622
rect 18622 46674 18674 46686
rect 18622 46610 18674 46622
rect 19630 46674 19682 46686
rect 23438 46674 23490 46686
rect 20066 46622 20078 46674
rect 20130 46622 20142 46674
rect 20402 46622 20414 46674
rect 20466 46622 20478 46674
rect 19630 46610 19682 46622
rect 23438 46610 23490 46622
rect 24334 46674 24386 46686
rect 24334 46610 24386 46622
rect 26910 46674 26962 46686
rect 26910 46610 26962 46622
rect 27134 46674 27186 46686
rect 27134 46610 27186 46622
rect 28142 46674 28194 46686
rect 29486 46674 29538 46686
rect 28578 46622 28590 46674
rect 28642 46622 28654 46674
rect 28142 46610 28194 46622
rect 29486 46610 29538 46622
rect 30046 46674 30098 46686
rect 30046 46610 30098 46622
rect 31278 46674 31330 46686
rect 31278 46610 31330 46622
rect 37214 46674 37266 46686
rect 37214 46610 37266 46622
rect 37438 46674 37490 46686
rect 37438 46610 37490 46622
rect 37886 46674 37938 46686
rect 40350 46674 40402 46686
rect 40002 46622 40014 46674
rect 40066 46622 40078 46674
rect 37886 46610 37938 46622
rect 40350 46610 40402 46622
rect 40574 46674 40626 46686
rect 44606 46674 44658 46686
rect 44146 46622 44158 46674
rect 44210 46622 44222 46674
rect 56130 46622 56142 46674
rect 56194 46622 56206 46674
rect 40574 46610 40626 46622
rect 44606 46610 44658 46622
rect 5070 46562 5122 46574
rect 5070 46498 5122 46510
rect 5854 46562 5906 46574
rect 5854 46498 5906 46510
rect 7534 46562 7586 46574
rect 7534 46498 7586 46510
rect 11566 46562 11618 46574
rect 11566 46498 11618 46510
rect 12462 46562 12514 46574
rect 12462 46498 12514 46510
rect 12910 46562 12962 46574
rect 12910 46498 12962 46510
rect 14478 46562 14530 46574
rect 14478 46498 14530 46510
rect 14926 46562 14978 46574
rect 14926 46498 14978 46510
rect 15374 46562 15426 46574
rect 15374 46498 15426 46510
rect 15822 46562 15874 46574
rect 15822 46498 15874 46510
rect 19742 46562 19794 46574
rect 19742 46498 19794 46510
rect 21422 46562 21474 46574
rect 21422 46498 21474 46510
rect 22206 46562 22258 46574
rect 22206 46498 22258 46510
rect 23886 46562 23938 46574
rect 23886 46498 23938 46510
rect 24782 46562 24834 46574
rect 24782 46498 24834 46510
rect 25678 46562 25730 46574
rect 25678 46498 25730 46510
rect 26686 46562 26738 46574
rect 26686 46498 26738 46510
rect 31726 46562 31778 46574
rect 31726 46498 31778 46510
rect 32062 46562 32114 46574
rect 32062 46498 32114 46510
rect 33966 46562 34018 46574
rect 33966 46498 34018 46510
rect 34862 46562 34914 46574
rect 34862 46498 34914 46510
rect 35310 46562 35362 46574
rect 35310 46498 35362 46510
rect 35758 46562 35810 46574
rect 55346 46510 55358 46562
rect 55410 46510 55422 46562
rect 35758 46498 35810 46510
rect 4174 46450 4226 46462
rect 6526 46450 6578 46462
rect 5170 46398 5182 46450
rect 5234 46447 5246 46450
rect 5730 46447 5742 46450
rect 5234 46401 5742 46447
rect 5234 46398 5246 46401
rect 5730 46398 5742 46401
rect 5794 46398 5806 46450
rect 4174 46386 4226 46398
rect 6526 46386 6578 46398
rect 8094 46450 8146 46462
rect 14030 46450 14082 46462
rect 10434 46398 10446 46450
rect 10498 46447 10510 46450
rect 10994 46447 11006 46450
rect 10498 46401 11006 46447
rect 10498 46398 10510 46401
rect 10994 46398 11006 46401
rect 11058 46398 11070 46450
rect 11442 46398 11454 46450
rect 11506 46447 11518 46450
rect 12898 46447 12910 46450
rect 11506 46401 12910 46447
rect 11506 46398 11518 46401
rect 12898 46398 12910 46401
rect 12962 46398 12974 46450
rect 8094 46386 8146 46398
rect 14030 46386 14082 46398
rect 28366 46450 28418 46462
rect 28366 46386 28418 46398
rect 29710 46450 29762 46462
rect 29710 46386 29762 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 3614 46114 3666 46126
rect 3614 46050 3666 46062
rect 17054 46114 17106 46126
rect 20414 46114 20466 46126
rect 18386 46111 18398 46114
rect 17054 46050 17106 46062
rect 17393 46065 18398 46111
rect 1934 46002 1986 46014
rect 1934 45938 1986 45950
rect 2606 46002 2658 46014
rect 2606 45938 2658 45950
rect 4510 46002 4562 46014
rect 15150 46002 15202 46014
rect 9874 45950 9886 46002
rect 9938 45950 9950 46002
rect 4510 45938 4562 45950
rect 15150 45938 15202 45950
rect 3390 45890 3442 45902
rect 4398 45890 4450 45902
rect 3826 45838 3838 45890
rect 3890 45838 3902 45890
rect 3390 45826 3442 45838
rect 4398 45826 4450 45838
rect 4622 45890 4674 45902
rect 6302 45890 6354 45902
rect 4946 45838 4958 45890
rect 5010 45838 5022 45890
rect 4622 45826 4674 45838
rect 6302 45826 6354 45838
rect 6862 45890 6914 45902
rect 11006 45890 11058 45902
rect 7970 45838 7982 45890
rect 8034 45838 8046 45890
rect 8418 45838 8430 45890
rect 8482 45838 8494 45890
rect 8978 45838 8990 45890
rect 9042 45838 9054 45890
rect 9538 45838 9550 45890
rect 9602 45838 9614 45890
rect 6862 45826 6914 45838
rect 11006 45826 11058 45838
rect 11342 45890 11394 45902
rect 11342 45826 11394 45838
rect 12686 45890 12738 45902
rect 13918 45890 13970 45902
rect 13682 45838 13694 45890
rect 13746 45838 13758 45890
rect 12686 45826 12738 45838
rect 13918 45826 13970 45838
rect 16158 45890 16210 45902
rect 17042 45838 17054 45890
rect 17106 45838 17118 45890
rect 16158 45826 16210 45838
rect 2494 45778 2546 45790
rect 2494 45714 2546 45726
rect 2718 45778 2770 45790
rect 11230 45778 11282 45790
rect 10098 45726 10110 45778
rect 10162 45726 10174 45778
rect 2718 45714 2770 45726
rect 11230 45714 11282 45726
rect 14030 45778 14082 45790
rect 14030 45714 14082 45726
rect 16718 45778 16770 45790
rect 17154 45726 17166 45778
rect 17218 45775 17230 45778
rect 17393 45775 17439 46065
rect 18386 46062 18398 46065
rect 18450 46062 18462 46114
rect 21858 46062 21870 46114
rect 21922 46111 21934 46114
rect 22194 46111 22206 46114
rect 21922 46065 22206 46111
rect 21922 46062 21934 46065
rect 22194 46062 22206 46065
rect 22258 46062 22270 46114
rect 30258 46062 30270 46114
rect 30322 46111 30334 46114
rect 30706 46111 30718 46114
rect 30322 46065 30718 46111
rect 30322 46062 30334 46065
rect 30706 46062 30718 46065
rect 30770 46062 30782 46114
rect 20414 46050 20466 46062
rect 17950 46002 18002 46014
rect 17950 45938 18002 45950
rect 18398 46002 18450 46014
rect 18398 45938 18450 45950
rect 21870 46002 21922 46014
rect 21870 45938 21922 45950
rect 27582 46002 27634 46014
rect 27582 45938 27634 45950
rect 29486 46002 29538 46014
rect 29486 45938 29538 45950
rect 30270 46002 30322 46014
rect 30270 45938 30322 45950
rect 32958 46002 33010 46014
rect 32958 45938 33010 45950
rect 39006 46002 39058 46014
rect 39006 45938 39058 45950
rect 39678 46002 39730 46014
rect 39678 45938 39730 45950
rect 44270 46002 44322 46014
rect 44270 45938 44322 45950
rect 23438 45890 23490 45902
rect 23438 45826 23490 45838
rect 25454 45890 25506 45902
rect 25454 45826 25506 45838
rect 31390 45890 31442 45902
rect 31390 45826 31442 45838
rect 31614 45890 31666 45902
rect 34190 45890 34242 45902
rect 31826 45838 31838 45890
rect 31890 45838 31902 45890
rect 31614 45826 31666 45838
rect 34190 45826 34242 45838
rect 34526 45890 34578 45902
rect 34526 45826 34578 45838
rect 36430 45890 36482 45902
rect 36430 45826 36482 45838
rect 36766 45890 36818 45902
rect 36766 45826 36818 45838
rect 39454 45890 39506 45902
rect 39454 45826 39506 45838
rect 40126 45890 40178 45902
rect 44034 45838 44046 45890
rect 44098 45838 44110 45890
rect 57362 45838 57374 45890
rect 57426 45838 57438 45890
rect 40126 45826 40178 45838
rect 17218 45729 17439 45775
rect 18846 45778 18898 45790
rect 17218 45726 17230 45729
rect 16718 45714 16770 45726
rect 18846 45714 18898 45726
rect 19518 45778 19570 45790
rect 19518 45714 19570 45726
rect 19854 45778 19906 45790
rect 19854 45714 19906 45726
rect 20526 45778 20578 45790
rect 20526 45714 20578 45726
rect 20750 45778 20802 45790
rect 20750 45714 20802 45726
rect 22430 45778 22482 45790
rect 22430 45714 22482 45726
rect 23998 45778 24050 45790
rect 23998 45714 24050 45726
rect 26014 45778 26066 45790
rect 26014 45714 26066 45726
rect 33518 45778 33570 45790
rect 33518 45714 33570 45726
rect 33630 45778 33682 45790
rect 33630 45714 33682 45726
rect 34862 45778 34914 45790
rect 34862 45714 34914 45726
rect 35310 45778 35362 45790
rect 35310 45714 35362 45726
rect 39902 45778 39954 45790
rect 39902 45714 39954 45726
rect 44382 45778 44434 45790
rect 44382 45714 44434 45726
rect 57150 45778 57202 45790
rect 57150 45714 57202 45726
rect 3726 45666 3778 45678
rect 3726 45602 3778 45614
rect 5854 45666 5906 45678
rect 5854 45602 5906 45614
rect 6750 45666 6802 45678
rect 6750 45602 6802 45614
rect 6974 45666 7026 45678
rect 6974 45602 7026 45614
rect 7422 45666 7474 45678
rect 7422 45602 7474 45614
rect 12126 45666 12178 45678
rect 12126 45602 12178 45614
rect 12798 45666 12850 45678
rect 12798 45602 12850 45614
rect 13022 45666 13074 45678
rect 15710 45666 15762 45678
rect 14466 45614 14478 45666
rect 14530 45614 14542 45666
rect 13022 45602 13074 45614
rect 15710 45602 15762 45614
rect 15934 45666 15986 45678
rect 15934 45602 15986 45614
rect 16046 45666 16098 45678
rect 16046 45602 16098 45614
rect 17502 45666 17554 45678
rect 17502 45602 17554 45614
rect 22766 45666 22818 45678
rect 28254 45666 28306 45678
rect 27010 45614 27022 45666
rect 27074 45614 27086 45666
rect 22766 45602 22818 45614
rect 28254 45602 28306 45614
rect 28702 45666 28754 45678
rect 28702 45602 28754 45614
rect 30718 45666 30770 45678
rect 30718 45602 30770 45614
rect 31726 45666 31778 45678
rect 31726 45602 31778 45614
rect 32286 45666 32338 45678
rect 32286 45602 32338 45614
rect 33854 45666 33906 45678
rect 33854 45602 33906 45614
rect 34526 45666 34578 45678
rect 34526 45602 34578 45614
rect 36542 45666 36594 45678
rect 36542 45602 36594 45614
rect 37550 45666 37602 45678
rect 37550 45602 37602 45614
rect 38334 45666 38386 45678
rect 38334 45602 38386 45614
rect 56702 45666 56754 45678
rect 56702 45602 56754 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 5294 45330 5346 45342
rect 5294 45266 5346 45278
rect 13582 45330 13634 45342
rect 13582 45266 13634 45278
rect 13694 45330 13746 45342
rect 13694 45266 13746 45278
rect 14030 45330 14082 45342
rect 14030 45266 14082 45278
rect 14254 45330 14306 45342
rect 21534 45330 21586 45342
rect 20626 45278 20638 45330
rect 20690 45278 20702 45330
rect 14254 45266 14306 45278
rect 21534 45266 21586 45278
rect 23102 45330 23154 45342
rect 23102 45266 23154 45278
rect 23662 45330 23714 45342
rect 23662 45266 23714 45278
rect 28926 45330 28978 45342
rect 28926 45266 28978 45278
rect 38110 45330 38162 45342
rect 38110 45266 38162 45278
rect 38894 45330 38946 45342
rect 38894 45266 38946 45278
rect 40126 45330 40178 45342
rect 40126 45266 40178 45278
rect 4286 45218 4338 45230
rect 4286 45154 4338 45166
rect 6974 45218 7026 45230
rect 6974 45154 7026 45166
rect 8206 45218 8258 45230
rect 8206 45154 8258 45166
rect 8878 45218 8930 45230
rect 11454 45218 11506 45230
rect 9762 45166 9774 45218
rect 9826 45166 9838 45218
rect 8878 45154 8930 45166
rect 11454 45154 11506 45166
rect 15150 45218 15202 45230
rect 15150 45154 15202 45166
rect 18846 45218 18898 45230
rect 18846 45154 18898 45166
rect 18958 45218 19010 45230
rect 21870 45218 21922 45230
rect 19730 45166 19742 45218
rect 19794 45166 19806 45218
rect 18958 45154 19010 45166
rect 21870 45154 21922 45166
rect 22766 45218 22818 45230
rect 22766 45154 22818 45166
rect 27358 45218 27410 45230
rect 27358 45154 27410 45166
rect 28030 45218 28082 45230
rect 28030 45154 28082 45166
rect 31054 45218 31106 45230
rect 31054 45154 31106 45166
rect 34302 45218 34354 45230
rect 34302 45154 34354 45166
rect 37214 45218 37266 45230
rect 37214 45154 37266 45166
rect 40014 45218 40066 45230
rect 40014 45154 40066 45166
rect 43038 45218 43090 45230
rect 43038 45154 43090 45166
rect 44494 45218 44546 45230
rect 44494 45154 44546 45166
rect 5630 45106 5682 45118
rect 2818 45054 2830 45106
rect 2882 45054 2894 45106
rect 3938 45054 3950 45106
rect 4002 45054 4014 45106
rect 5630 45042 5682 45054
rect 6862 45106 6914 45118
rect 6862 45042 6914 45054
rect 7086 45106 7138 45118
rect 8430 45106 8482 45118
rect 7522 45054 7534 45106
rect 7586 45054 7598 45106
rect 7086 45042 7138 45054
rect 8430 45042 8482 45054
rect 8654 45106 8706 45118
rect 11678 45106 11730 45118
rect 10098 45054 10110 45106
rect 10162 45054 10174 45106
rect 10882 45054 10894 45106
rect 10946 45054 10958 45106
rect 8654 45042 8706 45054
rect 11678 45042 11730 45054
rect 12014 45106 12066 45118
rect 12014 45042 12066 45054
rect 13022 45106 13074 45118
rect 14366 45106 14418 45118
rect 13346 45054 13358 45106
rect 13410 45054 13422 45106
rect 13022 45042 13074 45054
rect 14366 45042 14418 45054
rect 16942 45106 16994 45118
rect 21758 45106 21810 45118
rect 19618 45054 19630 45106
rect 19682 45054 19694 45106
rect 20738 45054 20750 45106
rect 20802 45054 20814 45106
rect 21298 45054 21310 45106
rect 21362 45054 21374 45106
rect 16942 45042 16994 45054
rect 21758 45042 21810 45054
rect 24446 45106 24498 45118
rect 24446 45042 24498 45054
rect 25790 45106 25842 45118
rect 25790 45042 25842 45054
rect 25902 45106 25954 45118
rect 25902 45042 25954 45054
rect 26126 45106 26178 45118
rect 26126 45042 26178 45054
rect 26238 45106 26290 45118
rect 26238 45042 26290 45054
rect 26686 45106 26738 45118
rect 26686 45042 26738 45054
rect 27134 45106 27186 45118
rect 27134 45042 27186 45054
rect 27918 45106 27970 45118
rect 27918 45042 27970 45054
rect 28142 45106 28194 45118
rect 28142 45042 28194 45054
rect 28590 45106 28642 45118
rect 28590 45042 28642 45054
rect 29598 45106 29650 45118
rect 32622 45106 32674 45118
rect 29922 45054 29934 45106
rect 29986 45054 29998 45106
rect 29598 45042 29650 45054
rect 32622 45042 32674 45054
rect 33630 45106 33682 45118
rect 33630 45042 33682 45054
rect 34414 45106 34466 45118
rect 34414 45042 34466 45054
rect 34526 45106 34578 45118
rect 35758 45106 35810 45118
rect 34962 45054 34974 45106
rect 35026 45054 35038 45106
rect 35522 45054 35534 45106
rect 35586 45054 35598 45106
rect 34526 45042 34578 45054
rect 35758 45042 35810 45054
rect 36654 45106 36706 45118
rect 42702 45106 42754 45118
rect 36978 45054 36990 45106
rect 37042 45054 37054 45106
rect 39554 45054 39566 45106
rect 39618 45054 39630 45106
rect 39778 45054 39790 45106
rect 39842 45054 39854 45106
rect 36654 45042 36706 45054
rect 42702 45042 42754 45054
rect 43934 45106 43986 45118
rect 43934 45042 43986 45054
rect 44158 45106 44210 45118
rect 44158 45042 44210 45054
rect 4174 44994 4226 45006
rect 1922 44942 1934 44994
rect 1986 44942 1998 44994
rect 4174 44930 4226 44942
rect 4846 44994 4898 45006
rect 4846 44930 4898 44942
rect 6302 44994 6354 45006
rect 6302 44930 6354 44942
rect 8990 44994 9042 45006
rect 11902 44994 11954 45006
rect 10322 44942 10334 44994
rect 10386 44942 10398 44994
rect 8990 44930 9042 44942
rect 11902 44930 11954 44942
rect 12574 44994 12626 45006
rect 12574 44930 12626 44942
rect 15598 44994 15650 45006
rect 15598 44930 15650 44942
rect 16046 44994 16098 45006
rect 16046 44930 16098 44942
rect 16494 44994 16546 45006
rect 16494 44930 16546 44942
rect 17950 44994 18002 45006
rect 17950 44930 18002 44942
rect 21646 44994 21698 45006
rect 21646 44930 21698 44942
rect 24222 44994 24274 45006
rect 24222 44930 24274 44942
rect 26910 44994 26962 45006
rect 26910 44930 26962 44942
rect 30494 44994 30546 45006
rect 37662 44994 37714 45006
rect 40462 44994 40514 45006
rect 31378 44942 31390 44994
rect 31442 44942 31454 44994
rect 38994 44942 39006 44994
rect 39058 44942 39070 44994
rect 30494 44930 30546 44942
rect 37662 44930 37714 44942
rect 40462 44930 40514 44942
rect 44382 44994 44434 45006
rect 44382 44930 44434 44942
rect 18958 44882 19010 44894
rect 32734 44882 32786 44894
rect 6066 44830 6078 44882
rect 6130 44879 6142 44882
rect 6290 44879 6302 44882
rect 6130 44833 6302 44879
rect 6130 44830 6142 44833
rect 6290 44830 6302 44833
rect 6354 44830 6366 44882
rect 15250 44830 15262 44882
rect 15314 44879 15326 44882
rect 15922 44879 15934 44882
rect 15314 44833 15934 44879
rect 15314 44830 15326 44833
rect 15922 44830 15934 44833
rect 15986 44879 15998 44882
rect 16482 44879 16494 44882
rect 15986 44833 16494 44879
rect 15986 44830 15998 44833
rect 16482 44830 16494 44833
rect 16546 44879 16558 44882
rect 17154 44879 17166 44882
rect 16546 44833 17166 44879
rect 16546 44830 16558 44833
rect 17154 44830 17166 44833
rect 17218 44830 17230 44882
rect 24770 44830 24782 44882
rect 24834 44830 24846 44882
rect 31266 44830 31278 44882
rect 31330 44830 31342 44882
rect 18958 44818 19010 44830
rect 32734 44818 32786 44830
rect 35982 44882 36034 44894
rect 35982 44818 36034 44830
rect 36094 44882 36146 44894
rect 36094 44818 36146 44830
rect 37326 44882 37378 44894
rect 37326 44818 37378 44830
rect 38670 44882 38722 44894
rect 38670 44818 38722 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 6302 44546 6354 44558
rect 12462 44546 12514 44558
rect 10770 44494 10782 44546
rect 10834 44543 10846 44546
rect 11554 44543 11566 44546
rect 10834 44497 11566 44543
rect 10834 44494 10846 44497
rect 11554 44494 11566 44497
rect 11618 44494 11630 44546
rect 6302 44482 6354 44494
rect 12462 44482 12514 44494
rect 12910 44546 12962 44558
rect 12910 44482 12962 44494
rect 15262 44546 15314 44558
rect 15262 44482 15314 44494
rect 17390 44546 17442 44558
rect 17390 44482 17442 44494
rect 20190 44546 20242 44558
rect 32958 44546 33010 44558
rect 25778 44494 25790 44546
rect 25842 44543 25854 44546
rect 26338 44543 26350 44546
rect 25842 44497 26350 44543
rect 25842 44494 25854 44497
rect 26338 44494 26350 44497
rect 26402 44494 26414 44546
rect 30706 44494 30718 44546
rect 30770 44543 30782 44546
rect 31378 44543 31390 44546
rect 30770 44497 31390 44543
rect 30770 44494 30782 44497
rect 31378 44494 31390 44497
rect 31442 44494 31454 44546
rect 20190 44482 20242 44494
rect 32958 44482 33010 44494
rect 38110 44546 38162 44558
rect 38110 44482 38162 44494
rect 38334 44546 38386 44558
rect 38334 44482 38386 44494
rect 39006 44546 39058 44558
rect 39006 44482 39058 44494
rect 45502 44546 45554 44558
rect 45502 44482 45554 44494
rect 2046 44434 2098 44446
rect 2046 44370 2098 44382
rect 2494 44434 2546 44446
rect 10782 44434 10834 44446
rect 6850 44382 6862 44434
rect 6914 44382 6926 44434
rect 2494 44370 2546 44382
rect 10782 44370 10834 44382
rect 18286 44434 18338 44446
rect 18286 44370 18338 44382
rect 18846 44434 18898 44446
rect 18846 44370 18898 44382
rect 25342 44434 25394 44446
rect 25342 44370 25394 44382
rect 25902 44434 25954 44446
rect 25902 44370 25954 44382
rect 26350 44434 26402 44446
rect 26350 44370 26402 44382
rect 27134 44434 27186 44446
rect 27134 44370 27186 44382
rect 31166 44434 31218 44446
rect 31166 44370 31218 44382
rect 35646 44434 35698 44446
rect 42366 44434 42418 44446
rect 40114 44382 40126 44434
rect 40178 44382 40190 44434
rect 35646 44370 35698 44382
rect 42366 44370 42418 44382
rect 43486 44434 43538 44446
rect 43486 44370 43538 44382
rect 2942 44322 2994 44334
rect 7534 44322 7586 44334
rect 9662 44322 9714 44334
rect 12014 44322 12066 44334
rect 6962 44270 6974 44322
rect 7026 44270 7038 44322
rect 8418 44270 8430 44322
rect 8482 44270 8494 44322
rect 9202 44270 9214 44322
rect 9266 44270 9278 44322
rect 9762 44270 9774 44322
rect 9826 44270 9838 44322
rect 2942 44258 2994 44270
rect 7534 44258 7586 44270
rect 9662 44258 9714 44270
rect 12014 44258 12066 44270
rect 12238 44322 12290 44334
rect 12238 44258 12290 44270
rect 15374 44322 15426 44334
rect 15374 44258 15426 44270
rect 15598 44322 15650 44334
rect 15598 44258 15650 44270
rect 18734 44322 18786 44334
rect 21870 44322 21922 44334
rect 19282 44270 19294 44322
rect 19346 44270 19358 44322
rect 18734 44258 18786 44270
rect 21870 44258 21922 44270
rect 23214 44322 23266 44334
rect 23214 44258 23266 44270
rect 23326 44322 23378 44334
rect 23326 44258 23378 44270
rect 24110 44322 24162 44334
rect 29934 44322 29986 44334
rect 32622 44322 32674 44334
rect 28018 44270 28030 44322
rect 28082 44270 28094 44322
rect 28578 44270 28590 44322
rect 28642 44270 28654 44322
rect 31938 44270 31950 44322
rect 32002 44270 32014 44322
rect 24110 44258 24162 44270
rect 29934 44258 29986 44270
rect 32622 44258 32674 44270
rect 36206 44322 36258 44334
rect 36206 44258 36258 44270
rect 36766 44322 36818 44334
rect 36766 44258 36818 44270
rect 38558 44322 38610 44334
rect 41806 44322 41858 44334
rect 39666 44270 39678 44322
rect 39730 44270 39742 44322
rect 41010 44270 41022 44322
rect 41074 44270 41086 44322
rect 38558 44258 38610 44270
rect 41806 44258 41858 44270
rect 42814 44322 42866 44334
rect 44046 44322 44098 44334
rect 43138 44270 43150 44322
rect 43202 44270 43214 44322
rect 42814 44258 42866 44270
rect 44046 44258 44098 44270
rect 44158 44322 44210 44334
rect 44158 44258 44210 44270
rect 44270 44322 44322 44334
rect 44706 44270 44718 44322
rect 44770 44270 44782 44322
rect 45490 44270 45502 44322
rect 45554 44270 45566 44322
rect 44270 44258 44322 44270
rect 5742 44210 5794 44222
rect 4162 44158 4174 44210
rect 4226 44158 4238 44210
rect 5742 44146 5794 44158
rect 6190 44210 6242 44222
rect 9438 44210 9490 44222
rect 8082 44158 8094 44210
rect 8146 44158 8158 44210
rect 6190 44146 6242 44158
rect 9438 44146 9490 44158
rect 11790 44210 11842 44222
rect 11790 44146 11842 44158
rect 13694 44210 13746 44222
rect 13694 44146 13746 44158
rect 15710 44210 15762 44222
rect 15710 44146 15762 44158
rect 16606 44210 16658 44222
rect 16606 44146 16658 44158
rect 16718 44210 16770 44222
rect 16718 44146 16770 44158
rect 17502 44210 17554 44222
rect 17502 44146 17554 44158
rect 19854 44210 19906 44222
rect 19854 44146 19906 44158
rect 20078 44210 20130 44222
rect 20078 44146 20130 44158
rect 21982 44210 22034 44222
rect 21982 44146 22034 44158
rect 22094 44210 22146 44222
rect 22094 44146 22146 44158
rect 23102 44210 23154 44222
rect 23102 44146 23154 44158
rect 23662 44210 23714 44222
rect 23662 44146 23714 44158
rect 26686 44210 26738 44222
rect 29598 44210 29650 44222
rect 35534 44210 35586 44222
rect 27682 44158 27694 44210
rect 27746 44158 27758 44210
rect 32050 44158 32062 44210
rect 32114 44158 32126 44210
rect 26686 44146 26738 44158
rect 29598 44146 29650 44158
rect 35534 44146 35586 44158
rect 35758 44210 35810 44222
rect 35758 44146 35810 44158
rect 37886 44210 37938 44222
rect 37886 44146 37938 44158
rect 45838 44210 45890 44222
rect 45838 44146 45890 44158
rect 3278 44098 3330 44110
rect 3278 44034 3330 44046
rect 3838 44098 3890 44110
rect 3838 44034 3890 44046
rect 5070 44098 5122 44110
rect 5070 44034 5122 44046
rect 5966 44098 6018 44110
rect 5966 44034 6018 44046
rect 11342 44098 11394 44110
rect 11342 44034 11394 44046
rect 14142 44098 14194 44110
rect 14142 44034 14194 44046
rect 14590 44098 14642 44110
rect 14590 44034 14642 44046
rect 16382 44098 16434 44110
rect 16382 44034 16434 44046
rect 17390 44098 17442 44110
rect 17390 44034 17442 44046
rect 18958 44098 19010 44110
rect 18958 44034 19010 44046
rect 20638 44098 20690 44110
rect 24558 44098 24610 44110
rect 29710 44098 29762 44110
rect 22530 44046 22542 44098
rect 22594 44046 22606 44098
rect 28578 44046 28590 44098
rect 28642 44046 28654 44098
rect 20638 44034 20690 44046
rect 24558 44034 24610 44046
rect 29710 44034 29762 44046
rect 30270 44098 30322 44110
rect 30270 44034 30322 44046
rect 30718 44098 30770 44110
rect 30718 44034 30770 44046
rect 33518 44098 33570 44110
rect 33518 44034 33570 44046
rect 43374 44098 43426 44110
rect 43374 44034 43426 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 7870 43762 7922 43774
rect 4498 43710 4510 43762
rect 4562 43710 4574 43762
rect 7870 43698 7922 43710
rect 9774 43762 9826 43774
rect 12574 43762 12626 43774
rect 10770 43710 10782 43762
rect 10834 43710 10846 43762
rect 9774 43698 9826 43710
rect 12574 43698 12626 43710
rect 27582 43762 27634 43774
rect 27582 43698 27634 43710
rect 28030 43762 28082 43774
rect 28030 43698 28082 43710
rect 28254 43762 28306 43774
rect 28254 43698 28306 43710
rect 29710 43762 29762 43774
rect 29710 43698 29762 43710
rect 37214 43762 37266 43774
rect 37214 43698 37266 43710
rect 37998 43762 38050 43774
rect 37998 43698 38050 43710
rect 43934 43762 43986 43774
rect 43934 43698 43986 43710
rect 46062 43762 46114 43774
rect 46062 43698 46114 43710
rect 2830 43650 2882 43662
rect 2830 43586 2882 43598
rect 3614 43650 3666 43662
rect 3614 43586 3666 43598
rect 7646 43650 7698 43662
rect 7646 43586 7698 43598
rect 7982 43650 8034 43662
rect 7982 43586 8034 43598
rect 8542 43650 8594 43662
rect 8542 43586 8594 43598
rect 13582 43650 13634 43662
rect 13582 43586 13634 43598
rect 13694 43650 13746 43662
rect 13694 43586 13746 43598
rect 15150 43650 15202 43662
rect 15150 43586 15202 43598
rect 16718 43650 16770 43662
rect 16718 43586 16770 43598
rect 18846 43650 18898 43662
rect 18846 43586 18898 43598
rect 19966 43650 20018 43662
rect 19966 43586 20018 43598
rect 20190 43650 20242 43662
rect 20190 43586 20242 43598
rect 20638 43650 20690 43662
rect 20638 43586 20690 43598
rect 22094 43650 22146 43662
rect 24222 43650 24274 43662
rect 23426 43598 23438 43650
rect 23490 43598 23502 43650
rect 22094 43586 22146 43598
rect 24222 43586 24274 43598
rect 26350 43650 26402 43662
rect 26350 43586 26402 43598
rect 27246 43650 27298 43662
rect 27246 43586 27298 43598
rect 27358 43650 27410 43662
rect 27358 43586 27410 43598
rect 28142 43650 28194 43662
rect 28142 43586 28194 43598
rect 29374 43650 29426 43662
rect 29374 43586 29426 43598
rect 39454 43650 39506 43662
rect 39454 43586 39506 43598
rect 39902 43650 39954 43662
rect 39902 43586 39954 43598
rect 40798 43650 40850 43662
rect 40798 43586 40850 43598
rect 42590 43650 42642 43662
rect 42590 43586 42642 43598
rect 43710 43650 43762 43662
rect 43710 43586 43762 43598
rect 44046 43650 44098 43662
rect 44046 43586 44098 43598
rect 46174 43650 46226 43662
rect 46174 43586 46226 43598
rect 3278 43538 3330 43550
rect 3278 43474 3330 43486
rect 4174 43538 4226 43550
rect 4174 43474 4226 43486
rect 7422 43538 7474 43550
rect 7422 43474 7474 43486
rect 11118 43538 11170 43550
rect 11118 43474 11170 43486
rect 11902 43538 11954 43550
rect 11902 43474 11954 43486
rect 12350 43538 12402 43550
rect 12350 43474 12402 43486
rect 12462 43538 12514 43550
rect 12462 43474 12514 43486
rect 13358 43538 13410 43550
rect 14590 43538 14642 43550
rect 14018 43486 14030 43538
rect 14082 43486 14094 43538
rect 13358 43474 13410 43486
rect 14590 43474 14642 43486
rect 15038 43538 15090 43550
rect 15038 43474 15090 43486
rect 15262 43538 15314 43550
rect 15262 43474 15314 43486
rect 16382 43538 16434 43550
rect 16382 43474 16434 43486
rect 16494 43538 16546 43550
rect 16494 43474 16546 43486
rect 16942 43538 16994 43550
rect 16942 43474 16994 43486
rect 17726 43538 17778 43550
rect 21534 43538 21586 43550
rect 19394 43486 19406 43538
rect 19458 43486 19470 43538
rect 19730 43486 19742 43538
rect 19794 43486 19806 43538
rect 17726 43474 17778 43486
rect 21534 43474 21586 43486
rect 22542 43538 22594 43550
rect 28702 43538 28754 43550
rect 34526 43538 34578 43550
rect 22978 43486 22990 43538
rect 23042 43486 23054 43538
rect 23986 43486 23998 43538
rect 24050 43486 24062 43538
rect 34290 43486 34302 43538
rect 34354 43486 34366 43538
rect 22542 43474 22594 43486
rect 28702 43474 28754 43486
rect 34526 43474 34578 43486
rect 34638 43538 34690 43550
rect 37662 43538 37714 43550
rect 35074 43486 35086 43538
rect 35138 43486 35150 43538
rect 35634 43486 35646 43538
rect 35698 43486 35710 43538
rect 34638 43474 34690 43486
rect 37662 43474 37714 43486
rect 38670 43538 38722 43550
rect 38670 43474 38722 43486
rect 39230 43538 39282 43550
rect 39230 43474 39282 43486
rect 41806 43538 41858 43550
rect 42702 43538 42754 43550
rect 42354 43486 42366 43538
rect 42418 43486 42430 43538
rect 41806 43474 41858 43486
rect 42702 43474 42754 43486
rect 44158 43538 44210 43550
rect 44158 43474 44210 43486
rect 44830 43538 44882 43550
rect 44830 43474 44882 43486
rect 45054 43538 45106 43550
rect 45054 43474 45106 43486
rect 45950 43538 46002 43550
rect 45950 43474 46002 43486
rect 1934 43426 1986 43438
rect 1934 43362 1986 43374
rect 2382 43426 2434 43438
rect 2382 43362 2434 43374
rect 5182 43426 5234 43438
rect 5182 43362 5234 43374
rect 5518 43426 5570 43438
rect 5518 43362 5570 43374
rect 6078 43426 6130 43438
rect 6078 43362 6130 43374
rect 6526 43426 6578 43438
rect 6526 43362 6578 43374
rect 6974 43426 7026 43438
rect 6974 43362 7026 43374
rect 8990 43426 9042 43438
rect 8990 43362 9042 43374
rect 10222 43426 10274 43438
rect 10222 43362 10274 43374
rect 12126 43426 12178 43438
rect 15822 43426 15874 43438
rect 14130 43374 14142 43426
rect 14194 43374 14206 43426
rect 12126 43362 12178 43374
rect 15822 43362 15874 43374
rect 17054 43426 17106 43438
rect 17054 43362 17106 43374
rect 18062 43426 18114 43438
rect 18062 43362 18114 43374
rect 20078 43426 20130 43438
rect 20078 43362 20130 43374
rect 21086 43426 21138 43438
rect 21086 43362 21138 43374
rect 25006 43426 25058 43438
rect 25006 43362 25058 43374
rect 25902 43426 25954 43438
rect 25902 43362 25954 43374
rect 30158 43426 30210 43438
rect 30158 43362 30210 43374
rect 30606 43426 30658 43438
rect 30606 43362 30658 43374
rect 31166 43426 31218 43438
rect 31166 43362 31218 43374
rect 31502 43426 31554 43438
rect 31502 43362 31554 43374
rect 32062 43426 32114 43438
rect 32062 43362 32114 43374
rect 32286 43426 32338 43438
rect 32286 43362 32338 43374
rect 32622 43426 32674 43438
rect 32622 43362 32674 43374
rect 33518 43426 33570 43438
rect 33518 43362 33570 43374
rect 36654 43426 36706 43438
rect 36654 43362 36706 43374
rect 40350 43426 40402 43438
rect 40350 43362 40402 43374
rect 26014 43314 26066 43326
rect 5170 43262 5182 43314
rect 5234 43311 5246 43314
rect 6626 43311 6638 43314
rect 5234 43265 6638 43311
rect 5234 43262 5246 43265
rect 6626 43262 6638 43265
rect 6690 43262 6702 43314
rect 26014 43250 26066 43262
rect 26238 43314 26290 43326
rect 26238 43250 26290 43262
rect 35870 43314 35922 43326
rect 35870 43250 35922 43262
rect 36094 43314 36146 43326
rect 36094 43250 36146 43262
rect 36206 43314 36258 43326
rect 36206 43250 36258 43262
rect 38894 43314 38946 43326
rect 38894 43250 38946 43262
rect 39342 43314 39394 43326
rect 45390 43314 45442 43326
rect 39666 43262 39678 43314
rect 39730 43311 39742 43314
rect 40338 43311 40350 43314
rect 39730 43265 40350 43311
rect 39730 43262 39742 43265
rect 40338 43262 40350 43265
rect 40402 43262 40414 43314
rect 43138 43262 43150 43314
rect 43202 43262 43214 43314
rect 39342 43250 39394 43262
rect 45390 43250 45442 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 4510 42978 4562 42990
rect 16382 42978 16434 42990
rect 18062 42978 18114 42990
rect 12674 42926 12686 42978
rect 12738 42926 12750 42978
rect 14242 42926 14254 42978
rect 14306 42926 14318 42978
rect 17042 42926 17054 42978
rect 17106 42975 17118 42978
rect 17106 42929 17663 42975
rect 17106 42926 17118 42929
rect 4510 42914 4562 42926
rect 16382 42914 16434 42926
rect 2606 42866 2658 42878
rect 5630 42866 5682 42878
rect 3826 42814 3838 42866
rect 3890 42814 3902 42866
rect 2606 42802 2658 42814
rect 5630 42802 5682 42814
rect 8990 42866 9042 42878
rect 16942 42866 16994 42878
rect 9874 42814 9886 42866
rect 9938 42814 9950 42866
rect 8990 42802 9042 42814
rect 16942 42802 16994 42814
rect 2382 42754 2434 42766
rect 2382 42690 2434 42702
rect 2718 42754 2770 42766
rect 6414 42754 6466 42766
rect 3602 42702 3614 42754
rect 3666 42702 3678 42754
rect 4610 42702 4622 42754
rect 4674 42702 4686 42754
rect 2718 42690 2770 42702
rect 6414 42690 6466 42702
rect 6750 42754 6802 42766
rect 12014 42754 12066 42766
rect 7522 42702 7534 42754
rect 7586 42702 7598 42754
rect 10658 42702 10670 42754
rect 10722 42702 10734 42754
rect 11330 42702 11342 42754
rect 11394 42702 11406 42754
rect 12114 42702 12126 42754
rect 12178 42702 12190 42754
rect 14242 42702 14254 42754
rect 14306 42702 14318 42754
rect 6750 42690 6802 42702
rect 12014 42690 12066 42702
rect 2158 42642 2210 42654
rect 2158 42578 2210 42590
rect 6526 42642 6578 42654
rect 6526 42578 6578 42590
rect 6638 42642 6690 42654
rect 6638 42578 6690 42590
rect 7758 42642 7810 42654
rect 7758 42578 7810 42590
rect 9550 42642 9602 42654
rect 13694 42642 13746 42654
rect 15822 42642 15874 42654
rect 10434 42590 10446 42642
rect 10498 42590 10510 42642
rect 13906 42590 13918 42642
rect 13970 42590 13982 42642
rect 17617 42639 17663 42929
rect 18062 42914 18114 42926
rect 18286 42978 18338 42990
rect 18286 42914 18338 42926
rect 18398 42978 18450 42990
rect 18398 42914 18450 42926
rect 18958 42978 19010 42990
rect 18958 42914 19010 42926
rect 26238 42978 26290 42990
rect 26238 42914 26290 42926
rect 26686 42978 26738 42990
rect 39902 42978 39954 42990
rect 27346 42926 27358 42978
rect 27410 42975 27422 42978
rect 28018 42975 28030 42978
rect 27410 42929 28030 42975
rect 27410 42926 27422 42929
rect 28018 42926 28030 42929
rect 28082 42926 28094 42978
rect 26686 42914 26738 42926
rect 39902 42914 39954 42926
rect 40350 42978 40402 42990
rect 40350 42914 40402 42926
rect 43934 42978 43986 42990
rect 43934 42914 43986 42926
rect 44158 42978 44210 42990
rect 44158 42914 44210 42926
rect 19406 42866 19458 42878
rect 20862 42866 20914 42878
rect 26014 42866 26066 42878
rect 19730 42814 19742 42866
rect 19794 42814 19806 42866
rect 22978 42814 22990 42866
rect 23042 42814 23054 42866
rect 19406 42802 19458 42814
rect 20862 42802 20914 42814
rect 26014 42802 26066 42814
rect 29486 42866 29538 42878
rect 29486 42802 29538 42814
rect 29934 42866 29986 42878
rect 29934 42802 29986 42814
rect 31726 42866 31778 42878
rect 31726 42802 31778 42814
rect 34862 42866 34914 42878
rect 34862 42802 34914 42814
rect 41022 42866 41074 42878
rect 41022 42802 41074 42814
rect 43262 42866 43314 42878
rect 43262 42802 43314 42814
rect 17950 42754 18002 42766
rect 17950 42690 18002 42702
rect 19182 42754 19234 42766
rect 19182 42690 19234 42702
rect 19854 42754 19906 42766
rect 19854 42690 19906 42702
rect 25790 42754 25842 42766
rect 31838 42754 31890 42766
rect 31490 42702 31502 42754
rect 31554 42702 31566 42754
rect 25790 42690 25842 42702
rect 31838 42690 31890 42702
rect 32062 42754 32114 42766
rect 32062 42690 32114 42702
rect 34638 42754 34690 42766
rect 40126 42754 40178 42766
rect 44270 42754 44322 42766
rect 39666 42702 39678 42754
rect 39730 42702 39742 42754
rect 43698 42702 43710 42754
rect 43762 42702 43774 42754
rect 34638 42690 34690 42702
rect 40126 42690 40178 42702
rect 44270 42690 44322 42702
rect 22430 42642 22482 42654
rect 17826 42639 17838 42642
rect 17617 42593 17838 42639
rect 17826 42590 17838 42593
rect 17890 42590 17902 42642
rect 9550 42578 9602 42590
rect 13694 42578 13746 42590
rect 15822 42578 15874 42590
rect 22430 42578 22482 42590
rect 22542 42642 22594 42654
rect 23662 42642 23714 42654
rect 22642 42590 22654 42642
rect 22706 42590 22718 42642
rect 22542 42578 22594 42590
rect 23662 42578 23714 42590
rect 23998 42642 24050 42654
rect 23998 42578 24050 42590
rect 28254 42642 28306 42654
rect 28254 42578 28306 42590
rect 28366 42642 28418 42654
rect 28366 42578 28418 42590
rect 30494 42642 30546 42654
rect 30494 42578 30546 42590
rect 30718 42642 30770 42654
rect 34414 42642 34466 42654
rect 33058 42590 33070 42642
rect 33122 42590 33134 42642
rect 30718 42578 30770 42590
rect 34414 42578 34466 42590
rect 34974 42642 35026 42654
rect 34974 42578 35026 42590
rect 35534 42642 35586 42654
rect 35534 42578 35586 42590
rect 35758 42642 35810 42654
rect 35758 42578 35810 42590
rect 35982 42642 36034 42654
rect 35982 42578 36034 42590
rect 37774 42642 37826 42654
rect 37774 42578 37826 42590
rect 38110 42642 38162 42654
rect 38110 42578 38162 42590
rect 6302 42530 6354 42542
rect 6302 42466 6354 42478
rect 8542 42530 8594 42542
rect 8542 42466 8594 42478
rect 9774 42530 9826 42542
rect 9774 42466 9826 42478
rect 14478 42530 14530 42542
rect 14478 42466 14530 42478
rect 15374 42530 15426 42542
rect 15374 42466 15426 42478
rect 16046 42530 16098 42542
rect 16046 42466 16098 42478
rect 16270 42530 16322 42542
rect 16270 42466 16322 42478
rect 17390 42530 17442 42542
rect 17390 42466 17442 42478
rect 19630 42530 19682 42542
rect 19630 42466 19682 42478
rect 20526 42530 20578 42542
rect 20526 42466 20578 42478
rect 21646 42530 21698 42542
rect 21646 42466 21698 42478
rect 22206 42530 22258 42542
rect 22206 42466 22258 42478
rect 24446 42530 24498 42542
rect 24446 42466 24498 42478
rect 25230 42530 25282 42542
rect 25230 42466 25282 42478
rect 27358 42530 27410 42542
rect 27358 42466 27410 42478
rect 27694 42530 27746 42542
rect 27694 42466 27746 42478
rect 28590 42530 28642 42542
rect 28590 42466 28642 42478
rect 30606 42530 30658 42542
rect 30606 42466 30658 42478
rect 35422 42530 35474 42542
rect 35422 42466 35474 42478
rect 38558 42530 38610 42542
rect 38558 42466 38610 42478
rect 39006 42530 39058 42542
rect 39006 42466 39058 42478
rect 40238 42530 40290 42542
rect 40238 42466 40290 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 2830 42194 2882 42206
rect 2830 42130 2882 42142
rect 3838 42194 3890 42206
rect 3838 42130 3890 42142
rect 7310 42194 7362 42206
rect 7310 42130 7362 42142
rect 8654 42194 8706 42206
rect 8654 42130 8706 42142
rect 10782 42194 10834 42206
rect 10782 42130 10834 42142
rect 10894 42194 10946 42206
rect 10894 42130 10946 42142
rect 12126 42194 12178 42206
rect 12126 42130 12178 42142
rect 12238 42194 12290 42206
rect 12238 42130 12290 42142
rect 13134 42194 13186 42206
rect 13134 42130 13186 42142
rect 15150 42194 15202 42206
rect 23326 42194 23378 42206
rect 16594 42142 16606 42194
rect 16658 42142 16670 42194
rect 15150 42130 15202 42142
rect 23326 42130 23378 42142
rect 27582 42194 27634 42206
rect 27582 42130 27634 42142
rect 30046 42194 30098 42206
rect 30046 42130 30098 42142
rect 34190 42194 34242 42206
rect 34190 42130 34242 42142
rect 34862 42194 34914 42206
rect 34862 42130 34914 42142
rect 6862 42082 6914 42094
rect 3154 42030 3166 42082
rect 3218 42030 3230 42082
rect 4162 42030 4174 42082
rect 4226 42030 4238 42082
rect 4834 42030 4846 42082
rect 4898 42030 4910 42082
rect 5506 42030 5518 42082
rect 5570 42030 5582 42082
rect 6862 42018 6914 42030
rect 7086 42082 7138 42094
rect 7086 42018 7138 42030
rect 7422 42082 7474 42094
rect 7422 42018 7474 42030
rect 8318 42082 8370 42094
rect 8318 42018 8370 42030
rect 11006 42082 11058 42094
rect 11006 42018 11058 42030
rect 14366 42082 14418 42094
rect 14366 42018 14418 42030
rect 17726 42082 17778 42094
rect 17726 42018 17778 42030
rect 25790 42082 25842 42094
rect 25790 42018 25842 42030
rect 26014 42082 26066 42094
rect 26014 42018 26066 42030
rect 26462 42082 26514 42094
rect 26462 42018 26514 42030
rect 26686 42082 26738 42094
rect 26686 42018 26738 42030
rect 26910 42082 26962 42094
rect 26910 42018 26962 42030
rect 27022 42082 27074 42094
rect 27022 42018 27074 42030
rect 29486 42082 29538 42094
rect 29486 42018 29538 42030
rect 31838 42082 31890 42094
rect 31838 42018 31890 42030
rect 31950 42082 32002 42094
rect 31950 42018 32002 42030
rect 33742 42082 33794 42094
rect 33742 42018 33794 42030
rect 33966 42082 34018 42094
rect 33966 42018 34018 42030
rect 34302 42082 34354 42094
rect 34302 42018 34354 42030
rect 35758 42082 35810 42094
rect 35758 42018 35810 42030
rect 35870 42082 35922 42094
rect 35870 42018 35922 42030
rect 36542 42082 36594 42094
rect 36542 42018 36594 42030
rect 36878 42082 36930 42094
rect 36878 42018 36930 42030
rect 37438 42082 37490 42094
rect 37438 42018 37490 42030
rect 37774 42082 37826 42094
rect 37774 42018 37826 42030
rect 40238 42082 40290 42094
rect 40238 42018 40290 42030
rect 40686 42082 40738 42094
rect 40686 42018 40738 42030
rect 10334 41970 10386 41982
rect 4722 41918 4734 41970
rect 4786 41918 4798 41970
rect 5954 41918 5966 41970
rect 6018 41918 6030 41970
rect 6290 41918 6302 41970
rect 6354 41918 6366 41970
rect 10334 41906 10386 41918
rect 14030 41970 14082 41982
rect 14030 41906 14082 41918
rect 16046 41970 16098 41982
rect 16046 41906 16098 41918
rect 16942 41970 16994 41982
rect 22094 41970 22146 41982
rect 17938 41918 17950 41970
rect 18002 41918 18014 41970
rect 18834 41918 18846 41970
rect 18898 41918 18910 41970
rect 16942 41906 16994 41918
rect 22094 41906 22146 41918
rect 22542 41970 22594 41982
rect 22542 41906 22594 41918
rect 23102 41970 23154 41982
rect 23102 41906 23154 41918
rect 23774 41970 23826 41982
rect 23774 41906 23826 41918
rect 24670 41970 24722 41982
rect 24670 41906 24722 41918
rect 25678 41970 25730 41982
rect 28590 41970 28642 41982
rect 30382 41970 30434 41982
rect 27794 41918 27806 41970
rect 27858 41918 27870 41970
rect 28802 41918 28814 41970
rect 28866 41918 28878 41970
rect 25678 41906 25730 41918
rect 28590 41906 28642 41918
rect 30382 41906 30434 41918
rect 31614 41970 31666 41982
rect 32846 41970 32898 41982
rect 38670 41970 38722 41982
rect 32274 41918 32286 41970
rect 32338 41918 32350 41970
rect 35074 41918 35086 41970
rect 35138 41918 35150 41970
rect 31614 41906 31666 41918
rect 32846 41906 32898 41918
rect 38670 41906 38722 41918
rect 38894 41970 38946 41982
rect 38894 41906 38946 41918
rect 39118 41970 39170 41982
rect 39118 41906 39170 41918
rect 40462 41970 40514 41982
rect 40462 41906 40514 41918
rect 40798 41970 40850 41982
rect 40798 41906 40850 41918
rect 41470 41970 41522 41982
rect 41470 41906 41522 41918
rect 44158 41970 44210 41982
rect 44158 41906 44210 41918
rect 44382 41970 44434 41982
rect 44382 41906 44434 41918
rect 1934 41858 1986 41870
rect 1934 41794 1986 41806
rect 2382 41858 2434 41870
rect 2382 41794 2434 41806
rect 9886 41858 9938 41870
rect 9886 41794 9938 41806
rect 11454 41858 11506 41870
rect 11454 41794 11506 41806
rect 15598 41858 15650 41870
rect 19966 41858 20018 41870
rect 18946 41806 18958 41858
rect 19010 41806 19022 41858
rect 15598 41794 15650 41806
rect 19966 41794 20018 41806
rect 20302 41858 20354 41870
rect 20302 41794 20354 41806
rect 20750 41858 20802 41870
rect 20750 41794 20802 41806
rect 21198 41858 21250 41870
rect 21198 41794 21250 41806
rect 21758 41858 21810 41870
rect 21758 41794 21810 41806
rect 23214 41858 23266 41870
rect 23214 41794 23266 41806
rect 24558 41858 24610 41870
rect 24558 41794 24610 41806
rect 31054 41858 31106 41870
rect 32386 41806 32398 41858
rect 32450 41806 32462 41858
rect 31054 41794 31106 41806
rect 12350 41746 12402 41758
rect 9874 41694 9886 41746
rect 9938 41743 9950 41746
rect 10210 41743 10222 41746
rect 9938 41697 10222 41743
rect 9938 41694 9950 41697
rect 10210 41694 10222 41697
rect 10274 41694 10286 41746
rect 12350 41682 12402 41694
rect 12910 41746 12962 41758
rect 12910 41682 12962 41694
rect 13246 41746 13298 41758
rect 13246 41682 13298 41694
rect 13918 41746 13970 41758
rect 13918 41682 13970 41694
rect 14254 41746 14306 41758
rect 35870 41746 35922 41758
rect 19058 41694 19070 41746
rect 19122 41694 19134 41746
rect 20962 41694 20974 41746
rect 21026 41743 21038 41746
rect 21746 41743 21758 41746
rect 21026 41697 21758 41743
rect 21026 41694 21038 41697
rect 21746 41694 21758 41697
rect 21810 41694 21822 41746
rect 14254 41682 14306 41694
rect 35870 41682 35922 41694
rect 39342 41746 39394 41758
rect 39342 41682 39394 41694
rect 39790 41746 39842 41758
rect 39790 41682 39842 41694
rect 43486 41746 43538 41758
rect 43486 41682 43538 41694
rect 43934 41746 43986 41758
rect 43934 41682 43986 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 17614 41410 17666 41422
rect 14018 41358 14030 41410
rect 14082 41358 14094 41410
rect 17614 41346 17666 41358
rect 19854 41410 19906 41422
rect 19854 41346 19906 41358
rect 21870 41410 21922 41422
rect 21870 41346 21922 41358
rect 22206 41410 22258 41422
rect 22206 41346 22258 41358
rect 25454 41410 25506 41422
rect 25454 41346 25506 41358
rect 27582 41410 27634 41422
rect 27582 41346 27634 41358
rect 39566 41410 39618 41422
rect 39566 41346 39618 41358
rect 39790 41410 39842 41422
rect 39790 41346 39842 41358
rect 5966 41298 6018 41310
rect 25230 41298 25282 41310
rect 2258 41246 2270 41298
rect 2322 41246 2334 41298
rect 7970 41246 7982 41298
rect 8034 41246 8046 41298
rect 10658 41246 10670 41298
rect 10722 41246 10734 41298
rect 13906 41246 13918 41298
rect 13970 41246 13982 41298
rect 20626 41246 20638 41298
rect 20690 41246 20702 41298
rect 24098 41246 24110 41298
rect 24162 41246 24174 41298
rect 5966 41234 6018 41246
rect 25230 41234 25282 41246
rect 26350 41298 26402 41310
rect 26350 41234 26402 41246
rect 32846 41298 32898 41310
rect 32846 41234 32898 41246
rect 35534 41298 35586 41310
rect 35534 41234 35586 41246
rect 36318 41298 36370 41310
rect 36318 41234 36370 41246
rect 38446 41298 38498 41310
rect 38446 41234 38498 41246
rect 39006 41298 39058 41310
rect 55346 41246 55358 41298
rect 55410 41246 55422 41298
rect 39006 41234 39058 41246
rect 4622 41186 4674 41198
rect 9662 41186 9714 41198
rect 11790 41186 11842 41198
rect 7522 41134 7534 41186
rect 7586 41134 7598 41186
rect 8418 41134 8430 41186
rect 8482 41134 8494 41186
rect 9874 41134 9886 41186
rect 9938 41134 9950 41186
rect 10770 41134 10782 41186
rect 10834 41134 10846 41186
rect 4622 41122 4674 41134
rect 9662 41122 9714 41134
rect 11790 41122 11842 41134
rect 12126 41186 12178 41198
rect 17278 41186 17330 41198
rect 14018 41134 14030 41186
rect 14082 41134 14094 41186
rect 14242 41134 14254 41186
rect 14306 41134 14318 41186
rect 16482 41134 16494 41186
rect 16546 41134 16558 41186
rect 12126 41122 12178 41134
rect 17278 41122 17330 41134
rect 20078 41186 20130 41198
rect 20750 41186 20802 41198
rect 28254 41186 28306 41198
rect 20402 41134 20414 41186
rect 20466 41134 20478 41186
rect 22978 41134 22990 41186
rect 23042 41134 23054 41186
rect 23762 41134 23774 41186
rect 23826 41134 23838 41186
rect 20078 41122 20130 41134
rect 20750 41122 20802 41134
rect 28254 41122 28306 41134
rect 28478 41186 28530 41198
rect 28478 41122 28530 41134
rect 29822 41186 29874 41198
rect 29822 41122 29874 41134
rect 32174 41186 32226 41198
rect 32174 41122 32226 41134
rect 32510 41186 32562 41198
rect 39230 41186 39282 41198
rect 37762 41134 37774 41186
rect 37826 41134 37838 41186
rect 32510 41122 32562 41134
rect 39230 41122 39282 41134
rect 42926 41186 42978 41198
rect 42926 41122 42978 41134
rect 43710 41186 43762 41198
rect 43710 41122 43762 41134
rect 43822 41186 43874 41198
rect 43822 41122 43874 41134
rect 45726 41186 45778 41198
rect 45726 41122 45778 41134
rect 46062 41186 46114 41198
rect 56130 41134 56142 41186
rect 56194 41134 56206 41186
rect 46062 41122 46114 41134
rect 2494 41074 2546 41086
rect 4062 41074 4114 41086
rect 12014 41074 12066 41086
rect 19294 41074 19346 41086
rect 3378 41022 3390 41074
rect 3442 41022 3454 41074
rect 4946 41022 4958 41074
rect 5010 41022 5022 41074
rect 7298 41022 7310 41074
rect 7362 41022 7374 41074
rect 11106 41022 11118 41074
rect 11170 41022 11182 41074
rect 16594 41022 16606 41074
rect 16658 41022 16670 41074
rect 18834 41022 18846 41074
rect 18898 41022 18910 41074
rect 2494 41010 2546 41022
rect 4062 41010 4114 41022
rect 12014 41010 12066 41022
rect 19294 41010 19346 41022
rect 21646 41074 21698 41086
rect 27694 41074 27746 41086
rect 24210 41022 24222 41074
rect 24274 41022 24286 41074
rect 25778 41022 25790 41074
rect 25842 41022 25854 41074
rect 21646 41010 21698 41022
rect 27694 41010 27746 41022
rect 32286 41074 32338 41086
rect 32286 41010 32338 41022
rect 37998 41074 38050 41086
rect 37998 41010 38050 41022
rect 40462 41074 40514 41086
rect 40462 41010 40514 41022
rect 40574 41074 40626 41086
rect 40574 41010 40626 41022
rect 43038 41074 43090 41086
rect 43038 41010 43090 41022
rect 44158 41074 44210 41086
rect 44158 41010 44210 41022
rect 45502 41074 45554 41086
rect 45502 41010 45554 41022
rect 2270 40962 2322 40974
rect 2270 40898 2322 40910
rect 3054 40962 3106 40974
rect 3054 40898 3106 40910
rect 12910 40962 12962 40974
rect 12910 40898 12962 40910
rect 15486 40962 15538 40974
rect 15486 40898 15538 40910
rect 15934 40962 15986 40974
rect 15934 40898 15986 40910
rect 18510 40962 18562 40974
rect 18510 40898 18562 40910
rect 20526 40962 20578 40974
rect 20526 40898 20578 40910
rect 23102 40962 23154 40974
rect 23102 40898 23154 40910
rect 27134 40962 27186 40974
rect 29598 40962 29650 40974
rect 28802 40910 28814 40962
rect 28866 40910 28878 40962
rect 27134 40898 27186 40910
rect 29598 40898 29650 40910
rect 29710 40962 29762 40974
rect 29710 40898 29762 40910
rect 30046 40962 30098 40974
rect 30046 40898 30098 40910
rect 30606 40962 30658 40974
rect 30606 40898 30658 40910
rect 31054 40962 31106 40974
rect 31054 40898 31106 40910
rect 39902 40962 39954 40974
rect 39902 40898 39954 40910
rect 40798 40962 40850 40974
rect 40798 40898 40850 40910
rect 43262 40962 43314 40974
rect 43262 40898 43314 40910
rect 43934 40962 43986 40974
rect 43934 40898 43986 40910
rect 45726 40962 45778 40974
rect 45726 40898 45778 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 1822 40626 1874 40638
rect 1822 40562 1874 40574
rect 8766 40626 8818 40638
rect 8766 40562 8818 40574
rect 8878 40626 8930 40638
rect 8878 40562 8930 40574
rect 10110 40626 10162 40638
rect 10110 40562 10162 40574
rect 10670 40626 10722 40638
rect 10670 40562 10722 40574
rect 12238 40626 12290 40638
rect 12238 40562 12290 40574
rect 13134 40626 13186 40638
rect 13134 40562 13186 40574
rect 13694 40626 13746 40638
rect 13694 40562 13746 40574
rect 16606 40626 16658 40638
rect 16606 40562 16658 40574
rect 17614 40626 17666 40638
rect 17614 40562 17666 40574
rect 17838 40626 17890 40638
rect 17838 40562 17890 40574
rect 20414 40626 20466 40638
rect 20414 40562 20466 40574
rect 21422 40626 21474 40638
rect 21422 40562 21474 40574
rect 21982 40626 22034 40638
rect 21982 40562 22034 40574
rect 24110 40626 24162 40638
rect 24110 40562 24162 40574
rect 24558 40626 24610 40638
rect 24558 40562 24610 40574
rect 26350 40626 26402 40638
rect 26350 40562 26402 40574
rect 26798 40626 26850 40638
rect 26798 40562 26850 40574
rect 27358 40626 27410 40638
rect 27358 40562 27410 40574
rect 28030 40626 28082 40638
rect 28030 40562 28082 40574
rect 28478 40626 28530 40638
rect 28478 40562 28530 40574
rect 28926 40626 28978 40638
rect 28926 40562 28978 40574
rect 34974 40626 35026 40638
rect 38670 40626 38722 40638
rect 36530 40574 36542 40626
rect 36594 40574 36606 40626
rect 34974 40562 35026 40574
rect 38670 40562 38722 40574
rect 40014 40626 40066 40638
rect 40014 40562 40066 40574
rect 40798 40626 40850 40638
rect 40798 40562 40850 40574
rect 43934 40626 43986 40638
rect 44930 40574 44942 40626
rect 44994 40574 45006 40626
rect 43934 40562 43986 40574
rect 7086 40514 7138 40526
rect 12910 40514 12962 40526
rect 2930 40462 2942 40514
rect 2994 40462 3006 40514
rect 8418 40462 8430 40514
rect 8482 40462 8494 40514
rect 7086 40450 7138 40462
rect 12910 40450 12962 40462
rect 17950 40514 18002 40526
rect 17950 40450 18002 40462
rect 20078 40514 20130 40526
rect 20078 40450 20130 40462
rect 22430 40514 22482 40526
rect 22430 40450 22482 40462
rect 23438 40514 23490 40526
rect 23438 40450 23490 40462
rect 29374 40514 29426 40526
rect 29374 40450 29426 40462
rect 31166 40514 31218 40526
rect 31166 40450 31218 40462
rect 33966 40514 34018 40526
rect 33966 40450 34018 40462
rect 34638 40514 34690 40526
rect 34638 40450 34690 40462
rect 37774 40514 37826 40526
rect 37774 40450 37826 40462
rect 43710 40514 43762 40526
rect 44482 40462 44494 40514
rect 44546 40462 44558 40514
rect 43710 40450 43762 40462
rect 2270 40402 2322 40414
rect 8990 40402 9042 40414
rect 3938 40350 3950 40402
rect 4002 40350 4014 40402
rect 4498 40350 4510 40402
rect 4562 40350 4574 40402
rect 5842 40350 5854 40402
rect 5906 40350 5918 40402
rect 8530 40350 8542 40402
rect 8594 40350 8606 40402
rect 2270 40338 2322 40350
rect 8990 40338 9042 40350
rect 9774 40402 9826 40414
rect 9774 40338 9826 40350
rect 11230 40402 11282 40414
rect 11230 40338 11282 40350
rect 11566 40402 11618 40414
rect 11566 40338 11618 40350
rect 12798 40402 12850 40414
rect 15822 40402 15874 40414
rect 15362 40350 15374 40402
rect 15426 40350 15438 40402
rect 12798 40338 12850 40350
rect 15822 40338 15874 40350
rect 16942 40402 16994 40414
rect 16942 40338 16994 40350
rect 19070 40402 19122 40414
rect 19070 40338 19122 40350
rect 20414 40402 20466 40414
rect 20414 40338 20466 40350
rect 20638 40402 20690 40414
rect 20638 40338 20690 40350
rect 22094 40402 22146 40414
rect 22094 40338 22146 40350
rect 22206 40402 22258 40414
rect 23550 40402 23602 40414
rect 23090 40350 23102 40402
rect 23154 40350 23166 40402
rect 22206 40338 22258 40350
rect 23550 40338 23602 40350
rect 23662 40402 23714 40414
rect 23662 40338 23714 40350
rect 29598 40402 29650 40414
rect 29598 40338 29650 40350
rect 29822 40402 29874 40414
rect 29822 40338 29874 40350
rect 33854 40402 33906 40414
rect 33854 40338 33906 40350
rect 36878 40402 36930 40414
rect 36878 40338 36930 40350
rect 37438 40402 37490 40414
rect 37438 40338 37490 40350
rect 41582 40402 41634 40414
rect 41582 40338 41634 40350
rect 41806 40402 41858 40414
rect 43598 40402 43650 40414
rect 46622 40402 46674 40414
rect 42130 40350 42142 40402
rect 42194 40350 42206 40402
rect 44370 40350 44382 40402
rect 44434 40350 44446 40402
rect 45378 40350 45390 40402
rect 45442 40350 45454 40402
rect 46834 40350 46846 40402
rect 46898 40350 46910 40402
rect 41806 40338 41858 40350
rect 43598 40338 43650 40350
rect 46622 40338 46674 40350
rect 7198 40290 7250 40302
rect 3042 40238 3054 40290
rect 3106 40238 3118 40290
rect 7198 40226 7250 40238
rect 14590 40290 14642 40302
rect 18734 40290 18786 40302
rect 15138 40238 15150 40290
rect 15202 40238 15214 40290
rect 14590 40226 14642 40238
rect 18734 40226 18786 40238
rect 19518 40290 19570 40302
rect 19518 40226 19570 40238
rect 26014 40290 26066 40302
rect 26014 40226 26066 40238
rect 29486 40290 29538 40302
rect 29486 40226 29538 40238
rect 45166 40290 45218 40302
rect 45166 40226 45218 40238
rect 47518 40290 47570 40302
rect 47518 40226 47570 40238
rect 7310 40178 7362 40190
rect 7310 40114 7362 40126
rect 11118 40178 11170 40190
rect 11118 40114 11170 40126
rect 11454 40178 11506 40190
rect 11454 40114 11506 40126
rect 13582 40178 13634 40190
rect 13582 40114 13634 40126
rect 13918 40178 13970 40190
rect 33966 40178 34018 40190
rect 23874 40126 23886 40178
rect 23938 40175 23950 40178
rect 24210 40175 24222 40178
rect 23938 40129 24222 40175
rect 23938 40126 23950 40129
rect 24210 40126 24222 40129
rect 24274 40126 24286 40178
rect 26114 40126 26126 40178
rect 26178 40175 26190 40178
rect 27234 40175 27246 40178
rect 26178 40129 27246 40175
rect 26178 40126 26190 40129
rect 27234 40126 27246 40129
rect 27298 40126 27310 40178
rect 13918 40114 13970 40126
rect 33966 40114 34018 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 16942 39842 16994 39854
rect 7522 39790 7534 39842
rect 7586 39839 7598 39842
rect 7746 39839 7758 39842
rect 7586 39793 7758 39839
rect 7586 39790 7598 39793
rect 7746 39790 7758 39793
rect 7810 39790 7822 39842
rect 14242 39790 14254 39842
rect 14306 39790 14318 39842
rect 16942 39778 16994 39790
rect 17502 39842 17554 39854
rect 17502 39778 17554 39790
rect 19854 39842 19906 39854
rect 19854 39778 19906 39790
rect 20190 39842 20242 39854
rect 20190 39778 20242 39790
rect 22094 39842 22146 39854
rect 22094 39778 22146 39790
rect 23102 39842 23154 39854
rect 23102 39778 23154 39790
rect 30942 39842 30994 39854
rect 30942 39778 30994 39790
rect 37550 39842 37602 39854
rect 37550 39778 37602 39790
rect 3726 39730 3778 39742
rect 3726 39666 3778 39678
rect 5966 39730 6018 39742
rect 5966 39666 6018 39678
rect 7534 39730 7586 39742
rect 7534 39666 7586 39678
rect 8990 39730 9042 39742
rect 8990 39666 9042 39678
rect 10446 39730 10498 39742
rect 10446 39666 10498 39678
rect 12462 39730 12514 39742
rect 12462 39666 12514 39678
rect 12910 39730 12962 39742
rect 12910 39666 12962 39678
rect 15038 39730 15090 39742
rect 15038 39666 15090 39678
rect 21646 39730 21698 39742
rect 25006 39730 25058 39742
rect 24210 39678 24222 39730
rect 24274 39678 24286 39730
rect 21646 39666 21698 39678
rect 25006 39666 25058 39678
rect 25454 39730 25506 39742
rect 25454 39666 25506 39678
rect 25902 39730 25954 39742
rect 25902 39666 25954 39678
rect 33630 39730 33682 39742
rect 33630 39666 33682 39678
rect 36878 39730 36930 39742
rect 36878 39666 36930 39678
rect 37662 39730 37714 39742
rect 43710 39730 43762 39742
rect 40674 39678 40686 39730
rect 40738 39678 40750 39730
rect 43922 39678 43934 39730
rect 43986 39678 43998 39730
rect 37662 39666 37714 39678
rect 43710 39666 43762 39678
rect 3502 39618 3554 39630
rect 2818 39566 2830 39618
rect 2882 39566 2894 39618
rect 3502 39554 3554 39566
rect 3838 39618 3890 39630
rect 3838 39554 3890 39566
rect 4174 39618 4226 39630
rect 4174 39554 4226 39566
rect 7982 39618 8034 39630
rect 7982 39554 8034 39566
rect 9550 39618 9602 39630
rect 9550 39554 9602 39566
rect 9998 39618 10050 39630
rect 9998 39554 10050 39566
rect 10222 39618 10274 39630
rect 10222 39554 10274 39566
rect 11118 39618 11170 39630
rect 11118 39554 11170 39566
rect 11342 39618 11394 39630
rect 17054 39618 17106 39630
rect 11666 39566 11678 39618
rect 11730 39566 11742 39618
rect 13906 39566 13918 39618
rect 13970 39566 13982 39618
rect 14242 39566 14254 39618
rect 14306 39566 14318 39618
rect 11342 39554 11394 39566
rect 17054 39554 17106 39566
rect 17726 39618 17778 39630
rect 17726 39554 17778 39566
rect 18398 39618 18450 39630
rect 18398 39554 18450 39566
rect 21870 39618 21922 39630
rect 21870 39554 21922 39566
rect 22542 39618 22594 39630
rect 22542 39554 22594 39566
rect 22990 39618 23042 39630
rect 31502 39618 31554 39630
rect 33742 39618 33794 39630
rect 39342 39618 39394 39630
rect 47518 39618 47570 39630
rect 26450 39566 26462 39618
rect 26514 39566 26526 39618
rect 27234 39566 27246 39618
rect 27298 39566 27310 39618
rect 27682 39566 27694 39618
rect 27746 39566 27758 39618
rect 32610 39566 32622 39618
rect 32674 39566 32686 39618
rect 34178 39566 34190 39618
rect 34242 39566 34254 39618
rect 38882 39566 38894 39618
rect 38946 39566 38958 39618
rect 40562 39566 40574 39618
rect 40626 39566 40638 39618
rect 42018 39566 42030 39618
rect 42082 39566 42094 39618
rect 44034 39566 44046 39618
rect 44098 39566 44110 39618
rect 57362 39566 57374 39618
rect 57426 39566 57438 39618
rect 22990 39554 23042 39566
rect 31502 39554 31554 39566
rect 33742 39554 33794 39566
rect 39342 39554 39394 39566
rect 47518 39554 47570 39566
rect 9102 39506 9154 39518
rect 1922 39454 1934 39506
rect 1986 39454 1998 39506
rect 6850 39454 6862 39506
rect 6914 39454 6926 39506
rect 8306 39454 8318 39506
rect 8370 39454 8382 39506
rect 9102 39442 9154 39454
rect 10558 39506 10610 39518
rect 10558 39442 10610 39454
rect 13694 39506 13746 39518
rect 13694 39442 13746 39454
rect 15934 39506 15986 39518
rect 19630 39506 19682 39518
rect 18722 39454 18734 39506
rect 18786 39454 18798 39506
rect 15934 39442 15986 39454
rect 19630 39442 19682 39454
rect 26686 39506 26738 39518
rect 26686 39442 26738 39454
rect 27806 39506 27858 39518
rect 27806 39442 27858 39454
rect 30830 39506 30882 39518
rect 57150 39506 57202 39518
rect 31826 39454 31838 39506
rect 31890 39454 31902 39506
rect 42466 39454 42478 39506
rect 42530 39454 42542 39506
rect 30830 39442 30882 39454
rect 57150 39442 57202 39454
rect 4958 39394 5010 39406
rect 4958 39330 5010 39342
rect 6526 39394 6578 39406
rect 6526 39330 6578 39342
rect 8878 39394 8930 39406
rect 8878 39330 8930 39342
rect 11230 39394 11282 39406
rect 11230 39330 11282 39342
rect 14478 39394 14530 39406
rect 14478 39330 14530 39342
rect 15598 39394 15650 39406
rect 15598 39330 15650 39342
rect 16494 39394 16546 39406
rect 16494 39330 16546 39342
rect 17838 39394 17890 39406
rect 17838 39330 17890 39342
rect 20974 39394 21026 39406
rect 20974 39330 21026 39342
rect 23102 39394 23154 39406
rect 23102 39330 23154 39342
rect 23774 39394 23826 39406
rect 23774 39330 23826 39342
rect 28366 39394 28418 39406
rect 28366 39330 28418 39342
rect 28814 39394 28866 39406
rect 28814 39330 28866 39342
rect 29934 39394 29986 39406
rect 29934 39330 29986 39342
rect 30382 39394 30434 39406
rect 30382 39330 30434 39342
rect 32398 39394 32450 39406
rect 32398 39330 32450 39342
rect 35086 39394 35138 39406
rect 35086 39330 35138 39342
rect 38110 39394 38162 39406
rect 38110 39330 38162 39342
rect 39230 39394 39282 39406
rect 39230 39330 39282 39342
rect 39454 39394 39506 39406
rect 39454 39330 39506 39342
rect 47854 39394 47906 39406
rect 47854 39330 47906 39342
rect 56702 39394 56754 39406
rect 56702 39330 56754 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 2158 39058 2210 39070
rect 2158 38994 2210 39006
rect 7758 39058 7810 39070
rect 7758 38994 7810 39006
rect 8094 39058 8146 39070
rect 8094 38994 8146 39006
rect 9998 39058 10050 39070
rect 9998 38994 10050 39006
rect 12350 39058 12402 39070
rect 12350 38994 12402 39006
rect 12574 39058 12626 39070
rect 12574 38994 12626 39006
rect 13358 39058 13410 39070
rect 13358 38994 13410 39006
rect 15710 39058 15762 39070
rect 15710 38994 15762 39006
rect 30046 39058 30098 39070
rect 30046 38994 30098 39006
rect 30494 39058 30546 39070
rect 39454 39058 39506 39070
rect 38882 39006 38894 39058
rect 38946 39006 38958 39058
rect 30494 38994 30546 39006
rect 39454 38994 39506 39006
rect 41694 39058 41746 39070
rect 41694 38994 41746 39006
rect 41918 39058 41970 39070
rect 41918 38994 41970 39006
rect 42814 39058 42866 39070
rect 42814 38994 42866 39006
rect 3838 38946 3890 38958
rect 7982 38946 8034 38958
rect 6066 38894 6078 38946
rect 6130 38894 6142 38946
rect 3838 38882 3890 38894
rect 7982 38882 8034 38894
rect 10110 38946 10162 38958
rect 10110 38882 10162 38894
rect 10782 38946 10834 38958
rect 10782 38882 10834 38894
rect 11118 38946 11170 38958
rect 11118 38882 11170 38894
rect 14254 38946 14306 38958
rect 14254 38882 14306 38894
rect 14590 38946 14642 38958
rect 14590 38882 14642 38894
rect 16382 38946 16434 38958
rect 16382 38882 16434 38894
rect 16494 38946 16546 38958
rect 16494 38882 16546 38894
rect 23214 38946 23266 38958
rect 23214 38882 23266 38894
rect 27806 38946 27858 38958
rect 27806 38882 27858 38894
rect 28702 38946 28754 38958
rect 28702 38882 28754 38894
rect 32510 38946 32562 38958
rect 36990 38946 37042 38958
rect 34626 38894 34638 38946
rect 34690 38894 34702 38946
rect 32510 38882 32562 38894
rect 36990 38882 37042 38894
rect 37214 38946 37266 38958
rect 37214 38882 37266 38894
rect 38334 38946 38386 38958
rect 38334 38882 38386 38894
rect 41582 38946 41634 38958
rect 41582 38882 41634 38894
rect 42478 38946 42530 38958
rect 42478 38882 42530 38894
rect 42590 38946 42642 38958
rect 42590 38882 42642 38894
rect 7422 38834 7474 38846
rect 1922 38782 1934 38834
rect 1986 38782 1998 38834
rect 3154 38782 3166 38834
rect 3218 38782 3230 38834
rect 5730 38782 5742 38834
rect 5794 38782 5806 38834
rect 6290 38782 6302 38834
rect 6354 38782 6366 38834
rect 6738 38782 6750 38834
rect 6802 38782 6814 38834
rect 7422 38770 7474 38782
rect 8654 38834 8706 38846
rect 8654 38770 8706 38782
rect 12686 38834 12738 38846
rect 12686 38770 12738 38782
rect 13694 38834 13746 38846
rect 24222 38834 24274 38846
rect 25790 38834 25842 38846
rect 27694 38834 27746 38846
rect 16146 38782 16158 38834
rect 16210 38782 16222 38834
rect 16930 38782 16942 38834
rect 16994 38782 17006 38834
rect 17714 38782 17726 38834
rect 17778 38782 17790 38834
rect 18050 38782 18062 38834
rect 18114 38782 18126 38834
rect 19618 38782 19630 38834
rect 19682 38782 19694 38834
rect 20738 38782 20750 38834
rect 20802 38782 20814 38834
rect 23762 38782 23774 38834
rect 23826 38782 23838 38834
rect 24546 38782 24558 38834
rect 24610 38782 24622 38834
rect 27346 38782 27358 38834
rect 27410 38782 27422 38834
rect 13694 38770 13746 38782
rect 24222 38770 24274 38782
rect 25790 38770 25842 38782
rect 27694 38770 27746 38782
rect 28366 38834 28418 38846
rect 28366 38770 28418 38782
rect 28478 38834 28530 38846
rect 28478 38770 28530 38782
rect 28814 38834 28866 38846
rect 28814 38770 28866 38782
rect 31054 38834 31106 38846
rect 31054 38770 31106 38782
rect 32622 38834 32674 38846
rect 36206 38834 36258 38846
rect 35522 38782 35534 38834
rect 35586 38782 35598 38834
rect 32622 38770 32674 38782
rect 36206 38770 36258 38782
rect 36878 38834 36930 38846
rect 36878 38770 36930 38782
rect 40014 38834 40066 38846
rect 40014 38770 40066 38782
rect 5182 38722 5234 38734
rect 2818 38670 2830 38722
rect 2882 38670 2894 38722
rect 4274 38670 4286 38722
rect 4338 38670 4350 38722
rect 5182 38658 5234 38670
rect 9102 38722 9154 38734
rect 9102 38658 9154 38670
rect 9886 38722 9938 38734
rect 9886 38658 9938 38670
rect 12014 38722 12066 38734
rect 12014 38658 12066 38670
rect 15262 38722 15314 38734
rect 22654 38722 22706 38734
rect 26350 38722 26402 38734
rect 21410 38670 21422 38722
rect 21474 38670 21486 38722
rect 24658 38670 24670 38722
rect 24722 38670 24734 38722
rect 15262 38658 15314 38670
rect 22654 38658 22706 38670
rect 26350 38658 26402 38670
rect 29598 38722 29650 38734
rect 34190 38722 34242 38734
rect 31378 38670 31390 38722
rect 31442 38670 31454 38722
rect 29598 38658 29650 38670
rect 34190 38658 34242 38670
rect 37662 38722 37714 38734
rect 37662 38658 37714 38670
rect 39566 38722 39618 38734
rect 39566 38658 39618 38670
rect 40462 38722 40514 38734
rect 40462 38658 40514 38670
rect 38558 38610 38610 38622
rect 21634 38558 21646 38610
rect 21698 38558 21710 38610
rect 31266 38558 31278 38610
rect 31330 38558 31342 38610
rect 38558 38546 38610 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 23662 38274 23714 38286
rect 26686 38274 26738 38286
rect 1810 38222 1822 38274
rect 1874 38271 1886 38274
rect 2258 38271 2270 38274
rect 1874 38225 2270 38271
rect 1874 38222 1886 38225
rect 2258 38222 2270 38225
rect 2322 38271 2334 38274
rect 2594 38271 2606 38274
rect 2322 38225 2606 38271
rect 2322 38222 2334 38225
rect 2594 38222 2606 38225
rect 2658 38222 2670 38274
rect 24210 38222 24222 38274
rect 24274 38271 24286 38274
rect 24546 38271 24558 38274
rect 24274 38225 24558 38271
rect 24274 38222 24286 38225
rect 24546 38222 24558 38225
rect 24610 38222 24622 38274
rect 23662 38210 23714 38222
rect 26686 38210 26738 38222
rect 31054 38274 31106 38286
rect 31054 38210 31106 38222
rect 31502 38274 31554 38286
rect 31502 38210 31554 38222
rect 32286 38274 32338 38286
rect 34178 38222 34190 38274
rect 34242 38271 34254 38274
rect 34514 38271 34526 38274
rect 34242 38225 34526 38271
rect 34242 38222 34254 38225
rect 34514 38222 34526 38225
rect 34578 38271 34590 38274
rect 35074 38271 35086 38274
rect 34578 38225 35086 38271
rect 34578 38222 34590 38225
rect 35074 38222 35086 38225
rect 35138 38222 35150 38274
rect 32286 38210 32338 38222
rect 1934 38162 1986 38174
rect 5070 38162 5122 38174
rect 18622 38162 18674 38174
rect 3266 38110 3278 38162
rect 3330 38110 3342 38162
rect 9986 38110 9998 38162
rect 10050 38110 10062 38162
rect 14466 38110 14478 38162
rect 14530 38110 14542 38162
rect 1934 38098 1986 38110
rect 5070 38098 5122 38110
rect 18622 38098 18674 38110
rect 18734 38162 18786 38174
rect 23214 38162 23266 38174
rect 20626 38110 20638 38162
rect 20690 38110 20702 38162
rect 22082 38110 22094 38162
rect 22146 38110 22158 38162
rect 18734 38098 18786 38110
rect 23214 38098 23266 38110
rect 23438 38162 23490 38174
rect 23438 38098 23490 38110
rect 24110 38162 24162 38174
rect 24110 38098 24162 38110
rect 28814 38162 28866 38174
rect 33518 38162 33570 38174
rect 31938 38110 31950 38162
rect 32002 38110 32014 38162
rect 28814 38098 28866 38110
rect 33518 38098 33570 38110
rect 34526 38162 34578 38174
rect 34526 38098 34578 38110
rect 34974 38162 35026 38174
rect 34974 38098 35026 38110
rect 36766 38162 36818 38174
rect 37986 38110 37998 38162
rect 38050 38110 38062 38162
rect 41906 38110 41918 38162
rect 41970 38110 41982 38162
rect 36766 38098 36818 38110
rect 2830 38050 2882 38062
rect 11790 38050 11842 38062
rect 24446 38050 24498 38062
rect 26574 38050 26626 38062
rect 5842 37998 5854 38050
rect 5906 37998 5918 38050
rect 7074 37998 7086 38050
rect 7138 37998 7150 38050
rect 7522 37998 7534 38050
rect 7586 37998 7598 38050
rect 9090 37998 9102 38050
rect 9154 37998 9166 38050
rect 14018 37998 14030 38050
rect 14082 37998 14094 38050
rect 14914 37998 14926 38050
rect 14978 37998 14990 38050
rect 20290 37998 20302 38050
rect 20354 37998 20366 38050
rect 25554 37998 25566 38050
rect 25618 37998 25630 38050
rect 2830 37986 2882 37998
rect 11790 37986 11842 37998
rect 24446 37986 24498 37998
rect 26574 37986 26626 37998
rect 27358 38050 27410 38062
rect 29598 38050 29650 38062
rect 27570 37998 27582 38050
rect 27634 37998 27646 38050
rect 27358 37986 27410 37998
rect 29598 37986 29650 37998
rect 30046 38050 30098 38062
rect 30046 37986 30098 37998
rect 30606 38050 30658 38062
rect 30606 37986 30658 37998
rect 30830 38050 30882 38062
rect 30830 37986 30882 37998
rect 33070 38050 33122 38062
rect 33070 37986 33122 37998
rect 33966 38050 34018 38062
rect 42142 38050 42194 38062
rect 39442 37998 39454 38050
rect 39506 37998 39518 38050
rect 33966 37986 34018 37998
rect 42142 37986 42194 37998
rect 42366 38050 42418 38062
rect 42366 37986 42418 37998
rect 2382 37938 2434 37950
rect 2382 37874 2434 37886
rect 4286 37938 4338 37950
rect 12686 37938 12738 37950
rect 16046 37938 16098 37950
rect 6402 37886 6414 37938
rect 6466 37886 6478 37938
rect 10098 37886 10110 37938
rect 10162 37886 10174 37938
rect 14354 37886 14366 37938
rect 14418 37886 14430 37938
rect 4286 37874 4338 37886
rect 12686 37874 12738 37886
rect 16046 37874 16098 37886
rect 16494 37938 16546 37950
rect 16494 37874 16546 37886
rect 16942 37938 16994 37950
rect 16942 37874 16994 37886
rect 17502 37938 17554 37950
rect 17502 37874 17554 37886
rect 19294 37938 19346 37950
rect 19294 37874 19346 37886
rect 19630 37938 19682 37950
rect 21646 37938 21698 37950
rect 20850 37886 20862 37938
rect 20914 37886 20926 37938
rect 19630 37874 19682 37886
rect 21646 37874 21698 37886
rect 22654 37938 22706 37950
rect 22654 37874 22706 37886
rect 28254 37938 28306 37950
rect 28254 37874 28306 37886
rect 32062 37938 32114 37950
rect 32062 37874 32114 37886
rect 32958 37938 33010 37950
rect 40126 37938 40178 37950
rect 38210 37886 38222 37938
rect 38274 37886 38286 37938
rect 32958 37874 33010 37886
rect 40126 37874 40178 37886
rect 41582 37938 41634 37950
rect 41582 37874 41634 37886
rect 41806 37938 41858 37950
rect 41806 37874 41858 37886
rect 3950 37826 4002 37838
rect 11230 37826 11282 37838
rect 5842 37774 5854 37826
rect 5906 37774 5918 37826
rect 3950 37762 4002 37774
rect 11230 37762 11282 37774
rect 12350 37826 12402 37838
rect 12350 37762 12402 37774
rect 15710 37826 15762 37838
rect 15710 37762 15762 37774
rect 17838 37826 17890 37838
rect 17838 37762 17890 37774
rect 18510 37826 18562 37838
rect 18510 37762 18562 37774
rect 24894 37826 24946 37838
rect 24894 37762 24946 37774
rect 25790 37826 25842 37838
rect 25790 37762 25842 37774
rect 26462 37826 26514 37838
rect 26462 37762 26514 37774
rect 32734 37826 32786 37838
rect 32734 37762 32786 37774
rect 41134 37826 41186 37838
rect 41134 37762 41186 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 2158 37490 2210 37502
rect 2158 37426 2210 37438
rect 3838 37490 3890 37502
rect 3838 37426 3890 37438
rect 4398 37490 4450 37502
rect 4398 37426 4450 37438
rect 9886 37490 9938 37502
rect 9886 37426 9938 37438
rect 14702 37490 14754 37502
rect 21534 37490 21586 37502
rect 16930 37438 16942 37490
rect 16994 37438 17006 37490
rect 14702 37426 14754 37438
rect 21534 37426 21586 37438
rect 22206 37490 22258 37502
rect 37550 37490 37602 37502
rect 22530 37438 22542 37490
rect 22594 37438 22606 37490
rect 27234 37438 27246 37490
rect 27298 37438 27310 37490
rect 27794 37438 27806 37490
rect 27858 37438 27870 37490
rect 38658 37438 38670 37490
rect 38722 37438 38734 37490
rect 22206 37426 22258 37438
rect 37550 37426 37602 37438
rect 1822 37378 1874 37390
rect 1822 37314 1874 37326
rect 7198 37378 7250 37390
rect 7198 37314 7250 37326
rect 8990 37378 9042 37390
rect 21422 37378 21474 37390
rect 10546 37326 10558 37378
rect 10610 37326 10622 37378
rect 14466 37326 14478 37378
rect 14530 37326 14542 37378
rect 8990 37314 9042 37326
rect 21422 37314 21474 37326
rect 21646 37378 21698 37390
rect 34414 37378 34466 37390
rect 23202 37326 23214 37378
rect 23266 37326 23278 37378
rect 21646 37314 21698 37326
rect 34414 37314 34466 37326
rect 34750 37378 34802 37390
rect 34750 37314 34802 37326
rect 35422 37378 35474 37390
rect 35422 37314 35474 37326
rect 2718 37266 2770 37278
rect 2718 37202 2770 37214
rect 3278 37266 3330 37278
rect 3278 37202 3330 37214
rect 4286 37266 4338 37278
rect 4286 37202 4338 37214
rect 4510 37266 4562 37278
rect 5742 37266 5794 37278
rect 4834 37214 4846 37266
rect 4898 37214 4910 37266
rect 4510 37202 4562 37214
rect 5742 37202 5794 37214
rect 6302 37266 6354 37278
rect 6302 37202 6354 37214
rect 6974 37266 7026 37278
rect 6974 37202 7026 37214
rect 7422 37266 7474 37278
rect 15150 37266 15202 37278
rect 8754 37214 8766 37266
rect 8818 37214 8830 37266
rect 10882 37214 10894 37266
rect 10946 37214 10958 37266
rect 12226 37214 12238 37266
rect 12290 37214 12302 37266
rect 14242 37214 14254 37266
rect 14306 37214 14318 37266
rect 7422 37202 7474 37214
rect 15150 37202 15202 37214
rect 15374 37266 15426 37278
rect 15374 37202 15426 37214
rect 16606 37266 16658 37278
rect 26238 37266 26290 37278
rect 18386 37214 18398 37266
rect 18450 37214 18462 37266
rect 18610 37214 18622 37266
rect 18674 37214 18686 37266
rect 20066 37214 20078 37266
rect 20130 37214 20142 37266
rect 23538 37214 23550 37266
rect 23602 37214 23614 37266
rect 24210 37214 24222 37266
rect 24274 37214 24286 37266
rect 16606 37202 16658 37214
rect 26238 37202 26290 37214
rect 26686 37266 26738 37278
rect 26686 37202 26738 37214
rect 28142 37266 28194 37278
rect 30606 37266 30658 37278
rect 29586 37214 29598 37266
rect 29650 37214 29662 37266
rect 28142 37202 28194 37214
rect 30606 37202 30658 37214
rect 31950 37266 32002 37278
rect 35646 37266 35698 37278
rect 32386 37214 32398 37266
rect 32450 37214 32462 37266
rect 31950 37202 32002 37214
rect 35646 37202 35698 37214
rect 35870 37266 35922 37278
rect 35870 37202 35922 37214
rect 38110 37266 38162 37278
rect 38110 37202 38162 37214
rect 38334 37266 38386 37278
rect 38334 37202 38386 37214
rect 42478 37266 42530 37278
rect 42802 37214 42814 37266
rect 42866 37214 42878 37266
rect 42478 37202 42530 37214
rect 17726 37154 17778 37166
rect 24782 37154 24834 37166
rect 18834 37102 18846 37154
rect 18898 37102 18910 37154
rect 19618 37102 19630 37154
rect 19682 37102 19694 37154
rect 23762 37102 23774 37154
rect 23826 37102 23838 37154
rect 17726 37090 17778 37102
rect 24782 37090 24834 37102
rect 25678 37154 25730 37166
rect 30046 37154 30098 37166
rect 29138 37102 29150 37154
rect 29202 37102 29214 37154
rect 25678 37090 25730 37102
rect 30046 37090 30098 37102
rect 32846 37154 32898 37166
rect 32846 37090 32898 37102
rect 33966 37154 34018 37166
rect 33966 37090 34018 37102
rect 35758 37154 35810 37166
rect 35758 37090 35810 37102
rect 41806 37154 41858 37166
rect 41806 37090 41858 37102
rect 42366 37154 42418 37166
rect 42366 37090 42418 37102
rect 6862 37042 6914 37054
rect 6862 36978 6914 36990
rect 7646 37042 7698 37054
rect 26910 37042 26962 37054
rect 15698 36990 15710 37042
rect 15762 36990 15774 37042
rect 19058 36990 19070 37042
rect 19122 36990 19134 37042
rect 7646 36978 7698 36990
rect 26910 36978 26962 36990
rect 30830 37042 30882 37054
rect 31154 36990 31166 37042
rect 31218 36990 31230 37042
rect 30830 36978 30882 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 2270 36706 2322 36718
rect 2270 36642 2322 36654
rect 4062 36706 4114 36718
rect 4062 36642 4114 36654
rect 9886 36706 9938 36718
rect 9886 36642 9938 36654
rect 12574 36706 12626 36718
rect 28478 36706 28530 36718
rect 27682 36654 27694 36706
rect 27746 36654 27758 36706
rect 12574 36642 12626 36654
rect 28478 36642 28530 36654
rect 31278 36706 31330 36718
rect 31278 36642 31330 36654
rect 41470 36706 41522 36718
rect 41470 36642 41522 36654
rect 1822 36594 1874 36606
rect 1822 36530 1874 36542
rect 6078 36594 6130 36606
rect 6078 36530 6130 36542
rect 6974 36594 7026 36606
rect 9214 36594 9266 36606
rect 26238 36594 26290 36606
rect 31390 36594 31442 36606
rect 7970 36542 7982 36594
rect 8034 36542 8046 36594
rect 10882 36542 10894 36594
rect 10946 36542 10958 36594
rect 27346 36542 27358 36594
rect 27410 36542 27422 36594
rect 28802 36542 28814 36594
rect 28866 36542 28878 36594
rect 6974 36530 7026 36542
rect 9214 36530 9266 36542
rect 26238 36530 26290 36542
rect 31390 36530 31442 36542
rect 31950 36594 32002 36606
rect 40798 36594 40850 36606
rect 43150 36594 43202 36606
rect 34850 36542 34862 36594
rect 34914 36542 34926 36594
rect 38658 36542 38670 36594
rect 38722 36542 38734 36594
rect 42354 36542 42366 36594
rect 42418 36542 42430 36594
rect 31950 36530 32002 36542
rect 40798 36530 40850 36542
rect 43150 36530 43202 36542
rect 4510 36482 4562 36494
rect 4510 36418 4562 36430
rect 4734 36482 4786 36494
rect 4734 36418 4786 36430
rect 4958 36482 5010 36494
rect 12350 36482 12402 36494
rect 13806 36482 13858 36494
rect 21982 36482 22034 36494
rect 7410 36430 7422 36482
rect 7474 36430 7486 36482
rect 8082 36430 8094 36482
rect 8146 36430 8158 36482
rect 10546 36430 10558 36482
rect 10610 36430 10622 36482
rect 11666 36430 11678 36482
rect 11730 36430 11742 36482
rect 12898 36430 12910 36482
rect 12962 36430 12974 36482
rect 15586 36430 15598 36482
rect 15650 36430 15662 36482
rect 16258 36430 16270 36482
rect 16322 36430 16334 36482
rect 17154 36430 17166 36482
rect 17218 36430 17230 36482
rect 19842 36430 19854 36482
rect 19906 36430 19918 36482
rect 4958 36418 5010 36430
rect 12350 36418 12402 36430
rect 13806 36418 13858 36430
rect 21982 36418 22034 36430
rect 22542 36482 22594 36494
rect 22542 36418 22594 36430
rect 22878 36482 22930 36494
rect 33630 36482 33682 36494
rect 41358 36482 41410 36494
rect 26898 36430 26910 36482
rect 26962 36430 26974 36482
rect 29586 36430 29598 36482
rect 29650 36430 29662 36482
rect 30482 36430 30494 36482
rect 30546 36430 30558 36482
rect 34626 36430 34638 36482
rect 34690 36430 34702 36482
rect 35970 36430 35982 36482
rect 36034 36430 36046 36482
rect 40114 36430 40126 36482
rect 40178 36430 40190 36482
rect 42466 36430 42478 36482
rect 42530 36430 42542 36482
rect 22878 36418 22930 36430
rect 33630 36418 33682 36430
rect 41358 36418 41410 36430
rect 2382 36370 2434 36382
rect 2382 36306 2434 36318
rect 2942 36370 2994 36382
rect 2942 36306 2994 36318
rect 3278 36370 3330 36382
rect 9774 36370 9826 36382
rect 14030 36370 14082 36382
rect 8306 36318 8318 36370
rect 8370 36318 8382 36370
rect 10658 36318 10670 36370
rect 10722 36318 10734 36370
rect 3278 36306 3330 36318
rect 9774 36306 9826 36318
rect 14030 36306 14082 36318
rect 14254 36370 14306 36382
rect 14254 36306 14306 36318
rect 14478 36370 14530 36382
rect 19630 36370 19682 36382
rect 15474 36318 15486 36370
rect 15538 36318 15550 36370
rect 16146 36318 16158 36370
rect 16210 36318 16222 36370
rect 18498 36318 18510 36370
rect 18562 36318 18574 36370
rect 14478 36306 14530 36318
rect 19630 36306 19682 36318
rect 20526 36370 20578 36382
rect 20526 36306 20578 36318
rect 21646 36370 21698 36382
rect 21646 36306 21698 36318
rect 21758 36370 21810 36382
rect 21758 36306 21810 36318
rect 23326 36370 23378 36382
rect 23326 36306 23378 36318
rect 23662 36370 23714 36382
rect 23662 36306 23714 36318
rect 24222 36370 24274 36382
rect 24222 36306 24274 36318
rect 24558 36370 24610 36382
rect 24558 36306 24610 36318
rect 28702 36370 28754 36382
rect 33182 36370 33234 36382
rect 29698 36318 29710 36370
rect 29762 36318 29774 36370
rect 28702 36306 28754 36318
rect 33182 36306 33234 36318
rect 33742 36370 33794 36382
rect 33742 36306 33794 36318
rect 36766 36370 36818 36382
rect 39106 36318 39118 36370
rect 39170 36318 39182 36370
rect 36766 36306 36818 36318
rect 6414 36258 6466 36270
rect 6414 36194 6466 36206
rect 9886 36258 9938 36270
rect 9886 36194 9938 36206
rect 17726 36258 17778 36270
rect 17726 36194 17778 36206
rect 18174 36258 18226 36270
rect 18174 36194 18226 36206
rect 19070 36258 19122 36270
rect 19070 36194 19122 36206
rect 20638 36258 20690 36270
rect 20638 36194 20690 36206
rect 20862 36258 20914 36270
rect 20862 36194 20914 36206
rect 22654 36258 22706 36270
rect 22654 36194 22706 36206
rect 25006 36258 25058 36270
rect 25006 36194 25058 36206
rect 25454 36258 25506 36270
rect 33966 36258 34018 36270
rect 30594 36206 30606 36258
rect 30658 36206 30670 36258
rect 25454 36194 25506 36206
rect 33966 36194 34018 36206
rect 41470 36258 41522 36270
rect 41470 36194 41522 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 1822 35922 1874 35934
rect 1822 35858 1874 35870
rect 2270 35922 2322 35934
rect 2270 35858 2322 35870
rect 3950 35922 4002 35934
rect 3950 35858 4002 35870
rect 4734 35922 4786 35934
rect 14590 35922 14642 35934
rect 8194 35870 8206 35922
rect 8258 35870 8270 35922
rect 4734 35858 4786 35870
rect 14590 35858 14642 35870
rect 16606 35922 16658 35934
rect 16606 35858 16658 35870
rect 21646 35922 21698 35934
rect 21646 35858 21698 35870
rect 22430 35922 22482 35934
rect 22430 35858 22482 35870
rect 23214 35922 23266 35934
rect 23214 35858 23266 35870
rect 23774 35922 23826 35934
rect 23774 35858 23826 35870
rect 26014 35922 26066 35934
rect 26014 35858 26066 35870
rect 27246 35922 27298 35934
rect 27246 35858 27298 35870
rect 27358 35922 27410 35934
rect 27358 35858 27410 35870
rect 27918 35922 27970 35934
rect 27918 35858 27970 35870
rect 32958 35922 33010 35934
rect 35086 35922 35138 35934
rect 34178 35870 34190 35922
rect 34242 35870 34254 35922
rect 32958 35858 33010 35870
rect 35086 35858 35138 35870
rect 35758 35922 35810 35934
rect 35758 35858 35810 35870
rect 36094 35922 36146 35934
rect 36094 35858 36146 35870
rect 37214 35922 37266 35934
rect 37214 35858 37266 35870
rect 38446 35922 38498 35934
rect 38446 35858 38498 35870
rect 39006 35922 39058 35934
rect 39006 35858 39058 35870
rect 39118 35922 39170 35934
rect 39118 35858 39170 35870
rect 41694 35922 41746 35934
rect 41694 35858 41746 35870
rect 41806 35922 41858 35934
rect 41806 35858 41858 35870
rect 54350 35922 54402 35934
rect 54350 35858 54402 35870
rect 3614 35810 3666 35822
rect 3614 35746 3666 35758
rect 4174 35810 4226 35822
rect 8878 35810 8930 35822
rect 11902 35810 11954 35822
rect 21534 35810 21586 35822
rect 5282 35758 5294 35810
rect 5346 35758 5358 35810
rect 10994 35758 11006 35810
rect 11058 35758 11070 35810
rect 12786 35758 12798 35810
rect 12850 35758 12862 35810
rect 13234 35758 13246 35810
rect 13298 35758 13310 35810
rect 17714 35758 17726 35810
rect 17778 35758 17790 35810
rect 20626 35758 20638 35810
rect 20690 35758 20702 35810
rect 4174 35746 4226 35758
rect 8878 35746 8930 35758
rect 11902 35746 11954 35758
rect 21534 35746 21586 35758
rect 27470 35810 27522 35822
rect 27470 35746 27522 35758
rect 32734 35810 32786 35822
rect 32734 35746 32786 35758
rect 35870 35810 35922 35822
rect 35870 35746 35922 35758
rect 39230 35810 39282 35822
rect 39230 35746 39282 35758
rect 41582 35810 41634 35822
rect 41582 35746 41634 35758
rect 3838 35698 3890 35710
rect 3042 35646 3054 35698
rect 3106 35646 3118 35698
rect 3838 35634 3890 35646
rect 5630 35698 5682 35710
rect 6750 35698 6802 35710
rect 6290 35646 6302 35698
rect 6354 35646 6366 35698
rect 5630 35634 5682 35646
rect 6750 35634 6802 35646
rect 8654 35698 8706 35710
rect 8654 35634 8706 35646
rect 8766 35698 8818 35710
rect 14926 35698 14978 35710
rect 10322 35646 10334 35698
rect 10386 35646 10398 35698
rect 11442 35646 11454 35698
rect 11506 35646 11518 35698
rect 12450 35646 12462 35698
rect 12514 35646 12526 35698
rect 13458 35646 13470 35698
rect 13522 35646 13534 35698
rect 14018 35646 14030 35698
rect 14082 35646 14094 35698
rect 8766 35634 8818 35646
rect 14926 35634 14978 35646
rect 16942 35698 16994 35710
rect 19294 35698 19346 35710
rect 29486 35698 29538 35710
rect 18274 35646 18286 35698
rect 18338 35646 18350 35698
rect 18946 35646 18958 35698
rect 19010 35646 19022 35698
rect 19394 35646 19406 35698
rect 19458 35646 19470 35698
rect 20850 35646 20862 35698
rect 20914 35646 20926 35698
rect 21858 35646 21870 35698
rect 21922 35646 21934 35698
rect 22642 35646 22654 35698
rect 22706 35646 22718 35698
rect 23986 35646 23998 35698
rect 24050 35646 24062 35698
rect 29026 35646 29038 35698
rect 29090 35646 29102 35698
rect 16942 35634 16994 35646
rect 19294 35634 19346 35646
rect 29486 35634 29538 35646
rect 32622 35698 32674 35710
rect 32622 35634 32674 35646
rect 33630 35698 33682 35710
rect 33630 35634 33682 35646
rect 33854 35698 33906 35710
rect 33854 35634 33906 35646
rect 34862 35698 34914 35710
rect 34862 35634 34914 35646
rect 34974 35698 35026 35710
rect 34974 35634 35026 35646
rect 35422 35698 35474 35710
rect 36306 35646 36318 35698
rect 36370 35646 36382 35698
rect 54898 35646 54910 35698
rect 54962 35646 54974 35698
rect 35422 35634 35474 35646
rect 7198 35586 7250 35598
rect 7198 35522 7250 35534
rect 7646 35586 7698 35598
rect 7646 35522 7698 35534
rect 9774 35586 9826 35598
rect 15598 35586 15650 35598
rect 11330 35534 11342 35586
rect 11394 35534 11406 35586
rect 9774 35522 9826 35534
rect 15598 35522 15650 35534
rect 16046 35586 16098 35598
rect 16046 35522 16098 35534
rect 24670 35586 24722 35598
rect 24670 35522 24722 35534
rect 25566 35586 25618 35598
rect 25566 35522 25618 35534
rect 28590 35586 28642 35598
rect 28590 35522 28642 35534
rect 30046 35586 30098 35598
rect 30046 35522 30098 35534
rect 30718 35586 30770 35598
rect 56018 35534 56030 35586
rect 56082 35534 56094 35586
rect 30718 35522 30770 35534
rect 2718 35474 2770 35486
rect 2718 35410 2770 35422
rect 3054 35474 3106 35486
rect 24782 35474 24834 35486
rect 7186 35422 7198 35474
rect 7250 35471 7262 35474
rect 7858 35471 7870 35474
rect 7250 35425 7870 35471
rect 7250 35422 7262 35425
rect 7858 35422 7870 35425
rect 7922 35422 7934 35474
rect 19954 35422 19966 35474
rect 20018 35422 20030 35474
rect 3054 35410 3106 35422
rect 24782 35410 24834 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 9102 35138 9154 35150
rect 28590 35138 28642 35150
rect 11554 35086 11566 35138
rect 11618 35086 11630 35138
rect 9102 35074 9154 35086
rect 28590 35074 28642 35086
rect 37550 35138 37602 35150
rect 37550 35074 37602 35086
rect 5630 35026 5682 35038
rect 7310 35026 7362 35038
rect 6626 34974 6638 35026
rect 6690 34974 6702 35026
rect 5630 34962 5682 34974
rect 7310 34962 7362 34974
rect 9326 35026 9378 35038
rect 12574 35026 12626 35038
rect 11442 34974 11454 35026
rect 11506 34974 11518 35026
rect 9326 34962 9378 34974
rect 12574 34962 12626 34974
rect 15710 35026 15762 35038
rect 26350 35026 26402 35038
rect 27918 35026 27970 35038
rect 25218 34974 25230 35026
rect 25282 34974 25294 35026
rect 26898 34974 26910 35026
rect 26962 34974 26974 35026
rect 15710 34962 15762 34974
rect 26350 34962 26402 34974
rect 27918 34962 27970 34974
rect 32062 35026 32114 35038
rect 32062 34962 32114 34974
rect 34526 35026 34578 35038
rect 34526 34962 34578 34974
rect 35646 35026 35698 35038
rect 37762 34974 37774 35026
rect 37826 34974 37838 35026
rect 35646 34962 35698 34974
rect 2158 34914 2210 34926
rect 2158 34850 2210 34862
rect 3838 34914 3890 34926
rect 6190 34914 6242 34926
rect 11118 34914 11170 34926
rect 16942 34914 16994 34926
rect 20862 34914 20914 34926
rect 26574 34914 26626 34926
rect 4722 34862 4734 34914
rect 4786 34862 4798 34914
rect 10322 34862 10334 34914
rect 10386 34862 10398 34914
rect 12898 34862 12910 34914
rect 12962 34862 12974 34914
rect 14914 34862 14926 34914
rect 14978 34862 14990 34914
rect 17826 34862 17838 34914
rect 17890 34862 17902 34914
rect 18274 34862 18286 34914
rect 18338 34862 18350 34914
rect 19170 34862 19182 34914
rect 19234 34862 19246 34914
rect 24658 34862 24670 34914
rect 24722 34862 24734 34914
rect 25778 34862 25790 34914
rect 25842 34862 25854 34914
rect 3838 34850 3890 34862
rect 6190 34850 6242 34862
rect 11118 34850 11170 34862
rect 16942 34850 16994 34862
rect 20862 34850 20914 34862
rect 26574 34850 26626 34862
rect 28478 34914 28530 34926
rect 28478 34850 28530 34862
rect 29934 34914 29986 34926
rect 32510 34914 32562 34926
rect 31378 34862 31390 34914
rect 31442 34862 31454 34914
rect 31826 34862 31838 34914
rect 31890 34862 31902 34914
rect 29934 34850 29986 34862
rect 32510 34850 32562 34862
rect 39902 34914 39954 34926
rect 40450 34862 40462 34914
rect 40514 34862 40526 34914
rect 39902 34850 39954 34862
rect 7870 34802 7922 34814
rect 7870 34738 7922 34750
rect 8206 34802 8258 34814
rect 13694 34802 13746 34814
rect 8754 34750 8766 34802
rect 8818 34750 8830 34802
rect 10546 34750 10558 34802
rect 10610 34750 10622 34802
rect 8206 34738 8258 34750
rect 13694 34738 13746 34750
rect 14030 34802 14082 34814
rect 15822 34802 15874 34814
rect 15138 34750 15150 34802
rect 15202 34750 15214 34802
rect 14030 34738 14082 34750
rect 15822 34738 15874 34750
rect 16606 34802 16658 34814
rect 16606 34738 16658 34750
rect 16718 34802 16770 34814
rect 29598 34802 29650 34814
rect 17490 34750 17502 34802
rect 17554 34750 17566 34802
rect 18386 34750 18398 34802
rect 18450 34750 18462 34802
rect 20514 34750 20526 34802
rect 20578 34750 20590 34802
rect 23874 34750 23886 34802
rect 23938 34750 23950 34802
rect 24770 34750 24782 34802
rect 24834 34750 24846 34802
rect 16718 34738 16770 34750
rect 29598 34738 29650 34750
rect 2606 34690 2658 34702
rect 4958 34690 5010 34702
rect 21534 34690 21586 34702
rect 2930 34638 2942 34690
rect 2994 34638 3006 34690
rect 3490 34638 3502 34690
rect 3554 34638 3566 34690
rect 18498 34638 18510 34690
rect 18562 34638 18574 34690
rect 2606 34626 2658 34638
rect 4958 34626 5010 34638
rect 21534 34626 21586 34638
rect 30606 34690 30658 34702
rect 30606 34626 30658 34638
rect 33742 34690 33794 34702
rect 33742 34626 33794 34638
rect 36766 34690 36818 34702
rect 36766 34626 36818 34638
rect 37774 34690 37826 34702
rect 37774 34626 37826 34638
rect 39006 34690 39058 34702
rect 39006 34626 39058 34638
rect 39454 34690 39506 34702
rect 43598 34690 43650 34702
rect 43026 34638 43038 34690
rect 43090 34638 43102 34690
rect 39454 34626 39506 34638
rect 43598 34626 43650 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 4398 34354 4450 34366
rect 4398 34290 4450 34302
rect 4958 34354 5010 34366
rect 4958 34290 5010 34302
rect 5406 34354 5458 34366
rect 5406 34290 5458 34302
rect 5742 34354 5794 34366
rect 8430 34354 8482 34366
rect 6290 34302 6302 34354
rect 6354 34302 6366 34354
rect 5742 34290 5794 34302
rect 8430 34290 8482 34302
rect 9886 34354 9938 34366
rect 9886 34290 9938 34302
rect 10334 34354 10386 34366
rect 10334 34290 10386 34302
rect 10782 34354 10834 34366
rect 10782 34290 10834 34302
rect 11230 34354 11282 34366
rect 11230 34290 11282 34302
rect 11678 34354 11730 34366
rect 11678 34290 11730 34302
rect 12126 34354 12178 34366
rect 12126 34290 12178 34302
rect 12574 34354 12626 34366
rect 12574 34290 12626 34302
rect 14030 34354 14082 34366
rect 15710 34354 15762 34366
rect 16942 34354 16994 34366
rect 21086 34354 21138 34366
rect 22766 34354 22818 34366
rect 25566 34354 25618 34366
rect 14914 34302 14926 34354
rect 14978 34302 14990 34354
rect 16146 34302 16158 34354
rect 16210 34302 16222 34354
rect 19282 34302 19294 34354
rect 19346 34302 19358 34354
rect 21634 34302 21646 34354
rect 21698 34302 21710 34354
rect 24210 34302 24222 34354
rect 24274 34302 24286 34354
rect 14030 34290 14082 34302
rect 15710 34290 15762 34302
rect 16942 34290 16994 34302
rect 21086 34290 21138 34302
rect 22766 34290 22818 34302
rect 25566 34290 25618 34302
rect 28254 34354 28306 34366
rect 28254 34290 28306 34302
rect 29262 34354 29314 34366
rect 29262 34290 29314 34302
rect 29710 34354 29762 34366
rect 29710 34290 29762 34302
rect 31726 34354 31778 34366
rect 31726 34290 31778 34302
rect 32734 34354 32786 34366
rect 32734 34290 32786 34302
rect 17950 34242 18002 34254
rect 3938 34190 3950 34242
rect 4002 34190 4014 34242
rect 7634 34190 7646 34242
rect 7698 34190 7710 34242
rect 17950 34178 18002 34190
rect 18622 34242 18674 34254
rect 18622 34178 18674 34190
rect 18734 34242 18786 34254
rect 18734 34178 18786 34190
rect 18846 34242 18898 34254
rect 18846 34178 18898 34190
rect 23102 34242 23154 34254
rect 32622 34242 32674 34254
rect 23874 34190 23886 34242
rect 23938 34190 23950 34242
rect 24434 34190 24446 34242
rect 24498 34190 24510 34242
rect 34066 34190 34078 34242
rect 34130 34190 34142 34242
rect 37090 34190 37102 34242
rect 37154 34190 37166 34242
rect 23102 34178 23154 34190
rect 32622 34178 32674 34190
rect 6862 34130 6914 34142
rect 2818 34078 2830 34130
rect 2882 34078 2894 34130
rect 3714 34078 3726 34130
rect 3778 34078 3790 34130
rect 6862 34066 6914 34078
rect 7982 34130 8034 34142
rect 7982 34066 8034 34078
rect 13470 34130 13522 34142
rect 14590 34130 14642 34142
rect 13794 34078 13806 34130
rect 13858 34078 13870 34130
rect 13470 34066 13522 34078
rect 14590 34066 14642 34078
rect 16494 34130 16546 34142
rect 16494 34066 16546 34078
rect 19742 34130 19794 34142
rect 19742 34066 19794 34078
rect 20750 34130 20802 34142
rect 22430 34130 22482 34142
rect 21858 34078 21870 34130
rect 21922 34078 21934 34130
rect 20750 34066 20802 34078
rect 22430 34066 22482 34078
rect 22766 34130 22818 34142
rect 27806 34130 27858 34142
rect 24658 34078 24670 34130
rect 24722 34078 24734 34130
rect 22766 34066 22818 34078
rect 27806 34066 27858 34078
rect 29934 34130 29986 34142
rect 29934 34066 29986 34078
rect 30382 34130 30434 34142
rect 30382 34066 30434 34078
rect 32958 34130 33010 34142
rect 32958 34066 33010 34078
rect 8878 34018 8930 34030
rect 1922 33966 1934 34018
rect 1986 33966 1998 34018
rect 8878 33954 8930 33966
rect 13022 34018 13074 34030
rect 13022 33954 13074 33966
rect 20190 34018 20242 34030
rect 20190 33954 20242 33966
rect 26014 34018 26066 34030
rect 26014 33954 26066 33966
rect 28702 34018 28754 34030
rect 28702 33954 28754 33966
rect 29822 34018 29874 34030
rect 29822 33954 29874 33966
rect 31166 34018 31218 34030
rect 31166 33954 31218 33966
rect 31614 34018 31666 34030
rect 36306 33966 36318 34018
rect 36370 33966 36382 34018
rect 38210 33966 38222 34018
rect 38274 33966 38286 34018
rect 31614 33954 31666 33966
rect 6638 33906 6690 33918
rect 6638 33842 6690 33854
rect 14142 33906 14194 33918
rect 14142 33842 14194 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 3726 33570 3778 33582
rect 3726 33506 3778 33518
rect 6638 33570 6690 33582
rect 6638 33506 6690 33518
rect 9550 33570 9602 33582
rect 9550 33506 9602 33518
rect 9886 33570 9938 33582
rect 28926 33570 28978 33582
rect 11218 33518 11230 33570
rect 11282 33567 11294 33570
rect 11778 33567 11790 33570
rect 11282 33521 11790 33567
rect 11282 33518 11294 33521
rect 11778 33518 11790 33521
rect 11842 33518 11854 33570
rect 17266 33518 17278 33570
rect 17330 33518 17342 33570
rect 23874 33518 23886 33570
rect 23938 33567 23950 33570
rect 24658 33567 24670 33570
rect 23938 33521 24670 33567
rect 23938 33518 23950 33521
rect 24658 33518 24670 33521
rect 24722 33518 24734 33570
rect 9886 33506 9938 33518
rect 28926 33506 28978 33518
rect 31726 33570 31778 33582
rect 31726 33506 31778 33518
rect 36878 33570 36930 33582
rect 36878 33506 36930 33518
rect 1934 33458 1986 33470
rect 1934 33394 1986 33406
rect 2382 33458 2434 33470
rect 2382 33394 2434 33406
rect 4622 33458 4674 33470
rect 4622 33394 4674 33406
rect 5742 33458 5794 33470
rect 5742 33394 5794 33406
rect 8094 33458 8146 33470
rect 8094 33394 8146 33406
rect 10558 33458 10610 33470
rect 10558 33394 10610 33406
rect 11006 33458 11058 33470
rect 11006 33394 11058 33406
rect 11454 33458 11506 33470
rect 11454 33394 11506 33406
rect 11902 33458 11954 33470
rect 11902 33394 11954 33406
rect 14366 33458 14418 33470
rect 14366 33394 14418 33406
rect 18734 33458 18786 33470
rect 18734 33394 18786 33406
rect 20414 33458 20466 33470
rect 20414 33394 20466 33406
rect 22094 33458 22146 33470
rect 22094 33394 22146 33406
rect 44494 33458 44546 33470
rect 44494 33394 44546 33406
rect 12910 33346 12962 33358
rect 2930 33294 2942 33346
rect 2994 33294 3006 33346
rect 8866 33294 8878 33346
rect 8930 33294 8942 33346
rect 12910 33282 12962 33294
rect 14926 33346 14978 33358
rect 16718 33346 16770 33358
rect 15922 33294 15934 33346
rect 15986 33294 15998 33346
rect 14926 33282 14978 33294
rect 16718 33282 16770 33294
rect 16942 33346 16994 33358
rect 16942 33282 16994 33294
rect 23438 33346 23490 33358
rect 23438 33282 23490 33294
rect 23774 33346 23826 33358
rect 23774 33282 23826 33294
rect 25454 33346 25506 33358
rect 29710 33346 29762 33358
rect 25890 33294 25902 33346
rect 25954 33294 25966 33346
rect 25454 33282 25506 33294
rect 29710 33282 29762 33294
rect 30046 33346 30098 33358
rect 30046 33282 30098 33294
rect 30382 33346 30434 33358
rect 30382 33282 30434 33294
rect 31054 33346 31106 33358
rect 31054 33282 31106 33294
rect 32734 33346 32786 33358
rect 32734 33282 32786 33294
rect 33406 33346 33458 33358
rect 37662 33346 37714 33358
rect 41470 33346 41522 33358
rect 33842 33294 33854 33346
rect 33906 33294 33918 33346
rect 37986 33294 37998 33346
rect 38050 33294 38062 33346
rect 33406 33282 33458 33294
rect 37662 33282 37714 33294
rect 41470 33282 41522 33294
rect 3166 33234 3218 33246
rect 3166 33170 3218 33182
rect 3838 33234 3890 33246
rect 3838 33170 3890 33182
rect 5854 33234 5906 33246
rect 5854 33170 5906 33182
rect 6750 33234 6802 33246
rect 6750 33170 6802 33182
rect 7310 33234 7362 33246
rect 7310 33170 7362 33182
rect 7422 33234 7474 33246
rect 13694 33234 13746 33246
rect 8978 33182 8990 33234
rect 9042 33182 9054 33234
rect 7422 33170 7474 33182
rect 13694 33170 13746 33182
rect 13806 33234 13858 33246
rect 13806 33170 13858 33182
rect 16158 33234 16210 33246
rect 16158 33170 16210 33182
rect 17838 33234 17890 33246
rect 17838 33170 17890 33182
rect 18174 33234 18226 33246
rect 18174 33170 18226 33182
rect 21646 33234 21698 33246
rect 21646 33170 21698 33182
rect 22654 33234 22706 33246
rect 22654 33170 22706 33182
rect 22766 33234 22818 33246
rect 22766 33170 22818 33182
rect 31838 33234 31890 33246
rect 42354 33182 42366 33234
rect 42418 33182 42430 33234
rect 31838 33170 31890 33182
rect 7646 33122 7698 33134
rect 7646 33058 7698 33070
rect 12238 33122 12290 33134
rect 12238 33058 12290 33070
rect 14030 33122 14082 33134
rect 14030 33058 14082 33070
rect 15262 33122 15314 33134
rect 15262 33058 15314 33070
rect 19294 33122 19346 33134
rect 19294 33058 19346 33070
rect 20862 33122 20914 33134
rect 20862 33058 20914 33070
rect 22990 33122 23042 33134
rect 22990 33058 23042 33070
rect 23550 33122 23602 33134
rect 23550 33058 23602 33070
rect 24110 33122 24162 33134
rect 24110 33058 24162 33070
rect 24558 33122 24610 33134
rect 29822 33122 29874 33134
rect 28242 33070 28254 33122
rect 28306 33070 28318 33122
rect 24558 33058 24610 33070
rect 29822 33058 29874 33070
rect 30830 33122 30882 33134
rect 30830 33058 30882 33070
rect 30942 33122 30994 33134
rect 30942 33058 30994 33070
rect 31726 33122 31778 33134
rect 31726 33058 31778 33070
rect 32398 33122 32450 33134
rect 41134 33122 41186 33134
rect 36306 33070 36318 33122
rect 36370 33070 36382 33122
rect 40338 33070 40350 33122
rect 40402 33070 40414 33122
rect 32398 33058 32450 33070
rect 41134 33058 41186 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 1934 32786 1986 32798
rect 1934 32722 1986 32734
rect 6078 32786 6130 32798
rect 6078 32722 6130 32734
rect 6414 32786 6466 32798
rect 11006 32786 11058 32798
rect 7186 32734 7198 32786
rect 7250 32734 7262 32786
rect 6414 32722 6466 32734
rect 11006 32722 11058 32734
rect 11230 32786 11282 32798
rect 11230 32722 11282 32734
rect 11678 32786 11730 32798
rect 14142 32786 14194 32798
rect 13122 32734 13134 32786
rect 13186 32734 13198 32786
rect 11678 32722 11730 32734
rect 14142 32722 14194 32734
rect 15150 32786 15202 32798
rect 15150 32722 15202 32734
rect 17614 32786 17666 32798
rect 17614 32722 17666 32734
rect 18174 32786 18226 32798
rect 18174 32722 18226 32734
rect 22094 32786 22146 32798
rect 22094 32722 22146 32734
rect 24110 32786 24162 32798
rect 24110 32722 24162 32734
rect 26910 32786 26962 32798
rect 26910 32722 26962 32734
rect 29374 32786 29426 32798
rect 29374 32722 29426 32734
rect 32062 32786 32114 32798
rect 32062 32722 32114 32734
rect 37214 32786 37266 32798
rect 37214 32722 37266 32734
rect 37550 32786 37602 32798
rect 37550 32722 37602 32734
rect 46622 32786 46674 32798
rect 46622 32722 46674 32734
rect 3950 32674 4002 32686
rect 3950 32610 4002 32622
rect 4958 32674 5010 32686
rect 4958 32610 5010 32622
rect 14814 32674 14866 32686
rect 14814 32610 14866 32622
rect 25678 32674 25730 32686
rect 25678 32610 25730 32622
rect 26014 32674 26066 32686
rect 26014 32610 26066 32622
rect 27806 32674 27858 32686
rect 36430 32674 36482 32686
rect 30370 32622 30382 32674
rect 30434 32622 30446 32674
rect 27806 32610 27858 32622
rect 36430 32610 36482 32622
rect 37998 32674 38050 32686
rect 51662 32674 51714 32686
rect 40338 32622 40350 32674
rect 40402 32622 40414 32674
rect 37998 32610 38050 32622
rect 51662 32610 51714 32622
rect 52670 32674 52722 32686
rect 52670 32610 52722 32622
rect 3278 32562 3330 32574
rect 2706 32510 2718 32562
rect 2770 32510 2782 32562
rect 3278 32498 3330 32510
rect 4286 32562 4338 32574
rect 4286 32498 4338 32510
rect 5406 32562 5458 32574
rect 8430 32562 8482 32574
rect 7410 32510 7422 32562
rect 7474 32510 7486 32562
rect 5406 32498 5458 32510
rect 8430 32498 8482 32510
rect 8766 32562 8818 32574
rect 8766 32498 8818 32510
rect 8990 32562 9042 32574
rect 8990 32498 9042 32510
rect 9998 32562 10050 32574
rect 9998 32498 10050 32510
rect 10894 32562 10946 32574
rect 12798 32562 12850 32574
rect 11890 32510 11902 32562
rect 11954 32510 11966 32562
rect 10894 32498 10946 32510
rect 12798 32498 12850 32510
rect 13582 32562 13634 32574
rect 13582 32498 13634 32510
rect 14030 32562 14082 32574
rect 14030 32498 14082 32510
rect 14254 32562 14306 32574
rect 16942 32562 16994 32574
rect 19518 32562 19570 32574
rect 28478 32562 28530 32574
rect 16258 32510 16270 32562
rect 16322 32510 16334 32562
rect 18946 32510 18958 32562
rect 19010 32510 19022 32562
rect 22866 32510 22878 32562
rect 22930 32510 22942 32562
rect 27122 32510 27134 32562
rect 27186 32510 27198 32562
rect 14254 32498 14306 32510
rect 16942 32498 16994 32510
rect 19518 32498 19570 32510
rect 28478 32498 28530 32510
rect 33518 32562 33570 32574
rect 48078 32562 48130 32574
rect 34178 32510 34190 32562
rect 34242 32510 34254 32562
rect 47506 32510 47518 32562
rect 47570 32510 47582 32562
rect 33518 32498 33570 32510
rect 48078 32498 48130 32510
rect 51998 32562 52050 32574
rect 51998 32498 52050 32510
rect 3390 32450 3442 32462
rect 3390 32386 3442 32398
rect 8542 32450 8594 32462
rect 8542 32386 8594 32398
rect 12574 32450 12626 32462
rect 19630 32450 19682 32462
rect 23550 32450 23602 32462
rect 16594 32398 16606 32450
rect 16658 32398 16670 32450
rect 23090 32398 23102 32450
rect 23154 32398 23166 32450
rect 12574 32386 12626 32398
rect 19630 32386 19682 32398
rect 23550 32386 23602 32398
rect 28926 32450 28978 32462
rect 28926 32386 28978 32398
rect 38670 32450 38722 32462
rect 41470 32450 41522 32462
rect 39106 32398 39118 32450
rect 39170 32398 39182 32450
rect 38670 32386 38722 32398
rect 41470 32386 41522 32398
rect 46174 32450 46226 32462
rect 46174 32386 46226 32398
rect 48190 32450 48242 32462
rect 48190 32386 48242 32398
rect 51102 32450 51154 32462
rect 51102 32386 51154 32398
rect 53230 32450 53282 32462
rect 53230 32386 53282 32398
rect 53678 32450 53730 32462
rect 53678 32386 53730 32398
rect 55022 32450 55074 32462
rect 55022 32386 55074 32398
rect 55918 32450 55970 32462
rect 55918 32386 55970 32398
rect 56366 32450 56418 32462
rect 56366 32386 56418 32398
rect 56814 32450 56866 32462
rect 56814 32386 56866 32398
rect 57374 32450 57426 32462
rect 57374 32386 57426 32398
rect 5182 32338 5234 32350
rect 5182 32274 5234 32286
rect 5630 32338 5682 32350
rect 5630 32274 5682 32286
rect 9886 32338 9938 32350
rect 9886 32274 9938 32286
rect 10222 32338 10274 32350
rect 10222 32274 10274 32286
rect 10334 32338 10386 32350
rect 10334 32274 10386 32286
rect 52558 32338 52610 32350
rect 52558 32274 52610 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 11118 32002 11170 32014
rect 11118 31938 11170 31950
rect 19518 32002 19570 32014
rect 19518 31938 19570 31950
rect 23326 32002 23378 32014
rect 23326 31938 23378 31950
rect 7758 31890 7810 31902
rect 7758 31826 7810 31838
rect 14590 31890 14642 31902
rect 14590 31826 14642 31838
rect 14926 31890 14978 31902
rect 14926 31826 14978 31838
rect 15710 31890 15762 31902
rect 15710 31826 15762 31838
rect 16158 31890 16210 31902
rect 16158 31826 16210 31838
rect 17054 31890 17106 31902
rect 17054 31826 17106 31838
rect 20302 31890 20354 31902
rect 20302 31826 20354 31838
rect 21982 31890 22034 31902
rect 29486 31890 29538 31902
rect 22418 31838 22430 31890
rect 22482 31838 22494 31890
rect 27346 31838 27358 31890
rect 27410 31838 27422 31890
rect 21982 31826 22034 31838
rect 29486 31826 29538 31838
rect 31390 31890 31442 31902
rect 53902 31890 53954 31902
rect 39442 31838 39454 31890
rect 39506 31838 39518 31890
rect 45714 31838 45726 31890
rect 45778 31838 45790 31890
rect 31390 31826 31442 31838
rect 53902 31826 53954 31838
rect 56926 31890 56978 31902
rect 56926 31826 56978 31838
rect 57262 31890 57314 31902
rect 57262 31826 57314 31838
rect 10110 31778 10162 31790
rect 2818 31726 2830 31778
rect 2882 31726 2894 31778
rect 4722 31726 4734 31778
rect 4786 31726 4798 31778
rect 5954 31726 5966 31778
rect 6018 31726 6030 31778
rect 6850 31726 6862 31778
rect 6914 31726 6926 31778
rect 10110 31714 10162 31726
rect 10782 31778 10834 31790
rect 12462 31778 12514 31790
rect 33854 31778 33906 31790
rect 11890 31726 11902 31778
rect 11954 31726 11966 31778
rect 19842 31726 19854 31778
rect 19906 31726 19918 31778
rect 23650 31726 23662 31778
rect 23714 31726 23726 31778
rect 10782 31714 10834 31726
rect 12462 31714 12514 31726
rect 33854 31714 33906 31726
rect 34190 31778 34242 31790
rect 34190 31714 34242 31726
rect 36766 31778 36818 31790
rect 36766 31714 36818 31726
rect 40126 31778 40178 31790
rect 47630 31778 47682 31790
rect 40450 31726 40462 31778
rect 40514 31726 40526 31778
rect 46050 31726 46062 31778
rect 46114 31726 46126 31778
rect 40126 31714 40178 31726
rect 47630 31714 47682 31726
rect 48190 31778 48242 31790
rect 48190 31714 48242 31726
rect 51550 31778 51602 31790
rect 51550 31714 51602 31726
rect 52446 31778 52498 31790
rect 55358 31778 55410 31790
rect 54674 31726 54686 31778
rect 54738 31726 54750 31778
rect 52446 31714 52498 31726
rect 55358 31714 55410 31726
rect 1822 31666 1874 31678
rect 1822 31602 1874 31614
rect 2158 31666 2210 31678
rect 2158 31602 2210 31614
rect 3054 31666 3106 31678
rect 3054 31602 3106 31614
rect 3614 31666 3666 31678
rect 3614 31602 3666 31614
rect 3950 31666 4002 31678
rect 3950 31602 4002 31614
rect 4958 31666 5010 31678
rect 4958 31602 5010 31614
rect 8430 31666 8482 31678
rect 8430 31602 8482 31614
rect 8766 31666 8818 31678
rect 8766 31602 8818 31614
rect 9550 31666 9602 31678
rect 9550 31602 9602 31614
rect 9998 31666 10050 31678
rect 9998 31602 10050 31614
rect 10558 31666 10610 31678
rect 14142 31666 14194 31678
rect 11666 31614 11678 31666
rect 11730 31614 11742 31666
rect 10558 31602 10610 31614
rect 14142 31602 14194 31614
rect 22542 31666 22594 31678
rect 22542 31602 22594 31614
rect 22766 31666 22818 31678
rect 33966 31666 34018 31678
rect 46510 31666 46562 31678
rect 28578 31614 28590 31666
rect 28642 31614 28654 31666
rect 36418 31614 36430 31666
rect 36482 31614 36494 31666
rect 38434 31614 38446 31666
rect 38498 31614 38510 31666
rect 22766 31602 22818 31614
rect 33966 31602 34018 31614
rect 46510 31602 46562 31614
rect 6638 31554 6690 31566
rect 5730 31502 5742 31554
rect 5794 31502 5806 31554
rect 6638 31490 6690 31502
rect 9774 31554 9826 31566
rect 9774 31490 9826 31502
rect 13022 31554 13074 31566
rect 13022 31490 13074 31502
rect 13582 31554 13634 31566
rect 13582 31490 13634 31502
rect 19630 31554 19682 31566
rect 19630 31490 19682 31502
rect 23438 31554 23490 31566
rect 23438 31490 23490 31502
rect 24110 31554 24162 31566
rect 24110 31490 24162 31502
rect 26574 31554 26626 31566
rect 43598 31554 43650 31566
rect 43026 31502 43038 31554
rect 43090 31502 43102 31554
rect 26574 31490 26626 31502
rect 43598 31490 43650 31502
rect 47294 31554 47346 31566
rect 47294 31490 47346 31502
rect 47518 31554 47570 31566
rect 47518 31490 47570 31502
rect 48526 31554 48578 31566
rect 48526 31490 48578 31502
rect 49086 31554 49138 31566
rect 49086 31490 49138 31502
rect 50206 31554 50258 31566
rect 50206 31490 50258 31502
rect 50766 31554 50818 31566
rect 50766 31490 50818 31502
rect 51214 31554 51266 31566
rect 53342 31554 53394 31566
rect 52098 31502 52110 31554
rect 52162 31502 52174 31554
rect 51214 31490 51266 31502
rect 53342 31490 53394 31502
rect 54462 31554 54514 31566
rect 54462 31490 54514 31502
rect 55694 31554 55746 31566
rect 55694 31490 55746 31502
rect 56254 31554 56306 31566
rect 56254 31490 56306 31502
rect 57710 31554 57762 31566
rect 57710 31490 57762 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 2046 31218 2098 31230
rect 2046 31154 2098 31166
rect 3166 31218 3218 31230
rect 3166 31154 3218 31166
rect 3614 31218 3666 31230
rect 3614 31154 3666 31166
rect 4734 31218 4786 31230
rect 7310 31218 7362 31230
rect 6402 31166 6414 31218
rect 6466 31166 6478 31218
rect 4734 31154 4786 31166
rect 7310 31154 7362 31166
rect 8094 31218 8146 31230
rect 8094 31154 8146 31166
rect 8542 31218 8594 31230
rect 8542 31154 8594 31166
rect 9998 31218 10050 31230
rect 14142 31218 14194 31230
rect 11442 31166 11454 31218
rect 11506 31166 11518 31218
rect 9998 31154 10050 31166
rect 14142 31154 14194 31166
rect 14590 31218 14642 31230
rect 14590 31154 14642 31166
rect 15486 31218 15538 31230
rect 15486 31154 15538 31166
rect 17614 31218 17666 31230
rect 17614 31154 17666 31166
rect 22654 31218 22706 31230
rect 22654 31154 22706 31166
rect 22766 31218 22818 31230
rect 22766 31154 22818 31166
rect 23774 31218 23826 31230
rect 23774 31154 23826 31166
rect 27134 31218 27186 31230
rect 27134 31154 27186 31166
rect 31278 31218 31330 31230
rect 45838 31218 45890 31230
rect 40338 31166 40350 31218
rect 40402 31166 40414 31218
rect 31278 31154 31330 31166
rect 45838 31154 45890 31166
rect 47854 31218 47906 31230
rect 47854 31154 47906 31166
rect 48638 31218 48690 31230
rect 48638 31154 48690 31166
rect 50654 31218 50706 31230
rect 50654 31154 50706 31166
rect 15262 31106 15314 31118
rect 13346 31054 13358 31106
rect 13410 31054 13422 31106
rect 15262 31042 15314 31054
rect 30494 31106 30546 31118
rect 30494 31042 30546 31054
rect 32062 31106 32114 31118
rect 32062 31042 32114 31054
rect 36206 31106 36258 31118
rect 44270 31106 44322 31118
rect 49534 31106 49586 31118
rect 42914 31054 42926 31106
rect 42978 31054 42990 31106
rect 48178 31054 48190 31106
rect 48242 31054 48254 31106
rect 36206 31042 36258 31054
rect 44270 31042 44322 31054
rect 49534 31042 49586 31054
rect 51326 31106 51378 31118
rect 51326 31042 51378 31054
rect 51662 31106 51714 31118
rect 51662 31042 51714 31054
rect 54910 31106 54962 31118
rect 54910 31042 54962 31054
rect 5070 30994 5122 31006
rect 5070 30930 5122 30942
rect 6750 30994 6802 31006
rect 6750 30930 6802 30942
rect 7646 30994 7698 31006
rect 7646 30930 7698 30942
rect 9102 30994 9154 31006
rect 9102 30930 9154 30942
rect 10334 30994 10386 31006
rect 10334 30930 10386 30942
rect 15038 30994 15090 31006
rect 27582 30994 27634 31006
rect 37438 30994 37490 31006
rect 45726 30994 45778 31006
rect 18386 30942 18398 30994
rect 18450 30942 18462 30994
rect 18834 30942 18846 30994
rect 18898 30942 18910 30994
rect 21074 30942 21086 30994
rect 21138 30942 21150 30994
rect 28130 30942 28142 30994
rect 28194 30942 28206 30994
rect 37762 30942 37774 30994
rect 37826 30942 37838 30994
rect 44034 30942 44046 30994
rect 44098 30942 44110 30994
rect 45378 30942 45390 30994
rect 45442 30942 45454 30994
rect 15038 30930 15090 30942
rect 27582 30930 27634 30942
rect 37438 30930 37490 30942
rect 45726 30930 45778 30942
rect 45950 30994 46002 31006
rect 45950 30930 46002 30942
rect 46510 30994 46562 31006
rect 46510 30930 46562 30942
rect 49870 30994 49922 31006
rect 55246 30994 55298 31006
rect 50418 30942 50430 30994
rect 50482 30942 50494 30994
rect 53106 30942 53118 30994
rect 53170 30942 53182 30994
rect 49870 30930 49922 30942
rect 55246 30930 55298 30942
rect 2382 30882 2434 30894
rect 2382 30818 2434 30830
rect 4174 30882 4226 30894
rect 4174 30818 4226 30830
rect 5518 30882 5570 30894
rect 5518 30818 5570 30830
rect 10894 30882 10946 30894
rect 10894 30818 10946 30830
rect 11118 30882 11170 30894
rect 15150 30882 15202 30894
rect 12002 30830 12014 30882
rect 12066 30830 12078 30882
rect 11118 30818 11170 30830
rect 15150 30818 15202 30830
rect 16046 30882 16098 30894
rect 16046 30818 16098 30830
rect 23438 30882 23490 30894
rect 23438 30818 23490 30830
rect 24334 30882 24386 30894
rect 24334 30818 24386 30830
rect 31614 30882 31666 30894
rect 31614 30818 31666 30830
rect 32622 30882 32674 30894
rect 32622 30818 32674 30830
rect 35422 30882 35474 30894
rect 35422 30818 35474 30830
rect 35870 30882 35922 30894
rect 44718 30882 44770 30894
rect 41570 30830 41582 30882
rect 41634 30830 41646 30882
rect 35870 30818 35922 30830
rect 44718 30818 44770 30830
rect 46846 30882 46898 30894
rect 46846 30818 46898 30830
rect 47294 30882 47346 30894
rect 53790 30882 53842 30894
rect 52658 30830 52670 30882
rect 52722 30830 52734 30882
rect 47294 30818 47346 30830
rect 53790 30818 53842 30830
rect 54350 30882 54402 30894
rect 54350 30818 54402 30830
rect 55694 30882 55746 30894
rect 55694 30818 55746 30830
rect 56142 30882 56194 30894
rect 56142 30818 56194 30830
rect 56702 30882 56754 30894
rect 56702 30818 56754 30830
rect 57486 30882 57538 30894
rect 57486 30818 57538 30830
rect 57822 30882 57874 30894
rect 57822 30818 57874 30830
rect 22878 30770 22930 30782
rect 40910 30770 40962 30782
rect 3602 30718 3614 30770
rect 3666 30767 3678 30770
rect 4162 30767 4174 30770
rect 3666 30721 4174 30767
rect 3666 30718 3678 30721
rect 4162 30718 4174 30721
rect 4226 30718 4238 30770
rect 21970 30718 21982 30770
rect 22034 30718 22046 30770
rect 23202 30718 23214 30770
rect 23266 30767 23278 30770
rect 23426 30767 23438 30770
rect 23266 30721 23438 30767
rect 23266 30718 23278 30721
rect 23426 30718 23438 30721
rect 23490 30718 23502 30770
rect 35410 30718 35422 30770
rect 35474 30767 35486 30770
rect 36082 30767 36094 30770
rect 35474 30721 36094 30767
rect 35474 30718 35486 30721
rect 36082 30718 36094 30721
rect 36146 30718 36158 30770
rect 22878 30706 22930 30718
rect 40910 30706 40962 30718
rect 50766 30770 50818 30782
rect 52322 30718 52334 30770
rect 52386 30718 52398 30770
rect 53890 30718 53902 30770
rect 53954 30767 53966 30770
rect 54674 30767 54686 30770
rect 53954 30721 54686 30767
rect 53954 30718 53966 30721
rect 54674 30718 54686 30721
rect 54738 30718 54750 30770
rect 55794 30718 55806 30770
rect 55858 30767 55870 30770
rect 56130 30767 56142 30770
rect 55858 30721 56142 30767
rect 55858 30718 55870 30721
rect 56130 30718 56142 30721
rect 56194 30718 56206 30770
rect 50766 30706 50818 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 14702 30434 14754 30446
rect 3714 30382 3726 30434
rect 3778 30431 3790 30434
rect 3938 30431 3950 30434
rect 3778 30385 3950 30431
rect 3778 30382 3790 30385
rect 3938 30382 3950 30385
rect 4002 30382 4014 30434
rect 14702 30370 14754 30382
rect 19182 30434 19234 30446
rect 33182 30434 33234 30446
rect 22866 30382 22878 30434
rect 22930 30431 22942 30434
rect 23202 30431 23214 30434
rect 22930 30385 23214 30431
rect 22930 30382 22942 30385
rect 23202 30382 23214 30385
rect 23266 30382 23278 30434
rect 19182 30370 19234 30382
rect 33182 30370 33234 30382
rect 34078 30434 34130 30446
rect 34078 30370 34130 30382
rect 38110 30434 38162 30446
rect 38110 30370 38162 30382
rect 3726 30322 3778 30334
rect 3726 30258 3778 30270
rect 19742 30322 19794 30334
rect 19742 30258 19794 30270
rect 21982 30322 22034 30334
rect 21982 30258 22034 30270
rect 33742 30322 33794 30334
rect 33742 30258 33794 30270
rect 36430 30322 36482 30334
rect 36430 30258 36482 30270
rect 36654 30322 36706 30334
rect 36654 30258 36706 30270
rect 43262 30322 43314 30334
rect 43262 30258 43314 30270
rect 50654 30322 50706 30334
rect 50654 30258 50706 30270
rect 1934 30210 1986 30222
rect 1934 30146 1986 30158
rect 5742 30210 5794 30222
rect 7982 30210 8034 30222
rect 7298 30158 7310 30210
rect 7362 30158 7374 30210
rect 5742 30146 5794 30158
rect 7982 30146 8034 30158
rect 11902 30210 11954 30222
rect 11902 30146 11954 30158
rect 14926 30210 14978 30222
rect 14926 30146 14978 30158
rect 15598 30210 15650 30222
rect 15598 30146 15650 30158
rect 15710 30210 15762 30222
rect 18958 30210 19010 30222
rect 16258 30158 16270 30210
rect 16322 30158 16334 30210
rect 16930 30158 16942 30210
rect 16994 30158 17006 30210
rect 17938 30158 17950 30210
rect 18002 30158 18014 30210
rect 15710 30146 15762 30158
rect 18958 30146 19010 30158
rect 19630 30210 19682 30222
rect 19630 30146 19682 30158
rect 20190 30210 20242 30222
rect 20190 30146 20242 30158
rect 20526 30210 20578 30222
rect 20526 30146 20578 30158
rect 23326 30210 23378 30222
rect 27022 30210 27074 30222
rect 23874 30158 23886 30210
rect 23938 30158 23950 30210
rect 23326 30146 23378 30158
rect 27022 30146 27074 30158
rect 30270 30210 30322 30222
rect 30270 30146 30322 30158
rect 31950 30210 32002 30222
rect 31950 30146 32002 30158
rect 41134 30210 41186 30222
rect 41134 30146 41186 30158
rect 43934 30210 43986 30222
rect 43934 30146 43986 30158
rect 44494 30210 44546 30222
rect 44494 30146 44546 30158
rect 46062 30210 46114 30222
rect 46062 30146 46114 30158
rect 50878 30210 50930 30222
rect 50878 30146 50930 30158
rect 52558 30210 52610 30222
rect 52558 30146 52610 30158
rect 53790 30210 53842 30222
rect 53790 30146 53842 30158
rect 57038 30210 57090 30222
rect 57038 30146 57090 30158
rect 2382 30098 2434 30110
rect 2382 30034 2434 30046
rect 2718 30098 2770 30110
rect 2718 30034 2770 30046
rect 6414 30098 6466 30110
rect 6414 30034 6466 30046
rect 8206 30098 8258 30110
rect 8206 30034 8258 30046
rect 8766 30098 8818 30110
rect 8766 30034 8818 30046
rect 9102 30098 9154 30110
rect 9102 30034 9154 30046
rect 10222 30098 10274 30110
rect 10222 30034 10274 30046
rect 10558 30098 10610 30110
rect 12910 30098 12962 30110
rect 19406 30098 19458 30110
rect 11442 30046 11454 30098
rect 11506 30046 11518 30098
rect 17154 30046 17166 30098
rect 17218 30046 17230 30098
rect 17714 30046 17726 30098
rect 17778 30046 17790 30098
rect 10558 30034 10610 30046
rect 12910 30034 12962 30046
rect 19406 30034 19458 30046
rect 20414 30098 20466 30110
rect 20414 30034 20466 30046
rect 29598 30098 29650 30110
rect 29598 30034 29650 30046
rect 29710 30098 29762 30110
rect 29710 30034 29762 30046
rect 32286 30098 32338 30110
rect 32286 30034 32338 30046
rect 32846 30098 32898 30110
rect 32846 30034 32898 30046
rect 35086 30098 35138 30110
rect 35086 30034 35138 30046
rect 35422 30098 35474 30110
rect 35422 30034 35474 30046
rect 35870 30098 35922 30110
rect 35870 30034 35922 30046
rect 36094 30098 36146 30110
rect 41694 30098 41746 30110
rect 40226 30046 40238 30098
rect 40290 30046 40302 30098
rect 36094 30034 36146 30046
rect 41694 30034 41746 30046
rect 42478 30098 42530 30110
rect 42478 30034 42530 30046
rect 44158 30098 44210 30110
rect 44158 30034 44210 30046
rect 46510 30098 46562 30110
rect 46510 30034 46562 30046
rect 46734 30098 46786 30110
rect 46734 30034 46786 30046
rect 48526 30098 48578 30110
rect 48526 30034 48578 30046
rect 49310 30098 49362 30110
rect 49310 30034 49362 30046
rect 49646 30098 49698 30110
rect 49646 30034 49698 30046
rect 50206 30098 50258 30110
rect 50206 30034 50258 30046
rect 50430 30098 50482 30110
rect 50430 30034 50482 30046
rect 55582 30098 55634 30110
rect 55582 30034 55634 30046
rect 56478 30098 56530 30110
rect 56478 30034 56530 30046
rect 3278 29986 3330 29998
rect 3278 29922 3330 29934
rect 4286 29986 4338 29998
rect 4286 29922 4338 29934
rect 4622 29986 4674 29998
rect 4622 29922 4674 29934
rect 9662 29986 9714 29998
rect 9662 29922 9714 29934
rect 11118 29986 11170 29998
rect 11118 29922 11170 29934
rect 12350 29986 12402 29998
rect 12350 29922 12402 29934
rect 13694 29986 13746 29998
rect 21534 29986 21586 29998
rect 14354 29934 14366 29986
rect 14418 29934 14430 29986
rect 13694 29922 13746 29934
rect 21534 29922 21586 29934
rect 22430 29986 22482 29998
rect 22430 29922 22482 29934
rect 22878 29986 22930 29998
rect 27358 29986 27410 29998
rect 26226 29934 26238 29986
rect 26290 29934 26302 29986
rect 22878 29922 22930 29934
rect 27358 29922 27410 29934
rect 29934 29986 29986 29998
rect 29934 29922 29986 29934
rect 30830 29986 30882 29998
rect 30830 29922 30882 29934
rect 31278 29986 31330 29998
rect 31278 29922 31330 29934
rect 32174 29986 32226 29998
rect 32174 29922 32226 29934
rect 33070 29986 33122 29998
rect 33070 29922 33122 29934
rect 33966 29986 34018 29998
rect 33966 29922 34018 29934
rect 34526 29986 34578 29998
rect 34526 29922 34578 29934
rect 35198 29986 35250 29998
rect 35198 29922 35250 29934
rect 36766 29986 36818 29998
rect 36766 29922 36818 29934
rect 37438 29986 37490 29998
rect 44270 29986 44322 29998
rect 42018 29934 42030 29986
rect 42082 29934 42094 29986
rect 37438 29922 37490 29934
rect 44270 29922 44322 29934
rect 45390 29986 45442 29998
rect 45390 29922 45442 29934
rect 46286 29986 46338 29998
rect 47630 29986 47682 29998
rect 47282 29934 47294 29986
rect 47346 29934 47358 29986
rect 46286 29922 46338 29934
rect 47630 29922 47682 29934
rect 48190 29986 48242 29998
rect 48190 29922 48242 29934
rect 51326 29986 51378 29998
rect 52222 29986 52274 29998
rect 51650 29934 51662 29986
rect 51714 29934 51726 29986
rect 51326 29922 51378 29934
rect 52222 29922 52274 29934
rect 53454 29986 53506 29998
rect 54910 29986 54962 29998
rect 54562 29934 54574 29986
rect 54626 29934 54638 29986
rect 53454 29922 53506 29934
rect 54910 29922 54962 29934
rect 55470 29986 55522 29998
rect 55470 29922 55522 29934
rect 56142 29986 56194 29998
rect 56142 29922 56194 29934
rect 57374 29986 57426 29998
rect 57374 29922 57426 29934
rect 57822 29986 57874 29998
rect 57822 29922 57874 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 2830 29650 2882 29662
rect 2830 29586 2882 29598
rect 3278 29650 3330 29662
rect 3278 29586 3330 29598
rect 4734 29650 4786 29662
rect 4734 29586 4786 29598
rect 6078 29650 6130 29662
rect 6078 29586 6130 29598
rect 6638 29650 6690 29662
rect 6638 29586 6690 29598
rect 7198 29650 7250 29662
rect 7198 29586 7250 29598
rect 7646 29650 7698 29662
rect 7646 29586 7698 29598
rect 8318 29650 8370 29662
rect 8318 29586 8370 29598
rect 8654 29650 8706 29662
rect 8654 29586 8706 29598
rect 16942 29650 16994 29662
rect 16942 29586 16994 29598
rect 18286 29650 18338 29662
rect 22318 29650 22370 29662
rect 21522 29598 21534 29650
rect 21586 29598 21598 29650
rect 18286 29586 18338 29598
rect 22318 29586 22370 29598
rect 22654 29650 22706 29662
rect 29262 29650 29314 29662
rect 28466 29598 28478 29650
rect 28530 29598 28542 29650
rect 22654 29586 22706 29598
rect 29262 29586 29314 29598
rect 30046 29650 30098 29662
rect 30046 29586 30098 29598
rect 30718 29650 30770 29662
rect 30718 29586 30770 29598
rect 35310 29650 35362 29662
rect 35310 29586 35362 29598
rect 37662 29650 37714 29662
rect 37662 29586 37714 29598
rect 41918 29650 41970 29662
rect 41918 29586 41970 29598
rect 42366 29650 42418 29662
rect 42366 29586 42418 29598
rect 43262 29650 43314 29662
rect 43262 29586 43314 29598
rect 43710 29650 43762 29662
rect 43710 29586 43762 29598
rect 44382 29650 44434 29662
rect 44382 29586 44434 29598
rect 44606 29650 44658 29662
rect 49646 29650 49698 29662
rect 47394 29598 47406 29650
rect 47458 29598 47470 29650
rect 44606 29586 44658 29598
rect 49646 29586 49698 29598
rect 54238 29650 54290 29662
rect 54238 29586 54290 29598
rect 56702 29650 56754 29662
rect 56702 29586 56754 29598
rect 4286 29538 4338 29550
rect 4286 29474 4338 29486
rect 5182 29538 5234 29550
rect 5182 29474 5234 29486
rect 9662 29538 9714 29550
rect 9662 29474 9714 29486
rect 15374 29538 15426 29550
rect 15374 29474 15426 29486
rect 23550 29538 23602 29550
rect 23550 29474 23602 29486
rect 32510 29538 32562 29550
rect 32510 29474 32562 29486
rect 35534 29538 35586 29550
rect 35534 29474 35586 29486
rect 36542 29538 36594 29550
rect 36542 29474 36594 29486
rect 38334 29538 38386 29550
rect 38334 29474 38386 29486
rect 38670 29538 38722 29550
rect 38670 29474 38722 29486
rect 39118 29538 39170 29550
rect 44830 29538 44882 29550
rect 51214 29538 51266 29550
rect 41570 29486 41582 29538
rect 41634 29486 41646 29538
rect 42914 29486 42926 29538
rect 42978 29486 42990 29538
rect 45938 29486 45950 29538
rect 46002 29486 46014 29538
rect 50306 29486 50318 29538
rect 50370 29486 50382 29538
rect 39118 29474 39170 29486
rect 44830 29474 44882 29486
rect 51214 29474 51266 29486
rect 54350 29538 54402 29550
rect 54350 29474 54402 29486
rect 57486 29538 57538 29550
rect 57486 29474 57538 29486
rect 57822 29538 57874 29550
rect 57822 29474 57874 29486
rect 10446 29426 10498 29438
rect 14702 29426 14754 29438
rect 11442 29374 11454 29426
rect 11506 29374 11518 29426
rect 14242 29374 14254 29426
rect 14306 29374 14318 29426
rect 10446 29362 10498 29374
rect 14702 29362 14754 29374
rect 14814 29426 14866 29438
rect 18622 29426 18674 29438
rect 25566 29426 25618 29438
rect 33518 29426 33570 29438
rect 15586 29374 15598 29426
rect 15650 29374 15662 29426
rect 19282 29374 19294 29426
rect 19346 29374 19358 29426
rect 23314 29374 23326 29426
rect 23378 29374 23390 29426
rect 26114 29374 26126 29426
rect 26178 29374 26190 29426
rect 31826 29374 31838 29426
rect 31890 29374 31902 29426
rect 14814 29362 14866 29374
rect 18622 29362 18674 29374
rect 25566 29362 25618 29374
rect 33518 29362 33570 29374
rect 34862 29426 34914 29438
rect 34862 29362 34914 29374
rect 35086 29426 35138 29438
rect 35086 29362 35138 29374
rect 36430 29426 36482 29438
rect 36430 29362 36482 29374
rect 36766 29426 36818 29438
rect 36766 29362 36818 29374
rect 37102 29426 37154 29438
rect 37102 29362 37154 29374
rect 37550 29426 37602 29438
rect 37550 29362 37602 29374
rect 37774 29426 37826 29438
rect 47742 29426 47794 29438
rect 46050 29374 46062 29426
rect 46114 29374 46126 29426
rect 46610 29374 46622 29426
rect 46674 29374 46686 29426
rect 37774 29362 37826 29374
rect 47742 29362 47794 29374
rect 49758 29426 49810 29438
rect 49758 29362 49810 29374
rect 50654 29426 50706 29438
rect 51774 29426 51826 29438
rect 51426 29374 51438 29426
rect 51490 29374 51502 29426
rect 50654 29362 50706 29374
rect 51774 29362 51826 29374
rect 53566 29426 53618 29438
rect 54898 29374 54910 29426
rect 54962 29374 54974 29426
rect 53566 29362 53618 29374
rect 1934 29314 1986 29326
rect 1934 29250 1986 29262
rect 2270 29314 2322 29326
rect 2270 29250 2322 29262
rect 3726 29314 3778 29326
rect 3726 29250 3778 29262
rect 5742 29314 5794 29326
rect 5742 29250 5794 29262
rect 10894 29314 10946 29326
rect 13358 29314 13410 29326
rect 11666 29262 11678 29314
rect 11730 29262 11742 29314
rect 10894 29250 10946 29262
rect 13358 29250 13410 29262
rect 16270 29314 16322 29326
rect 16270 29250 16322 29262
rect 17614 29314 17666 29326
rect 17614 29250 17666 29262
rect 23998 29314 24050 29326
rect 23998 29250 24050 29262
rect 24894 29314 24946 29326
rect 24894 29250 24946 29262
rect 30606 29314 30658 29326
rect 34078 29314 34130 29326
rect 48190 29314 48242 29326
rect 32050 29262 32062 29314
rect 32114 29262 32126 29314
rect 45938 29262 45950 29314
rect 46002 29262 46014 29314
rect 30606 29250 30658 29262
rect 34078 29250 34130 29262
rect 48190 29250 48242 29262
rect 48862 29314 48914 29326
rect 52110 29314 52162 29326
rect 51314 29262 51326 29314
rect 51378 29262 51390 29314
rect 48862 29250 48914 29262
rect 52110 29250 52162 29262
rect 52558 29314 52610 29326
rect 52558 29250 52610 29262
rect 53006 29314 53058 29326
rect 56018 29262 56030 29314
rect 56082 29262 56094 29314
rect 53006 29250 53058 29262
rect 30494 29202 30546 29214
rect 2258 29150 2270 29202
rect 2322 29199 2334 29202
rect 3042 29199 3054 29202
rect 2322 29153 3054 29199
rect 2322 29150 2334 29153
rect 3042 29150 3054 29153
rect 3106 29150 3118 29202
rect 3378 29150 3390 29202
rect 3442 29199 3454 29202
rect 4946 29199 4958 29202
rect 3442 29153 4958 29199
rect 3442 29150 3454 29153
rect 4946 29150 4958 29153
rect 5010 29150 5022 29202
rect 5394 29150 5406 29202
rect 5458 29199 5470 29202
rect 5730 29199 5742 29202
rect 5458 29153 5742 29199
rect 5458 29150 5470 29153
rect 5730 29150 5742 29153
rect 5794 29150 5806 29202
rect 30494 29138 30546 29150
rect 35422 29202 35474 29214
rect 35422 29138 35474 29150
rect 44718 29202 44770 29214
rect 44718 29138 44770 29150
rect 49646 29202 49698 29214
rect 54238 29202 54290 29214
rect 52546 29150 52558 29202
rect 52610 29199 52622 29202
rect 53890 29199 53902 29202
rect 52610 29153 53902 29199
rect 52610 29150 52622 29153
rect 53890 29150 53902 29153
rect 53954 29150 53966 29202
rect 49646 29138 49698 29150
rect 54238 29138 54290 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 42478 28866 42530 28878
rect 3490 28814 3502 28866
rect 3554 28863 3566 28866
rect 4050 28863 4062 28866
rect 3554 28817 4062 28863
rect 3554 28814 3566 28817
rect 4050 28814 4062 28817
rect 4114 28814 4126 28866
rect 35634 28814 35646 28866
rect 35698 28863 35710 28866
rect 35970 28863 35982 28866
rect 35698 28817 35982 28863
rect 35698 28814 35710 28817
rect 35970 28814 35982 28817
rect 36034 28863 36046 28866
rect 36530 28863 36542 28866
rect 36034 28817 36542 28863
rect 36034 28814 36046 28817
rect 36530 28814 36542 28817
rect 36594 28814 36606 28866
rect 42478 28802 42530 28814
rect 48750 28866 48802 28878
rect 48750 28802 48802 28814
rect 2606 28754 2658 28766
rect 2606 28690 2658 28702
rect 3054 28754 3106 28766
rect 3054 28690 3106 28702
rect 3614 28754 3666 28766
rect 3614 28690 3666 28702
rect 4062 28754 4114 28766
rect 4062 28690 4114 28702
rect 19966 28754 20018 28766
rect 19966 28690 20018 28702
rect 22430 28754 22482 28766
rect 22430 28690 22482 28702
rect 25902 28754 25954 28766
rect 25902 28690 25954 28702
rect 26462 28754 26514 28766
rect 26462 28690 26514 28702
rect 28814 28754 28866 28766
rect 28814 28690 28866 28702
rect 29822 28754 29874 28766
rect 35758 28754 35810 28766
rect 30594 28702 30606 28754
rect 30658 28702 30670 28754
rect 32050 28702 32062 28754
rect 32114 28702 32126 28754
rect 29822 28690 29874 28702
rect 35758 28690 35810 28702
rect 36094 28754 36146 28766
rect 36094 28690 36146 28702
rect 36542 28754 36594 28766
rect 36542 28690 36594 28702
rect 40350 28754 40402 28766
rect 40350 28690 40402 28702
rect 46174 28754 46226 28766
rect 46174 28690 46226 28702
rect 46622 28754 46674 28766
rect 49870 28754 49922 28766
rect 48402 28702 48414 28754
rect 48466 28702 48478 28754
rect 46622 28690 46674 28702
rect 49870 28690 49922 28702
rect 50430 28754 50482 28766
rect 50430 28690 50482 28702
rect 52558 28754 52610 28766
rect 52558 28690 52610 28702
rect 4510 28642 4562 28654
rect 4510 28578 4562 28590
rect 4958 28642 5010 28654
rect 31726 28642 31778 28654
rect 14018 28590 14030 28642
rect 14082 28590 14094 28642
rect 14466 28590 14478 28642
rect 14530 28590 14542 28642
rect 16594 28590 16606 28642
rect 16658 28590 16670 28642
rect 30930 28590 30942 28642
rect 30994 28590 31006 28642
rect 4958 28578 5010 28590
rect 31726 28578 31778 28590
rect 32734 28642 32786 28654
rect 35198 28642 35250 28654
rect 34626 28590 34638 28642
rect 34690 28590 34702 28642
rect 32734 28578 32786 28590
rect 35198 28578 35250 28590
rect 37774 28642 37826 28654
rect 37774 28578 37826 28590
rect 38222 28642 38274 28654
rect 38222 28578 38274 28590
rect 40798 28642 40850 28654
rect 40798 28578 40850 28590
rect 41470 28642 41522 28654
rect 41470 28578 41522 28590
rect 42590 28642 42642 28654
rect 42590 28578 42642 28590
rect 42814 28642 42866 28654
rect 42814 28578 42866 28590
rect 49310 28642 49362 28654
rect 49310 28578 49362 28590
rect 50878 28642 50930 28654
rect 50878 28578 50930 28590
rect 52110 28642 52162 28654
rect 52110 28578 52162 28590
rect 53678 28642 53730 28654
rect 53678 28578 53730 28590
rect 54574 28642 54626 28654
rect 54574 28578 54626 28590
rect 55358 28642 55410 28654
rect 57598 28642 57650 28654
rect 56578 28590 56590 28642
rect 56642 28590 56654 28642
rect 55358 28578 55410 28590
rect 57598 28578 57650 28590
rect 58046 28642 58098 28654
rect 58046 28578 58098 28590
rect 25118 28530 25170 28542
rect 25118 28466 25170 28478
rect 25454 28530 25506 28542
rect 25454 28466 25506 28478
rect 27022 28530 27074 28542
rect 27022 28466 27074 28478
rect 27358 28530 27410 28542
rect 27358 28466 27410 28478
rect 30270 28530 30322 28542
rect 30270 28466 30322 28478
rect 32286 28530 32338 28542
rect 35086 28530 35138 28542
rect 33394 28478 33406 28530
rect 33458 28478 33470 28530
rect 32286 28466 32338 28478
rect 35086 28466 35138 28478
rect 41358 28530 41410 28542
rect 41358 28466 41410 28478
rect 43486 28530 43538 28542
rect 43486 28466 43538 28478
rect 44718 28530 44770 28542
rect 44718 28466 44770 28478
rect 45614 28530 45666 28542
rect 45614 28466 45666 28478
rect 45726 28530 45778 28542
rect 45726 28466 45778 28478
rect 48526 28530 48578 28542
rect 48526 28466 48578 28478
rect 51662 28530 51714 28542
rect 51662 28466 51714 28478
rect 53454 28530 53506 28542
rect 53454 28466 53506 28478
rect 54014 28530 54066 28542
rect 54014 28466 54066 28478
rect 56366 28530 56418 28542
rect 56366 28466 56418 28478
rect 57262 28530 57314 28542
rect 57262 28466 57314 28478
rect 2158 28418 2210 28430
rect 2158 28354 2210 28366
rect 17614 28418 17666 28430
rect 17614 28354 17666 28366
rect 18062 28418 18114 28430
rect 18062 28354 18114 28366
rect 32062 28418 32114 28430
rect 32062 28354 32114 28366
rect 33742 28418 33794 28430
rect 33742 28354 33794 28366
rect 34974 28418 35026 28430
rect 34974 28354 35026 28366
rect 37438 28418 37490 28430
rect 37438 28354 37490 28366
rect 37662 28418 37714 28430
rect 37662 28354 37714 28366
rect 41134 28418 41186 28430
rect 41134 28354 41186 28366
rect 42478 28418 42530 28430
rect 42478 28354 42530 28366
rect 43822 28418 43874 28430
rect 43822 28354 43874 28366
rect 44382 28418 44434 28430
rect 44382 28354 44434 28366
rect 45390 28418 45442 28430
rect 45390 28354 45442 28366
rect 47182 28418 47234 28430
rect 47182 28354 47234 28366
rect 47630 28418 47682 28430
rect 47630 28354 47682 28366
rect 51326 28418 51378 28430
rect 51326 28354 51378 28366
rect 53566 28418 53618 28430
rect 53566 28354 53618 28366
rect 55694 28418 55746 28430
rect 55694 28354 55746 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 3502 28082 3554 28094
rect 3502 28018 3554 28030
rect 4062 28082 4114 28094
rect 4062 28018 4114 28030
rect 10334 28082 10386 28094
rect 10334 28018 10386 28030
rect 15486 28082 15538 28094
rect 15486 28018 15538 28030
rect 16942 28082 16994 28094
rect 26686 28082 26738 28094
rect 23986 28030 23998 28082
rect 24050 28030 24062 28082
rect 25666 28030 25678 28082
rect 25730 28030 25742 28082
rect 16942 28018 16994 28030
rect 26686 28018 26738 28030
rect 29710 28082 29762 28094
rect 29710 28018 29762 28030
rect 32510 28082 32562 28094
rect 32510 28018 32562 28030
rect 33630 28082 33682 28094
rect 33630 28018 33682 28030
rect 37550 28082 37602 28094
rect 37550 28018 37602 28030
rect 44046 28082 44098 28094
rect 44046 28018 44098 28030
rect 47854 28082 47906 28094
rect 47854 28018 47906 28030
rect 49646 28082 49698 28094
rect 49646 28018 49698 28030
rect 50206 28082 50258 28094
rect 50206 28018 50258 28030
rect 51774 28082 51826 28094
rect 51774 28018 51826 28030
rect 53902 28082 53954 28094
rect 53902 28018 53954 28030
rect 54686 28082 54738 28094
rect 54686 28018 54738 28030
rect 19182 27970 19234 27982
rect 14578 27918 14590 27970
rect 14642 27918 14654 27970
rect 19182 27906 19234 27918
rect 28142 27970 28194 27982
rect 28142 27906 28194 27918
rect 28478 27970 28530 27982
rect 38446 27970 38498 27982
rect 29362 27918 29374 27970
rect 29426 27918 29438 27970
rect 31266 27918 31278 27970
rect 31330 27918 31342 27970
rect 35746 27918 35758 27970
rect 35810 27918 35822 27970
rect 28478 27906 28530 27918
rect 38446 27906 38498 27918
rect 39678 27970 39730 27982
rect 39678 27906 39730 27918
rect 40686 27970 40738 27982
rect 40686 27906 40738 27918
rect 40798 27970 40850 27982
rect 40798 27906 40850 27918
rect 41582 27970 41634 27982
rect 41582 27906 41634 27918
rect 42478 27970 42530 27982
rect 42478 27906 42530 27918
rect 46958 27970 47010 27982
rect 46958 27906 47010 27918
rect 47966 27970 48018 27982
rect 47966 27906 48018 27918
rect 48190 27970 48242 27982
rect 48190 27906 48242 27918
rect 49758 27970 49810 27982
rect 56366 27970 56418 27982
rect 52994 27918 53006 27970
rect 53058 27918 53070 27970
rect 55458 27918 55470 27970
rect 55522 27918 55534 27970
rect 49758 27906 49810 27918
rect 56366 27906 56418 27918
rect 57374 27970 57426 27982
rect 57374 27906 57426 27918
rect 14926 27858 14978 27870
rect 3042 27806 3054 27858
rect 3106 27806 3118 27858
rect 11330 27806 11342 27858
rect 11394 27806 11406 27858
rect 13458 27806 13470 27858
rect 13522 27806 13534 27858
rect 14018 27806 14030 27858
rect 14082 27806 14094 27858
rect 14926 27794 14978 27806
rect 17726 27858 17778 27870
rect 17726 27794 17778 27806
rect 17950 27858 18002 27870
rect 18846 27858 18898 27870
rect 18274 27806 18286 27858
rect 18338 27806 18350 27858
rect 17950 27794 18002 27806
rect 18846 27794 18898 27806
rect 21310 27858 21362 27870
rect 26238 27858 26290 27870
rect 21634 27806 21646 27858
rect 21698 27806 21710 27858
rect 21310 27794 21362 27806
rect 26238 27794 26290 27806
rect 33966 27858 34018 27870
rect 33966 27794 34018 27806
rect 35086 27858 35138 27870
rect 38110 27858 38162 27870
rect 35970 27806 35982 27858
rect 36034 27806 36046 27858
rect 35086 27794 35138 27806
rect 38110 27794 38162 27806
rect 40014 27858 40066 27870
rect 40014 27794 40066 27806
rect 40462 27858 40514 27870
rect 40462 27794 40514 27806
rect 41918 27858 41970 27870
rect 43822 27858 43874 27870
rect 42690 27806 42702 27858
rect 42754 27806 42766 27858
rect 43250 27806 43262 27858
rect 43314 27806 43326 27858
rect 41918 27794 41970 27806
rect 43822 27794 43874 27806
rect 44494 27858 44546 27870
rect 46846 27858 46898 27870
rect 45602 27806 45614 27858
rect 45666 27806 45678 27858
rect 46386 27806 46398 27858
rect 46450 27806 46462 27858
rect 44494 27794 44546 27806
rect 46846 27794 46898 27806
rect 47630 27858 47682 27870
rect 47630 27794 47682 27806
rect 49422 27858 49474 27870
rect 51886 27858 51938 27870
rect 56702 27858 56754 27870
rect 51650 27806 51662 27858
rect 51714 27806 51726 27858
rect 53218 27806 53230 27858
rect 53282 27806 53294 27858
rect 55682 27806 55694 27858
rect 55746 27806 55758 27858
rect 49422 27794 49474 27806
rect 51886 27794 51938 27806
rect 56702 27794 56754 27806
rect 15822 27746 15874 27758
rect 1922 27694 1934 27746
rect 1986 27694 1998 27746
rect 15822 27682 15874 27694
rect 16270 27746 16322 27758
rect 36542 27746 36594 27758
rect 30258 27694 30270 27746
rect 30322 27694 30334 27746
rect 16270 27682 16322 27694
rect 36542 27682 36594 27694
rect 36990 27746 37042 27758
rect 36990 27682 37042 27694
rect 39006 27746 39058 27758
rect 39006 27682 39058 27694
rect 42590 27746 42642 27758
rect 42590 27682 42642 27694
rect 43934 27746 43986 27758
rect 48638 27746 48690 27758
rect 45714 27694 45726 27746
rect 45778 27694 45790 27746
rect 43934 27682 43986 27694
rect 48638 27682 48690 27694
rect 52334 27746 52386 27758
rect 52334 27682 52386 27694
rect 54238 27746 54290 27758
rect 54238 27682 54290 27694
rect 57822 27746 57874 27758
rect 57822 27682 57874 27694
rect 24782 27634 24834 27646
rect 24782 27570 24834 27582
rect 26014 27634 26066 27646
rect 26014 27570 26066 27582
rect 34638 27634 34690 27646
rect 34638 27570 34690 27582
rect 34750 27634 34802 27646
rect 34750 27570 34802 27582
rect 34974 27634 35026 27646
rect 46958 27634 47010 27646
rect 43026 27582 43038 27634
rect 43090 27582 43102 27634
rect 45490 27582 45502 27634
rect 45554 27582 45566 27634
rect 34974 27570 35026 27582
rect 46958 27570 47010 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 56590 27298 56642 27310
rect 43698 27246 43710 27298
rect 43762 27295 43774 27298
rect 44034 27295 44046 27298
rect 43762 27249 44046 27295
rect 43762 27246 43774 27249
rect 44034 27246 44046 27249
rect 44098 27246 44110 27298
rect 56242 27246 56254 27298
rect 56306 27246 56318 27298
rect 56590 27234 56642 27246
rect 2158 27186 2210 27198
rect 18510 27186 18562 27198
rect 15138 27134 15150 27186
rect 15202 27134 15214 27186
rect 2158 27122 2210 27134
rect 18510 27122 18562 27134
rect 26126 27186 26178 27198
rect 26126 27122 26178 27134
rect 28142 27186 28194 27198
rect 28142 27122 28194 27134
rect 28590 27186 28642 27198
rect 28590 27122 28642 27134
rect 30046 27186 30098 27198
rect 30046 27122 30098 27134
rect 30382 27186 30434 27198
rect 30382 27122 30434 27134
rect 30942 27186 30994 27198
rect 30942 27122 30994 27134
rect 31390 27186 31442 27198
rect 31390 27122 31442 27134
rect 32734 27186 32786 27198
rect 32734 27122 32786 27134
rect 39678 27186 39730 27198
rect 39678 27122 39730 27134
rect 43150 27186 43202 27198
rect 43150 27122 43202 27134
rect 43598 27186 43650 27198
rect 43598 27122 43650 27134
rect 44158 27186 44210 27198
rect 56814 27186 56866 27198
rect 48178 27134 48190 27186
rect 48242 27134 48254 27186
rect 44158 27122 44210 27134
rect 56814 27122 56866 27134
rect 11006 27074 11058 27086
rect 11006 27010 11058 27022
rect 25678 27074 25730 27086
rect 25678 27010 25730 27022
rect 26686 27074 26738 27086
rect 26686 27010 26738 27022
rect 27470 27074 27522 27086
rect 27470 27010 27522 27022
rect 28030 27074 28082 27086
rect 37662 27074 37714 27086
rect 34066 27022 34078 27074
rect 34130 27022 34142 27074
rect 34850 27022 34862 27074
rect 34914 27022 34926 27074
rect 35746 27022 35758 27074
rect 35810 27022 35822 27074
rect 28030 27010 28082 27022
rect 37662 27010 37714 27022
rect 37998 27074 38050 27086
rect 37998 27010 38050 27022
rect 38222 27074 38274 27086
rect 38222 27010 38274 27022
rect 38894 27074 38946 27086
rect 38894 27010 38946 27022
rect 41582 27074 41634 27086
rect 41582 27010 41634 27022
rect 41918 27074 41970 27086
rect 41918 27010 41970 27022
rect 46062 27074 46114 27086
rect 49086 27074 49138 27086
rect 47058 27022 47070 27074
rect 47122 27022 47134 27074
rect 46062 27010 46114 27022
rect 49086 27010 49138 27022
rect 49310 27074 49362 27086
rect 51662 27074 51714 27086
rect 50194 27022 50206 27074
rect 50258 27022 50270 27074
rect 49310 27010 49362 27022
rect 51662 27010 51714 27022
rect 52670 27074 52722 27086
rect 54350 27074 54402 27086
rect 53554 27022 53566 27074
rect 53618 27022 53630 27074
rect 52670 27010 52722 27022
rect 54350 27010 54402 27022
rect 57710 27074 57762 27086
rect 57710 27010 57762 27022
rect 13022 26962 13074 26974
rect 17166 26962 17218 26974
rect 13794 26910 13806 26962
rect 13858 26910 13870 26962
rect 13022 26898 13074 26910
rect 17166 26898 17218 26910
rect 21982 26962 22034 26974
rect 21982 26898 22034 26910
rect 24558 26962 24610 26974
rect 24558 26898 24610 26910
rect 27246 26962 27298 26974
rect 36878 26962 36930 26974
rect 33954 26910 33966 26962
rect 34018 26910 34030 26962
rect 34626 26910 34638 26962
rect 34690 26910 34702 26962
rect 27246 26898 27298 26910
rect 36878 26898 36930 26910
rect 37774 26962 37826 26974
rect 37774 26898 37826 26910
rect 38670 26962 38722 26974
rect 38670 26898 38722 26910
rect 39230 26962 39282 26974
rect 39230 26898 39282 26910
rect 41358 26962 41410 26974
rect 41358 26898 41410 26910
rect 42366 26962 42418 26974
rect 42366 26898 42418 26910
rect 42702 26962 42754 26974
rect 42702 26898 42754 26910
rect 44494 26962 44546 26974
rect 44494 26898 44546 26910
rect 45614 26962 45666 26974
rect 45614 26898 45666 26910
rect 47742 26962 47794 26974
rect 47742 26898 47794 26910
rect 49198 26962 49250 26974
rect 55582 26962 55634 26974
rect 50418 26910 50430 26962
rect 50482 26910 50494 26962
rect 49198 26898 49250 26910
rect 55582 26898 55634 26910
rect 11342 26850 11394 26862
rect 25342 26850 25394 26862
rect 21634 26798 21646 26850
rect 21698 26798 21710 26850
rect 24882 26798 24894 26850
rect 24946 26798 24958 26850
rect 11342 26786 11394 26798
rect 25342 26786 25394 26798
rect 25566 26850 25618 26862
rect 25566 26786 25618 26798
rect 32174 26850 32226 26862
rect 36318 26850 36370 26862
rect 34290 26798 34302 26850
rect 34354 26798 34366 26850
rect 32174 26786 32226 26798
rect 36318 26786 36370 26798
rect 39006 26850 39058 26862
rect 39006 26786 39058 26798
rect 40126 26850 40178 26862
rect 40126 26786 40178 26798
rect 40798 26850 40850 26862
rect 40798 26786 40850 26798
rect 41582 26850 41634 26862
rect 41582 26786 41634 26798
rect 42590 26850 42642 26862
rect 42590 26786 42642 26798
rect 45838 26850 45890 26862
rect 45838 26786 45890 26798
rect 45950 26850 46002 26862
rect 51326 26850 51378 26862
rect 46834 26798 46846 26850
rect 46898 26798 46910 26850
rect 50194 26798 50206 26850
rect 50258 26798 50270 26850
rect 45950 26786 46002 26798
rect 51326 26786 51378 26798
rect 52334 26850 52386 26862
rect 52334 26786 52386 26798
rect 53790 26850 53842 26862
rect 53790 26786 53842 26798
rect 54686 26850 54738 26862
rect 54686 26786 54738 26798
rect 55246 26850 55298 26862
rect 55246 26786 55298 26798
rect 57374 26850 57426 26862
rect 57374 26786 57426 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 25006 26514 25058 26526
rect 16258 26462 16270 26514
rect 16322 26462 16334 26514
rect 24434 26462 24446 26514
rect 24498 26462 24510 26514
rect 25006 26450 25058 26462
rect 25678 26514 25730 26526
rect 25678 26450 25730 26462
rect 26350 26514 26402 26526
rect 33518 26514 33570 26526
rect 27682 26462 27694 26514
rect 27746 26462 27758 26514
rect 31490 26462 31502 26514
rect 31554 26462 31566 26514
rect 26350 26450 26402 26462
rect 33518 26450 33570 26462
rect 34750 26514 34802 26526
rect 34750 26450 34802 26462
rect 35422 26514 35474 26526
rect 35422 26450 35474 26462
rect 37102 26514 37154 26526
rect 37102 26450 37154 26462
rect 37662 26514 37714 26526
rect 37662 26450 37714 26462
rect 38446 26514 38498 26526
rect 38446 26450 38498 26462
rect 38894 26514 38946 26526
rect 38894 26450 38946 26462
rect 41582 26514 41634 26526
rect 41582 26450 41634 26462
rect 43374 26514 43426 26526
rect 43374 26450 43426 26462
rect 46622 26514 46674 26526
rect 46622 26450 46674 26462
rect 47518 26514 47570 26526
rect 47518 26450 47570 26462
rect 48526 26514 48578 26526
rect 48526 26450 48578 26462
rect 18062 26402 18114 26414
rect 35982 26402 36034 26414
rect 32050 26350 32062 26402
rect 32114 26350 32126 26402
rect 18062 26338 18114 26350
rect 35982 26338 36034 26350
rect 37998 26402 38050 26414
rect 37998 26338 38050 26350
rect 39790 26402 39842 26414
rect 48750 26402 48802 26414
rect 43922 26350 43934 26402
rect 43986 26350 43998 26402
rect 39790 26338 39842 26350
rect 48750 26338 48802 26350
rect 54910 26402 54962 26414
rect 57374 26402 57426 26414
rect 56018 26350 56030 26402
rect 56082 26350 56094 26402
rect 54910 26338 54962 26350
rect 57374 26338 57426 26350
rect 13582 26290 13634 26302
rect 18398 26290 18450 26302
rect 14018 26238 14030 26290
rect 14082 26238 14094 26290
rect 13582 26226 13634 26238
rect 18398 26226 18450 26238
rect 18958 26290 19010 26302
rect 19854 26290 19906 26302
rect 19618 26238 19630 26290
rect 19682 26238 19694 26290
rect 18958 26226 19010 26238
rect 19854 26226 19906 26238
rect 20414 26290 20466 26302
rect 20414 26226 20466 26238
rect 21310 26290 21362 26302
rect 30606 26290 30658 26302
rect 35534 26290 35586 26302
rect 21858 26238 21870 26290
rect 21922 26238 21934 26290
rect 29922 26238 29934 26290
rect 29986 26238 29998 26290
rect 31602 26238 31614 26290
rect 31666 26238 31678 26290
rect 32498 26238 32510 26290
rect 32562 26238 32574 26290
rect 34514 26238 34526 26290
rect 34578 26238 34590 26290
rect 21310 26226 21362 26238
rect 30606 26226 30658 26238
rect 35534 26226 35586 26238
rect 36542 26290 36594 26302
rect 39342 26290 39394 26302
rect 47070 26290 47122 26302
rect 50766 26290 50818 26302
rect 36866 26238 36878 26290
rect 36930 26238 36942 26290
rect 44258 26238 44270 26290
rect 44322 26238 44334 26290
rect 44818 26238 44830 26290
rect 44882 26238 44894 26290
rect 45826 26238 45838 26290
rect 45890 26238 45902 26290
rect 46162 26238 46174 26290
rect 46226 26238 46238 26290
rect 48290 26238 48302 26290
rect 48354 26238 48366 26290
rect 36542 26226 36594 26238
rect 39342 26226 39394 26238
rect 47070 26226 47122 26238
rect 50766 26226 50818 26238
rect 52670 26290 52722 26302
rect 53442 26238 53454 26290
rect 53506 26238 53518 26290
rect 53666 26238 53678 26290
rect 53730 26238 53742 26290
rect 56242 26238 56254 26290
rect 56306 26238 56318 26290
rect 52670 26226 52722 26238
rect 20862 26178 20914 26190
rect 20862 26114 20914 26126
rect 40350 26178 40402 26190
rect 40350 26114 40402 26126
rect 40686 26178 40738 26190
rect 40686 26114 40738 26126
rect 42142 26178 42194 26190
rect 42142 26114 42194 26126
rect 42590 26178 42642 26190
rect 42590 26114 42642 26126
rect 49422 26178 49474 26190
rect 49422 26114 49474 26126
rect 49870 26178 49922 26190
rect 49870 26114 49922 26126
rect 50990 26178 51042 26190
rect 50990 26114 51042 26126
rect 51550 26178 51602 26190
rect 54462 26178 54514 26190
rect 53106 26126 53118 26178
rect 53170 26126 53182 26178
rect 51550 26114 51602 26126
rect 54462 26114 54514 26126
rect 55358 26178 55410 26190
rect 55358 26114 55410 26126
rect 57822 26178 57874 26190
rect 57822 26114 57874 26126
rect 17054 26066 17106 26078
rect 17054 26002 17106 26014
rect 26126 26066 26178 26078
rect 26126 26002 26178 26014
rect 26910 26066 26962 26078
rect 26910 26002 26962 26014
rect 35422 26066 35474 26078
rect 35422 26002 35474 26014
rect 37214 26066 37266 26078
rect 37214 26002 37266 26014
rect 44270 26066 44322 26078
rect 44270 26002 44322 26014
rect 48862 26066 48914 26078
rect 48862 26002 48914 26014
rect 50430 26066 50482 26078
rect 50430 26002 50482 26014
rect 51774 26066 51826 26078
rect 51774 26002 51826 26014
rect 52110 26066 52162 26078
rect 57922 26014 57934 26066
rect 57986 26063 57998 26066
rect 58258 26063 58270 26066
rect 57986 26017 58270 26063
rect 57986 26014 57998 26017
rect 58258 26014 58270 26017
rect 58322 26014 58334 26066
rect 52110 26002 52162 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 20974 25730 21026 25742
rect 20974 25666 21026 25678
rect 28142 25730 28194 25742
rect 28142 25666 28194 25678
rect 35646 25730 35698 25742
rect 35646 25666 35698 25678
rect 35870 25730 35922 25742
rect 35870 25666 35922 25678
rect 37550 25730 37602 25742
rect 37550 25666 37602 25678
rect 38110 25730 38162 25742
rect 38110 25666 38162 25678
rect 38334 25730 38386 25742
rect 57598 25730 57650 25742
rect 48850 25678 48862 25730
rect 48914 25727 48926 25730
rect 49634 25727 49646 25730
rect 48914 25681 49646 25727
rect 48914 25678 48926 25681
rect 49634 25678 49646 25681
rect 49698 25678 49710 25730
rect 50866 25678 50878 25730
rect 50930 25727 50942 25730
rect 51426 25727 51438 25730
rect 50930 25681 51438 25727
rect 50930 25678 50942 25681
rect 51426 25678 51438 25681
rect 51490 25678 51502 25730
rect 38334 25666 38386 25678
rect 57598 25666 57650 25678
rect 16046 25618 16098 25630
rect 27022 25618 27074 25630
rect 41806 25618 41858 25630
rect 26002 25566 26014 25618
rect 26066 25566 26078 25618
rect 31490 25566 31502 25618
rect 31554 25566 31566 25618
rect 16046 25554 16098 25566
rect 27022 25554 27074 25566
rect 41806 25554 41858 25566
rect 43150 25618 43202 25630
rect 49534 25618 49586 25630
rect 47394 25566 47406 25618
rect 47458 25566 47470 25618
rect 43150 25554 43202 25566
rect 49534 25554 49586 25566
rect 51326 25618 51378 25630
rect 51326 25554 51378 25566
rect 51774 25618 51826 25630
rect 51774 25554 51826 25566
rect 52334 25618 52386 25630
rect 52334 25554 52386 25566
rect 52670 25618 52722 25630
rect 56354 25566 56366 25618
rect 56418 25566 56430 25618
rect 52670 25554 52722 25566
rect 15598 25506 15650 25518
rect 14578 25454 14590 25506
rect 14642 25454 14654 25506
rect 15598 25442 15650 25454
rect 17502 25506 17554 25518
rect 27806 25506 27858 25518
rect 17938 25454 17950 25506
rect 18002 25454 18014 25506
rect 27570 25454 27582 25506
rect 27634 25454 27646 25506
rect 17502 25442 17554 25454
rect 27806 25442 27858 25454
rect 28030 25506 28082 25518
rect 33966 25506 34018 25518
rect 31154 25454 31166 25506
rect 31218 25454 31230 25506
rect 28030 25442 28082 25454
rect 33966 25442 34018 25454
rect 35422 25506 35474 25518
rect 35422 25442 35474 25454
rect 37662 25506 37714 25518
rect 37662 25442 37714 25454
rect 38894 25506 38946 25518
rect 38894 25442 38946 25454
rect 39118 25506 39170 25518
rect 39118 25442 39170 25454
rect 39342 25506 39394 25518
rect 39342 25442 39394 25454
rect 40574 25506 40626 25518
rect 40574 25442 40626 25454
rect 43822 25506 43874 25518
rect 43822 25442 43874 25454
rect 44158 25506 44210 25518
rect 53790 25506 53842 25518
rect 47730 25454 47742 25506
rect 47794 25454 47806 25506
rect 44158 25442 44210 25454
rect 53790 25442 53842 25454
rect 55134 25506 55186 25518
rect 56466 25454 56478 25506
rect 56530 25454 56542 25506
rect 57922 25454 57934 25506
rect 57986 25454 57998 25506
rect 55134 25442 55186 25454
rect 14366 25394 14418 25406
rect 31838 25394 31890 25406
rect 15250 25342 15262 25394
rect 15314 25342 15326 25394
rect 24658 25342 24670 25394
rect 24722 25342 24734 25394
rect 14366 25330 14418 25342
rect 31838 25330 31890 25342
rect 32398 25394 32450 25406
rect 32398 25330 32450 25342
rect 32622 25394 32674 25406
rect 32622 25330 32674 25342
rect 32734 25394 32786 25406
rect 33742 25394 33794 25406
rect 32834 25342 32846 25394
rect 32898 25342 32910 25394
rect 32734 25330 32786 25342
rect 33742 25330 33794 25342
rect 34302 25394 34354 25406
rect 34302 25330 34354 25342
rect 36430 25394 36482 25406
rect 36430 25330 36482 25342
rect 36766 25394 36818 25406
rect 36766 25330 36818 25342
rect 37886 25394 37938 25406
rect 37886 25330 37938 25342
rect 39566 25394 39618 25406
rect 39566 25330 39618 25342
rect 40238 25394 40290 25406
rect 40238 25330 40290 25342
rect 41134 25394 41186 25406
rect 41134 25330 41186 25342
rect 43038 25394 43090 25406
rect 43038 25330 43090 25342
rect 43262 25394 43314 25406
rect 43262 25330 43314 25342
rect 44494 25394 44546 25406
rect 44494 25330 44546 25342
rect 46174 25394 46226 25406
rect 46174 25330 46226 25342
rect 46846 25394 46898 25406
rect 47966 25394 48018 25406
rect 47618 25342 47630 25394
rect 47682 25342 47694 25394
rect 46846 25330 46898 25342
rect 47966 25330 48018 25342
rect 50430 25394 50482 25406
rect 50430 25330 50482 25342
rect 50878 25394 50930 25406
rect 50878 25330 50930 25342
rect 54238 25394 54290 25406
rect 54238 25330 54290 25342
rect 56030 25394 56082 25406
rect 56030 25330 56082 25342
rect 21534 25282 21586 25294
rect 20402 25230 20414 25282
rect 20466 25230 20478 25282
rect 21534 25218 21586 25230
rect 24110 25282 24162 25294
rect 24110 25218 24162 25230
rect 26462 25282 26514 25294
rect 26462 25218 26514 25230
rect 28590 25282 28642 25294
rect 28590 25218 28642 25230
rect 30046 25282 30098 25294
rect 30046 25218 30098 25230
rect 32510 25282 32562 25294
rect 32510 25218 32562 25230
rect 33966 25282 34018 25294
rect 33966 25218 34018 25230
rect 34974 25282 35026 25294
rect 34974 25218 35026 25230
rect 35086 25282 35138 25294
rect 35086 25218 35138 25230
rect 35198 25282 35250 25294
rect 35198 25218 35250 25230
rect 41246 25282 41298 25294
rect 41246 25218 41298 25230
rect 41470 25282 41522 25294
rect 41470 25218 41522 25230
rect 42254 25282 42306 25294
rect 42254 25218 42306 25230
rect 44046 25282 44098 25294
rect 44046 25218 44098 25230
rect 45838 25282 45890 25294
rect 45838 25218 45890 25230
rect 46734 25282 46786 25294
rect 46734 25218 46786 25230
rect 48190 25282 48242 25294
rect 48190 25218 48242 25230
rect 48638 25282 48690 25294
rect 48638 25218 48690 25230
rect 49086 25282 49138 25294
rect 49086 25218 49138 25230
rect 50094 25282 50146 25294
rect 54798 25282 54850 25294
rect 53442 25230 53454 25282
rect 53506 25230 53518 25282
rect 50094 25218 50146 25230
rect 54798 25218 54850 25230
rect 57710 25282 57762 25294
rect 57710 25218 57762 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 14366 24946 14418 24958
rect 14366 24882 14418 24894
rect 21422 24946 21474 24958
rect 21422 24882 21474 24894
rect 21870 24946 21922 24958
rect 21870 24882 21922 24894
rect 25902 24946 25954 24958
rect 25902 24882 25954 24894
rect 27582 24946 27634 24958
rect 27582 24882 27634 24894
rect 29710 24946 29762 24958
rect 29710 24882 29762 24894
rect 30270 24946 30322 24958
rect 30270 24882 30322 24894
rect 31390 24946 31442 24958
rect 31390 24882 31442 24894
rect 32734 24946 32786 24958
rect 32734 24882 32786 24894
rect 34302 24946 34354 24958
rect 34302 24882 34354 24894
rect 37774 24946 37826 24958
rect 37774 24882 37826 24894
rect 38222 24946 38274 24958
rect 38222 24882 38274 24894
rect 40574 24946 40626 24958
rect 40574 24882 40626 24894
rect 43822 24946 43874 24958
rect 43822 24882 43874 24894
rect 46846 24946 46898 24958
rect 46846 24882 46898 24894
rect 48078 24946 48130 24958
rect 48078 24882 48130 24894
rect 51774 24946 51826 24958
rect 51774 24882 51826 24894
rect 52334 24946 52386 24958
rect 52334 24882 52386 24894
rect 52782 24946 52834 24958
rect 52782 24882 52834 24894
rect 57486 24946 57538 24958
rect 57486 24882 57538 24894
rect 14702 24834 14754 24846
rect 14702 24770 14754 24782
rect 15262 24834 15314 24846
rect 24670 24834 24722 24846
rect 18834 24782 18846 24834
rect 18898 24782 18910 24834
rect 22866 24782 22878 24834
rect 22930 24782 22942 24834
rect 15262 24770 15314 24782
rect 24670 24770 24722 24782
rect 26910 24834 26962 24846
rect 26910 24770 26962 24782
rect 27022 24834 27074 24846
rect 27022 24770 27074 24782
rect 29822 24834 29874 24846
rect 29822 24770 29874 24782
rect 36766 24834 36818 24846
rect 36766 24770 36818 24782
rect 37326 24834 37378 24846
rect 37326 24770 37378 24782
rect 38670 24834 38722 24846
rect 38670 24770 38722 24782
rect 40126 24834 40178 24846
rect 40126 24770 40178 24782
rect 46062 24834 46114 24846
rect 47182 24834 47234 24846
rect 46946 24782 46958 24834
rect 47010 24782 47022 24834
rect 46062 24770 46114 24782
rect 47182 24770 47234 24782
rect 49982 24834 50034 24846
rect 49982 24770 50034 24782
rect 51102 24834 51154 24846
rect 54798 24834 54850 24846
rect 53890 24782 53902 24834
rect 53954 24782 53966 24834
rect 51102 24770 51154 24782
rect 54798 24770 54850 24782
rect 55134 24834 55186 24846
rect 55134 24770 55186 24782
rect 56030 24834 56082 24846
rect 56030 24770 56082 24782
rect 25678 24722 25730 24734
rect 25678 24658 25730 24670
rect 26350 24722 26402 24734
rect 26350 24658 26402 24670
rect 26686 24722 26738 24734
rect 26686 24658 26738 24670
rect 27918 24722 27970 24734
rect 27918 24658 27970 24670
rect 31950 24722 32002 24734
rect 31950 24658 32002 24670
rect 33630 24722 33682 24734
rect 34078 24722 34130 24734
rect 35646 24722 35698 24734
rect 33954 24670 33966 24722
rect 34018 24670 34030 24722
rect 35186 24670 35198 24722
rect 35250 24670 35262 24722
rect 33630 24658 33682 24670
rect 34078 24658 34130 24670
rect 35646 24658 35698 24670
rect 35870 24722 35922 24734
rect 39678 24722 39730 24734
rect 39442 24670 39454 24722
rect 39506 24670 39518 24722
rect 35870 24658 35922 24670
rect 39678 24658 39730 24670
rect 39902 24722 39954 24734
rect 39902 24658 39954 24670
rect 42254 24722 42306 24734
rect 42254 24658 42306 24670
rect 42926 24722 42978 24734
rect 42926 24658 42978 24670
rect 43934 24722 43986 24734
rect 43934 24658 43986 24670
rect 44158 24722 44210 24734
rect 45726 24722 45778 24734
rect 44370 24670 44382 24722
rect 44434 24670 44446 24722
rect 45490 24670 45502 24722
rect 45554 24670 45566 24722
rect 44158 24658 44210 24670
rect 45726 24658 45778 24670
rect 46734 24722 46786 24734
rect 46734 24658 46786 24670
rect 49646 24722 49698 24734
rect 49646 24658 49698 24670
rect 49758 24722 49810 24734
rect 49758 24658 49810 24670
rect 50206 24722 50258 24734
rect 51886 24722 51938 24734
rect 56366 24722 56418 24734
rect 50866 24670 50878 24722
rect 50930 24670 50942 24722
rect 54114 24670 54126 24722
rect 54178 24670 54190 24722
rect 50206 24658 50258 24670
rect 51886 24658 51938 24670
rect 56366 24658 56418 24670
rect 56590 24722 56642 24734
rect 56590 24658 56642 24670
rect 58046 24722 58098 24734
rect 58046 24658 58098 24670
rect 20638 24610 20690 24622
rect 20638 24546 20690 24558
rect 25790 24610 25842 24622
rect 25790 24546 25842 24558
rect 30830 24610 30882 24622
rect 30830 24546 30882 24558
rect 34190 24610 34242 24622
rect 34190 24546 34242 24558
rect 36654 24610 36706 24622
rect 36654 24546 36706 24558
rect 39790 24610 39842 24622
rect 39790 24546 39842 24558
rect 41470 24610 41522 24622
rect 44046 24610 44098 24622
rect 42690 24558 42702 24610
rect 42754 24558 42766 24610
rect 41470 24546 41522 24558
rect 44046 24546 44098 24558
rect 45950 24610 46002 24622
rect 45950 24546 46002 24558
rect 47630 24610 47682 24622
rect 47630 24546 47682 24558
rect 48526 24610 48578 24622
rect 48526 24546 48578 24558
rect 53230 24610 53282 24622
rect 56130 24558 56142 24610
rect 56194 24558 56206 24610
rect 53230 24546 53282 24558
rect 29710 24498 29762 24510
rect 29710 24434 29762 24446
rect 31838 24498 31890 24510
rect 31838 24434 31890 24446
rect 32398 24498 32450 24510
rect 32398 24434 32450 24446
rect 32622 24498 32674 24510
rect 32622 24434 32674 24446
rect 35422 24498 35474 24510
rect 35422 24434 35474 24446
rect 35982 24498 36034 24510
rect 35982 24434 36034 24446
rect 36542 24498 36594 24510
rect 42478 24498 42530 24510
rect 37538 24446 37550 24498
rect 37602 24495 37614 24498
rect 37986 24495 37998 24498
rect 37602 24449 37998 24495
rect 37602 24446 37614 24449
rect 37986 24446 37998 24449
rect 38050 24446 38062 24498
rect 36542 24434 36594 24446
rect 42478 24434 42530 24446
rect 43038 24498 43090 24510
rect 43038 24434 43090 24446
rect 45614 24498 45666 24510
rect 45614 24434 45666 24446
rect 47518 24498 47570 24510
rect 47518 24434 47570 24446
rect 49646 24498 49698 24510
rect 49646 24434 49698 24446
rect 51774 24498 51826 24510
rect 55806 24498 55858 24510
rect 52098 24446 52110 24498
rect 52162 24495 52174 24498
rect 52994 24495 53006 24498
rect 52162 24449 53006 24495
rect 52162 24446 52174 24449
rect 52994 24446 53006 24449
rect 53058 24495 53070 24498
rect 53666 24495 53678 24498
rect 53058 24449 53678 24495
rect 53058 24446 53070 24449
rect 53666 24446 53678 24449
rect 53730 24446 53742 24498
rect 51774 24434 51826 24446
rect 55806 24434 55858 24446
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 38894 24162 38946 24174
rect 57150 24162 57202 24174
rect 39890 24110 39902 24162
rect 39954 24110 39966 24162
rect 38894 24098 38946 24110
rect 57150 24098 57202 24110
rect 57598 24162 57650 24174
rect 57598 24098 57650 24110
rect 22542 24050 22594 24062
rect 22542 23986 22594 23998
rect 23102 24050 23154 24062
rect 23102 23986 23154 23998
rect 24334 24050 24386 24062
rect 24334 23986 24386 23998
rect 27918 24050 27970 24062
rect 27918 23986 27970 23998
rect 30606 24050 30658 24062
rect 34190 24050 34242 24062
rect 47630 24050 47682 24062
rect 32162 23998 32174 24050
rect 32226 23998 32238 24050
rect 32946 23998 32958 24050
rect 33010 23998 33022 24050
rect 34962 23998 34974 24050
rect 35026 23998 35038 24050
rect 30606 23986 30658 23998
rect 34190 23986 34242 23998
rect 47630 23986 47682 23998
rect 50766 24050 50818 24062
rect 50766 23986 50818 23998
rect 56702 24050 56754 24062
rect 56702 23986 56754 23998
rect 17502 23938 17554 23950
rect 23214 23938 23266 23950
rect 17826 23886 17838 23938
rect 17890 23886 17902 23938
rect 21746 23886 21758 23938
rect 21810 23886 21822 23938
rect 17502 23874 17554 23886
rect 23214 23874 23266 23886
rect 29934 23938 29986 23950
rect 34078 23938 34130 23950
rect 31714 23886 31726 23938
rect 31778 23886 31790 23938
rect 32722 23886 32734 23938
rect 32786 23886 32798 23938
rect 29934 23874 29986 23886
rect 34078 23874 34130 23886
rect 35198 23938 35250 23950
rect 35198 23874 35250 23886
rect 38446 23938 38498 23950
rect 38446 23874 38498 23886
rect 38670 23938 38722 23950
rect 39454 23938 39506 23950
rect 39106 23886 39118 23938
rect 39170 23886 39182 23938
rect 38670 23874 38722 23886
rect 39454 23874 39506 23886
rect 40238 23938 40290 23950
rect 40238 23874 40290 23886
rect 40462 23938 40514 23950
rect 40462 23874 40514 23886
rect 40910 23938 40962 23950
rect 40910 23874 40962 23886
rect 41246 23938 41298 23950
rect 41246 23874 41298 23886
rect 41918 23938 41970 23950
rect 43710 23938 43762 23950
rect 42354 23886 42366 23938
rect 42418 23886 42430 23938
rect 42690 23886 42702 23938
rect 42754 23886 42766 23938
rect 41918 23874 41970 23886
rect 43710 23874 43762 23886
rect 46622 23938 46674 23950
rect 46622 23874 46674 23886
rect 46734 23938 46786 23950
rect 46734 23874 46786 23886
rect 46958 23938 47010 23950
rect 46958 23874 47010 23886
rect 48638 23938 48690 23950
rect 48638 23874 48690 23886
rect 49870 23938 49922 23950
rect 49870 23874 49922 23886
rect 50990 23938 51042 23950
rect 53454 23938 53506 23950
rect 52098 23886 52110 23938
rect 52162 23886 52174 23938
rect 52658 23886 52670 23938
rect 52722 23886 52734 23938
rect 50990 23874 51042 23886
rect 53454 23874 53506 23886
rect 53678 23938 53730 23950
rect 56926 23938 56978 23950
rect 55010 23886 55022 23938
rect 55074 23886 55086 23938
rect 53678 23874 53730 23886
rect 56926 23874 56978 23886
rect 22990 23826 23042 23838
rect 22990 23762 23042 23774
rect 23550 23826 23602 23838
rect 27470 23826 27522 23838
rect 26114 23774 26126 23826
rect 26178 23774 26190 23826
rect 23550 23762 23602 23774
rect 27470 23762 27522 23774
rect 33182 23826 33234 23838
rect 33182 23762 33234 23774
rect 35422 23826 35474 23838
rect 35422 23762 35474 23774
rect 35982 23826 36034 23838
rect 35982 23762 36034 23774
rect 36318 23826 36370 23838
rect 36318 23762 36370 23774
rect 37550 23826 37602 23838
rect 37550 23762 37602 23774
rect 37886 23826 37938 23838
rect 37886 23762 37938 23774
rect 43822 23826 43874 23838
rect 43822 23762 43874 23774
rect 43934 23826 43986 23838
rect 46286 23826 46338 23838
rect 44034 23774 44046 23826
rect 44098 23774 44110 23826
rect 43934 23762 43986 23774
rect 46286 23762 46338 23774
rect 47182 23826 47234 23838
rect 47182 23762 47234 23774
rect 48974 23826 49026 23838
rect 54014 23826 54066 23838
rect 51874 23774 51886 23826
rect 51938 23774 51950 23826
rect 56018 23774 56030 23826
rect 56082 23774 56094 23826
rect 48974 23762 49026 23774
rect 54014 23762 54066 23774
rect 20974 23714 21026 23726
rect 20402 23662 20414 23714
rect 20466 23662 20478 23714
rect 20974 23650 21026 23662
rect 21982 23714 22034 23726
rect 21982 23650 22034 23662
rect 27134 23714 27186 23726
rect 27134 23650 27186 23662
rect 28926 23714 28978 23726
rect 28926 23650 28978 23662
rect 30046 23714 30098 23726
rect 30046 23650 30098 23662
rect 30270 23714 30322 23726
rect 30270 23650 30322 23662
rect 34862 23714 34914 23726
rect 34862 23650 34914 23662
rect 34974 23714 35026 23726
rect 34974 23650 35026 23662
rect 36766 23714 36818 23726
rect 36766 23650 36818 23662
rect 38894 23714 38946 23726
rect 38894 23650 38946 23662
rect 41134 23714 41186 23726
rect 41134 23650 41186 23662
rect 42030 23714 42082 23726
rect 42030 23650 42082 23662
rect 42142 23714 42194 23726
rect 42142 23650 42194 23662
rect 43598 23714 43650 23726
rect 43598 23650 43650 23662
rect 45390 23714 45442 23726
rect 48190 23714 48242 23726
rect 46610 23662 46622 23714
rect 46674 23662 46686 23714
rect 45390 23650 45442 23662
rect 48190 23650 48242 23662
rect 48862 23714 48914 23726
rect 48862 23650 48914 23662
rect 49534 23714 49586 23726
rect 53902 23714 53954 23726
rect 50418 23662 50430 23714
rect 50482 23662 50494 23714
rect 52434 23662 52446 23714
rect 52498 23662 52510 23714
rect 49534 23650 49586 23662
rect 53902 23650 53954 23662
rect 57934 23714 57986 23726
rect 57934 23650 57986 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 17950 23378 18002 23390
rect 17950 23314 18002 23326
rect 20302 23378 20354 23390
rect 20302 23314 20354 23326
rect 23774 23378 23826 23390
rect 23774 23314 23826 23326
rect 24670 23378 24722 23390
rect 24670 23314 24722 23326
rect 30382 23378 30434 23390
rect 30382 23314 30434 23326
rect 31054 23378 31106 23390
rect 31054 23314 31106 23326
rect 33966 23378 34018 23390
rect 33966 23314 34018 23326
rect 36542 23378 36594 23390
rect 36542 23314 36594 23326
rect 37102 23378 37154 23390
rect 37102 23314 37154 23326
rect 37438 23378 37490 23390
rect 37438 23314 37490 23326
rect 38782 23378 38834 23390
rect 38782 23314 38834 23326
rect 39566 23378 39618 23390
rect 39566 23314 39618 23326
rect 41470 23378 41522 23390
rect 41470 23314 41522 23326
rect 44718 23378 44770 23390
rect 44718 23314 44770 23326
rect 45950 23378 46002 23390
rect 45950 23314 46002 23326
rect 46846 23378 46898 23390
rect 46846 23314 46898 23326
rect 47294 23378 47346 23390
rect 47294 23314 47346 23326
rect 47742 23378 47794 23390
rect 47742 23314 47794 23326
rect 48750 23378 48802 23390
rect 48750 23314 48802 23326
rect 51886 23378 51938 23390
rect 51886 23314 51938 23326
rect 52110 23378 52162 23390
rect 52110 23314 52162 23326
rect 55022 23378 55074 23390
rect 55022 23314 55074 23326
rect 55470 23378 55522 23390
rect 57486 23378 57538 23390
rect 56130 23326 56142 23378
rect 56194 23326 56206 23378
rect 55470 23314 55522 23326
rect 57486 23314 57538 23326
rect 24894 23266 24946 23278
rect 21298 23214 21310 23266
rect 21362 23214 21374 23266
rect 24894 23202 24946 23214
rect 27358 23266 27410 23278
rect 35870 23266 35922 23278
rect 53790 23266 53842 23278
rect 29138 23214 29150 23266
rect 29202 23214 29214 23266
rect 42802 23214 42814 23266
rect 42866 23214 42878 23266
rect 27358 23202 27410 23214
rect 35870 23202 35922 23214
rect 53790 23202 53842 23214
rect 19406 23154 19458 23166
rect 19170 23102 19182 23154
rect 19234 23102 19246 23154
rect 19406 23090 19458 23102
rect 20750 23154 20802 23166
rect 20750 23090 20802 23102
rect 25678 23154 25730 23166
rect 27246 23154 27298 23166
rect 26114 23102 26126 23154
rect 26178 23102 26190 23154
rect 25678 23090 25730 23102
rect 27246 23090 27298 23102
rect 27582 23154 27634 23166
rect 27582 23090 27634 23102
rect 28478 23154 28530 23166
rect 29934 23154 29986 23166
rect 29250 23102 29262 23154
rect 29314 23102 29326 23154
rect 28478 23090 28530 23102
rect 29934 23090 29986 23102
rect 30158 23154 30210 23166
rect 30158 23090 30210 23102
rect 31390 23154 31442 23166
rect 31390 23090 31442 23102
rect 34638 23154 34690 23166
rect 34638 23090 34690 23102
rect 34974 23154 35026 23166
rect 34974 23090 35026 23102
rect 35086 23154 35138 23166
rect 40350 23154 40402 23166
rect 40114 23102 40126 23154
rect 40178 23102 40190 23154
rect 35086 23090 35138 23102
rect 40350 23090 40402 23102
rect 40574 23154 40626 23166
rect 42478 23154 42530 23166
rect 40786 23102 40798 23154
rect 40850 23102 40862 23154
rect 40574 23090 40626 23102
rect 42478 23090 42530 23102
rect 49534 23154 49586 23166
rect 49534 23090 49586 23102
rect 49758 23154 49810 23166
rect 49758 23090 49810 23102
rect 50094 23154 50146 23166
rect 50094 23090 50146 23102
rect 50990 23154 51042 23166
rect 50990 23090 51042 23102
rect 51662 23154 51714 23166
rect 55246 23154 55298 23166
rect 53330 23102 53342 23154
rect 53394 23102 53406 23154
rect 54002 23102 54014 23154
rect 54066 23102 54078 23154
rect 51662 23090 51714 23102
rect 55246 23090 55298 23102
rect 56478 23154 56530 23166
rect 56478 23090 56530 23102
rect 18510 23042 18562 23054
rect 30046 23042 30098 23054
rect 24546 22990 24558 23042
rect 24610 22990 24622 23042
rect 26450 22990 26462 23042
rect 26514 22990 26526 23042
rect 18510 22978 18562 22990
rect 30046 22978 30098 22990
rect 31838 23042 31890 23054
rect 31838 22978 31890 22990
rect 32398 23042 32450 23054
rect 32398 22978 32450 22990
rect 32846 23042 32898 23054
rect 32846 22978 32898 22990
rect 33518 23042 33570 23054
rect 33518 22978 33570 22990
rect 34750 23042 34802 23054
rect 37886 23042 37938 23054
rect 35746 22990 35758 23042
rect 35810 22990 35822 23042
rect 34750 22978 34802 22990
rect 37886 22978 37938 22990
rect 38334 23042 38386 23054
rect 38334 22978 38386 22990
rect 40462 23042 40514 23054
rect 40462 22978 40514 22990
rect 41918 23042 41970 23054
rect 41918 22978 41970 22990
rect 43262 23042 43314 23054
rect 43262 22978 43314 22990
rect 43710 23042 43762 23054
rect 43710 22978 43762 22990
rect 44158 23042 44210 23054
rect 44158 22978 44210 22990
rect 45054 23042 45106 23054
rect 45054 22978 45106 22990
rect 45502 23042 45554 23054
rect 45502 22978 45554 22990
rect 46398 23042 46450 23054
rect 46398 22978 46450 22990
rect 48190 23042 48242 23054
rect 48190 22978 48242 22990
rect 49646 23042 49698 23054
rect 49646 22978 49698 22990
rect 50542 23042 50594 23054
rect 50542 22978 50594 22990
rect 51774 23042 51826 23054
rect 55134 23042 55186 23054
rect 53442 22990 53454 23042
rect 53506 22990 53518 23042
rect 51774 22978 51826 22990
rect 55134 22978 55186 22990
rect 56702 23042 56754 23054
rect 57922 22990 57934 23042
rect 57986 22990 57998 23042
rect 56702 22978 56754 22990
rect 28142 22930 28194 22942
rect 28142 22866 28194 22878
rect 36094 22930 36146 22942
rect 36306 22878 36318 22930
rect 36370 22927 36382 22930
rect 36642 22927 36654 22930
rect 36370 22881 36654 22927
rect 36370 22878 36382 22881
rect 36642 22878 36654 22881
rect 36706 22927 36718 22930
rect 37874 22927 37886 22930
rect 36706 22881 37886 22927
rect 36706 22878 36718 22881
rect 37874 22878 37886 22881
rect 37938 22927 37950 22930
rect 38434 22927 38446 22930
rect 37938 22881 38446 22927
rect 37938 22878 37950 22881
rect 38434 22878 38446 22881
rect 38498 22878 38510 22930
rect 47618 22878 47630 22930
rect 47682 22927 47694 22930
rect 48514 22927 48526 22930
rect 47682 22881 48526 22927
rect 47682 22878 47694 22881
rect 48514 22878 48526 22881
rect 48578 22878 48590 22930
rect 53330 22878 53342 22930
rect 53394 22878 53406 22930
rect 36094 22866 36146 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 26014 22594 26066 22606
rect 52558 22594 52610 22606
rect 32386 22542 32398 22594
rect 32450 22591 32462 22594
rect 33394 22591 33406 22594
rect 32450 22545 33406 22591
rect 32450 22542 32462 22545
rect 33394 22542 33406 22545
rect 33458 22542 33470 22594
rect 34962 22542 34974 22594
rect 35026 22591 35038 22594
rect 36082 22591 36094 22594
rect 35026 22545 36094 22591
rect 35026 22542 35038 22545
rect 36082 22542 36094 22545
rect 36146 22542 36158 22594
rect 42130 22542 42142 22594
rect 42194 22591 42206 22594
rect 43250 22591 43262 22594
rect 42194 22545 43262 22591
rect 42194 22542 42206 22545
rect 43250 22542 43262 22545
rect 43314 22542 43326 22594
rect 26014 22530 26066 22542
rect 52558 22530 52610 22542
rect 19742 22482 19794 22494
rect 19742 22418 19794 22430
rect 23774 22482 23826 22494
rect 23774 22418 23826 22430
rect 24782 22482 24834 22494
rect 24782 22418 24834 22430
rect 25118 22482 25170 22494
rect 25118 22418 25170 22430
rect 26238 22482 26290 22494
rect 26238 22418 26290 22430
rect 26798 22482 26850 22494
rect 26798 22418 26850 22430
rect 27470 22482 27522 22494
rect 27470 22418 27522 22430
rect 27582 22482 27634 22494
rect 27582 22418 27634 22430
rect 32174 22482 32226 22494
rect 32174 22418 32226 22430
rect 35198 22482 35250 22494
rect 35198 22418 35250 22430
rect 35758 22482 35810 22494
rect 35758 22418 35810 22430
rect 36094 22482 36146 22494
rect 36094 22418 36146 22430
rect 36542 22482 36594 22494
rect 40014 22482 40066 22494
rect 37986 22430 37998 22482
rect 38050 22430 38062 22482
rect 36542 22418 36594 22430
rect 40014 22418 40066 22430
rect 41806 22482 41858 22494
rect 41806 22418 41858 22430
rect 42142 22482 42194 22494
rect 42142 22418 42194 22430
rect 43598 22482 43650 22494
rect 43598 22418 43650 22430
rect 50430 22482 50482 22494
rect 50430 22418 50482 22430
rect 57038 22482 57090 22494
rect 57038 22418 57090 22430
rect 28926 22370 28978 22382
rect 33742 22370 33794 22382
rect 2818 22318 2830 22370
rect 2882 22318 2894 22370
rect 18946 22318 18958 22370
rect 19010 22318 19022 22370
rect 27234 22318 27246 22370
rect 27298 22318 27310 22370
rect 27682 22318 27694 22370
rect 27746 22367 27758 22370
rect 27906 22367 27918 22370
rect 27746 22321 27918 22367
rect 27746 22318 27758 22321
rect 27906 22318 27918 22321
rect 27970 22318 27982 22370
rect 29698 22318 29710 22370
rect 29762 22318 29774 22370
rect 28926 22306 28978 22318
rect 33742 22306 33794 22318
rect 37662 22370 37714 22382
rect 37662 22306 37714 22318
rect 39902 22370 39954 22382
rect 39902 22306 39954 22318
rect 40350 22370 40402 22382
rect 40350 22306 40402 22318
rect 42590 22370 42642 22382
rect 42590 22306 42642 22318
rect 44382 22370 44434 22382
rect 44382 22306 44434 22318
rect 46286 22370 46338 22382
rect 46286 22306 46338 22318
rect 47294 22370 47346 22382
rect 47294 22306 47346 22318
rect 47406 22370 47458 22382
rect 48414 22370 48466 22382
rect 47618 22318 47630 22370
rect 47682 22318 47694 22370
rect 47406 22306 47458 22318
rect 48414 22306 48466 22318
rect 48638 22370 48690 22382
rect 48638 22306 48690 22318
rect 53902 22370 53954 22382
rect 53902 22306 53954 22318
rect 54014 22370 54066 22382
rect 56814 22370 56866 22382
rect 54226 22318 54238 22370
rect 54290 22318 54302 22370
rect 54014 22306 54066 22318
rect 56814 22306 56866 22318
rect 57934 22370 57986 22382
rect 57934 22306 57986 22318
rect 18734 22258 18786 22270
rect 1922 22206 1934 22258
rect 1986 22206 1998 22258
rect 18734 22194 18786 22206
rect 22094 22258 22146 22270
rect 22094 22194 22146 22206
rect 22430 22258 22482 22270
rect 22430 22194 22482 22206
rect 23214 22258 23266 22270
rect 23214 22194 23266 22206
rect 23326 22258 23378 22270
rect 23326 22194 23378 22206
rect 28030 22258 28082 22270
rect 28030 22194 28082 22206
rect 31390 22258 31442 22270
rect 31390 22194 31442 22206
rect 31726 22258 31778 22270
rect 31726 22194 31778 22206
rect 34078 22258 34130 22270
rect 34078 22194 34130 22206
rect 34302 22258 34354 22270
rect 34302 22194 34354 22206
rect 39230 22258 39282 22270
rect 39230 22194 39282 22206
rect 40238 22258 40290 22270
rect 40238 22194 40290 22206
rect 40910 22258 40962 22270
rect 40910 22194 40962 22206
rect 41246 22258 41298 22270
rect 41246 22194 41298 22206
rect 45390 22258 45442 22270
rect 45390 22194 45442 22206
rect 48190 22258 48242 22270
rect 49086 22258 49138 22270
rect 48850 22206 48862 22258
rect 48914 22206 48926 22258
rect 48190 22194 48242 22206
rect 49086 22194 49138 22206
rect 52558 22258 52610 22270
rect 52558 22194 52610 22206
rect 52670 22258 52722 22270
rect 52670 22194 52722 22206
rect 54798 22258 54850 22270
rect 54798 22194 54850 22206
rect 57598 22258 57650 22270
rect 57598 22194 57650 22206
rect 22990 22146 23042 22158
rect 29934 22146 29986 22158
rect 25666 22094 25678 22146
rect 25730 22094 25742 22146
rect 22990 22082 23042 22094
rect 29934 22082 29986 22094
rect 30718 22146 30770 22158
rect 30718 22082 30770 22094
rect 32734 22146 32786 22158
rect 32734 22082 32786 22094
rect 33182 22146 33234 22158
rect 33182 22082 33234 22094
rect 33854 22146 33906 22158
rect 33854 22082 33906 22094
rect 34862 22146 34914 22158
rect 37998 22146 38050 22158
rect 37314 22094 37326 22146
rect 37378 22143 37390 22146
rect 37538 22143 37550 22146
rect 37378 22097 37550 22143
rect 37378 22094 37390 22097
rect 37538 22094 37550 22097
rect 37602 22094 37614 22146
rect 34862 22082 34914 22094
rect 37998 22082 38050 22094
rect 38222 22146 38274 22158
rect 38222 22082 38274 22094
rect 38670 22146 38722 22158
rect 38670 22082 38722 22094
rect 38782 22146 38834 22158
rect 38782 22082 38834 22094
rect 39006 22146 39058 22158
rect 39006 22082 39058 22094
rect 41134 22146 41186 22158
rect 41134 22082 41186 22094
rect 43038 22146 43090 22158
rect 43038 22082 43090 22094
rect 44046 22146 44098 22158
rect 44046 22082 44098 22094
rect 45950 22146 46002 22158
rect 45950 22082 46002 22094
rect 46174 22146 46226 22158
rect 48638 22146 48690 22158
rect 46834 22094 46846 22146
rect 46898 22094 46910 22146
rect 46174 22082 46226 22094
rect 48638 22082 48690 22094
rect 49534 22146 49586 22158
rect 49534 22082 49586 22094
rect 49982 22146 50034 22158
rect 49982 22082 50034 22094
rect 50878 22146 50930 22158
rect 50878 22082 50930 22094
rect 51326 22146 51378 22158
rect 51326 22082 51378 22094
rect 51774 22146 51826 22158
rect 55134 22146 55186 22158
rect 53442 22094 53454 22146
rect 53506 22094 53518 22146
rect 51774 22082 51826 22094
rect 55134 22082 55186 22094
rect 55582 22146 55634 22158
rect 56466 22094 56478 22146
rect 56530 22094 56542 22146
rect 55582 22082 55634 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 23550 21810 23602 21822
rect 23550 21746 23602 21758
rect 26126 21810 26178 21822
rect 26126 21746 26178 21758
rect 30718 21810 30770 21822
rect 30718 21746 30770 21758
rect 34078 21810 34130 21822
rect 34078 21746 34130 21758
rect 34638 21810 34690 21822
rect 34638 21746 34690 21758
rect 35982 21810 36034 21822
rect 35982 21746 36034 21758
rect 37326 21810 37378 21822
rect 37326 21746 37378 21758
rect 39454 21810 39506 21822
rect 39454 21746 39506 21758
rect 40238 21810 40290 21822
rect 40238 21746 40290 21758
rect 41694 21810 41746 21822
rect 41694 21746 41746 21758
rect 42142 21810 42194 21822
rect 42142 21746 42194 21758
rect 42702 21810 42754 21822
rect 42702 21746 42754 21758
rect 48190 21810 48242 21822
rect 48190 21746 48242 21758
rect 49646 21810 49698 21822
rect 49646 21746 49698 21758
rect 52894 21810 52946 21822
rect 52894 21746 52946 21758
rect 53678 21810 53730 21822
rect 53678 21746 53730 21758
rect 23326 21698 23378 21710
rect 23326 21634 23378 21646
rect 24782 21698 24834 21710
rect 24782 21634 24834 21646
rect 29150 21698 29202 21710
rect 29150 21634 29202 21646
rect 29486 21698 29538 21710
rect 29486 21634 29538 21646
rect 30606 21698 30658 21710
rect 30606 21634 30658 21646
rect 30942 21698 30994 21710
rect 30942 21634 30994 21646
rect 31950 21698 32002 21710
rect 31950 21634 32002 21646
rect 37102 21698 37154 21710
rect 37102 21634 37154 21646
rect 39342 21698 39394 21710
rect 39342 21634 39394 21646
rect 39566 21698 39618 21710
rect 39566 21634 39618 21646
rect 43486 21698 43538 21710
rect 45166 21698 45218 21710
rect 43486 21634 43538 21646
rect 43598 21642 43650 21654
rect 22654 21586 22706 21598
rect 22418 21534 22430 21586
rect 22482 21534 22494 21586
rect 22654 21522 22706 21534
rect 23998 21586 24050 21598
rect 32174 21586 32226 21598
rect 31378 21534 31390 21586
rect 31442 21534 31454 21586
rect 31714 21534 31726 21586
rect 31778 21534 31790 21586
rect 23998 21522 24050 21534
rect 32174 21522 32226 21534
rect 33742 21586 33794 21598
rect 33742 21522 33794 21534
rect 35422 21586 35474 21598
rect 35422 21522 35474 21534
rect 36990 21586 37042 21598
rect 36990 21522 37042 21534
rect 37998 21586 38050 21598
rect 37998 21522 38050 21534
rect 40462 21586 40514 21598
rect 40462 21522 40514 21534
rect 40910 21586 40962 21598
rect 40910 21522 40962 21534
rect 41918 21586 41970 21598
rect 45166 21634 45218 21646
rect 45390 21698 45442 21710
rect 50654 21698 50706 21710
rect 45938 21646 45950 21698
rect 46002 21646 46014 21698
rect 45390 21634 45442 21646
rect 50654 21634 50706 21646
rect 54798 21698 54850 21710
rect 54798 21634 54850 21646
rect 55022 21698 55074 21710
rect 55022 21634 55074 21646
rect 55918 21698 55970 21710
rect 55918 21634 55970 21646
rect 57822 21698 57874 21710
rect 57822 21634 57874 21646
rect 43598 21578 43650 21590
rect 44046 21586 44098 21598
rect 41918 21522 41970 21534
rect 44046 21522 44098 21534
rect 45054 21586 45106 21598
rect 48750 21586 48802 21598
rect 46274 21534 46286 21586
rect 46338 21534 46350 21586
rect 46946 21534 46958 21586
rect 47010 21534 47022 21586
rect 47954 21534 47966 21586
rect 48018 21534 48030 21586
rect 45054 21522 45106 21534
rect 48750 21522 48802 21534
rect 49534 21586 49586 21598
rect 49534 21522 49586 21534
rect 49758 21586 49810 21598
rect 49758 21522 49810 21534
rect 50094 21586 50146 21598
rect 50094 21522 50146 21534
rect 50990 21586 51042 21598
rect 50990 21522 51042 21534
rect 51886 21586 51938 21598
rect 51886 21522 51938 21534
rect 54126 21586 54178 21598
rect 54126 21522 54178 21534
rect 55470 21586 55522 21598
rect 55470 21522 55522 21534
rect 56030 21586 56082 21598
rect 57922 21534 57934 21586
rect 57986 21583 57998 21586
rect 58258 21583 58270 21586
rect 57986 21537 58270 21583
rect 57986 21534 57998 21537
rect 58258 21534 58270 21537
rect 58322 21534 58334 21586
rect 56030 21522 56082 21534
rect 21758 21474 21810 21486
rect 21758 21410 21810 21422
rect 23438 21474 23490 21486
rect 23438 21410 23490 21422
rect 24334 21474 24386 21486
rect 24334 21410 24386 21422
rect 28254 21474 28306 21486
rect 28254 21410 28306 21422
rect 28702 21474 28754 21486
rect 28702 21410 28754 21422
rect 30046 21474 30098 21486
rect 32622 21474 32674 21486
rect 31938 21422 31950 21474
rect 32002 21422 32014 21474
rect 30046 21410 30098 21422
rect 32622 21410 32674 21422
rect 34078 21474 34130 21486
rect 34078 21410 34130 21422
rect 36430 21474 36482 21486
rect 36430 21410 36482 21422
rect 37774 21474 37826 21486
rect 37774 21410 37826 21422
rect 38782 21474 38834 21486
rect 38782 21410 38834 21422
rect 40350 21474 40402 21486
rect 40350 21410 40402 21422
rect 41806 21474 41858 21486
rect 41806 21410 41858 21422
rect 44494 21474 44546 21486
rect 44494 21410 44546 21422
rect 46510 21474 46562 21486
rect 51438 21474 51490 21486
rect 46722 21422 46734 21474
rect 46786 21422 46798 21474
rect 46510 21410 46562 21422
rect 51438 21410 51490 21422
rect 52334 21474 52386 21486
rect 52334 21410 52386 21422
rect 53230 21474 53282 21486
rect 53230 21410 53282 21422
rect 54910 21474 54962 21486
rect 54910 21410 54962 21422
rect 55694 21474 55746 21486
rect 55694 21410 55746 21422
rect 56590 21474 56642 21486
rect 57474 21422 57486 21474
rect 57538 21422 57550 21474
rect 56590 21410 56642 21422
rect 33966 21362 34018 21374
rect 24322 21310 24334 21362
rect 24386 21359 24398 21362
rect 24658 21359 24670 21362
rect 24386 21313 24670 21359
rect 24386 21310 24398 21313
rect 24658 21310 24670 21313
rect 24722 21359 24734 21362
rect 25106 21359 25118 21362
rect 24722 21313 25118 21359
rect 24722 21310 24734 21313
rect 25106 21310 25118 21313
rect 25170 21310 25182 21362
rect 33966 21298 34018 21310
rect 35534 21362 35586 21374
rect 43486 21362 43538 21374
rect 35746 21310 35758 21362
rect 35810 21359 35822 21362
rect 36754 21359 36766 21362
rect 35810 21313 36766 21359
rect 35810 21310 35822 21313
rect 36754 21310 36766 21313
rect 36818 21310 36830 21362
rect 38322 21310 38334 21362
rect 38386 21310 38398 21362
rect 35534 21298 35586 21310
rect 43486 21298 43538 21310
rect 48302 21362 48354 21374
rect 52322 21310 52334 21362
rect 52386 21359 52398 21362
rect 52882 21359 52894 21362
rect 52386 21313 52894 21359
rect 52386 21310 52398 21313
rect 52882 21310 52894 21313
rect 52946 21310 52958 21362
rect 48302 21298 48354 21310
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 34862 21026 34914 21038
rect 49534 21026 49586 21038
rect 33282 20974 33294 21026
rect 33346 21023 33358 21026
rect 33506 21023 33518 21026
rect 33346 20977 33518 21023
rect 33346 20974 33358 20977
rect 33506 20974 33518 20977
rect 33570 20974 33582 21026
rect 39330 20974 39342 21026
rect 39394 21023 39406 21026
rect 40226 21023 40238 21026
rect 39394 20977 40238 21023
rect 39394 20974 39406 20977
rect 40226 20974 40238 20977
rect 40290 20974 40302 21026
rect 34862 20962 34914 20974
rect 49534 20962 49586 20974
rect 50542 21026 50594 21038
rect 51426 20974 51438 21026
rect 51490 21023 51502 21026
rect 51986 21023 51998 21026
rect 51490 20977 51998 21023
rect 51490 20974 51502 20977
rect 51986 20974 51998 20977
rect 52050 20974 52062 21026
rect 52322 20974 52334 21026
rect 52386 21023 52398 21026
rect 52770 21023 52782 21026
rect 52386 20977 52782 21023
rect 52386 20974 52398 20977
rect 52770 20974 52782 20977
rect 52834 20974 52846 21026
rect 50542 20962 50594 20974
rect 21758 20914 21810 20926
rect 31054 20914 31106 20926
rect 22194 20862 22206 20914
rect 22258 20862 22270 20914
rect 21758 20850 21810 20862
rect 31054 20850 31106 20862
rect 31278 20914 31330 20926
rect 31278 20850 31330 20862
rect 32622 20914 32674 20926
rect 32622 20850 32674 20862
rect 33182 20914 33234 20926
rect 33182 20850 33234 20862
rect 33518 20914 33570 20926
rect 33518 20850 33570 20862
rect 36766 20914 36818 20926
rect 36766 20850 36818 20862
rect 38446 20914 38498 20926
rect 38446 20850 38498 20862
rect 39454 20914 39506 20926
rect 39454 20850 39506 20862
rect 40238 20914 40290 20926
rect 40238 20850 40290 20862
rect 44718 20914 44770 20926
rect 44718 20850 44770 20862
rect 45390 20914 45442 20926
rect 45390 20850 45442 20862
rect 51438 20914 51490 20926
rect 51438 20850 51490 20862
rect 52222 20914 52274 20926
rect 52222 20850 52274 20862
rect 54686 20914 54738 20926
rect 54686 20850 54738 20862
rect 23774 20802 23826 20814
rect 22530 20750 22542 20802
rect 22594 20750 22606 20802
rect 23774 20738 23826 20750
rect 25902 20802 25954 20814
rect 28478 20802 28530 20814
rect 32174 20802 32226 20814
rect 26674 20750 26686 20802
rect 26738 20750 26750 20802
rect 29922 20750 29934 20802
rect 29986 20750 29998 20802
rect 30706 20750 30718 20802
rect 30770 20750 30782 20802
rect 25902 20738 25954 20750
rect 28478 20738 28530 20750
rect 32174 20738 32226 20750
rect 34414 20802 34466 20814
rect 34414 20738 34466 20750
rect 34750 20802 34802 20814
rect 34750 20738 34802 20750
rect 34974 20802 35026 20814
rect 34974 20738 35026 20750
rect 38110 20802 38162 20814
rect 38110 20738 38162 20750
rect 38222 20802 38274 20814
rect 38222 20738 38274 20750
rect 38670 20802 38722 20814
rect 38670 20738 38722 20750
rect 38894 20802 38946 20814
rect 38894 20738 38946 20750
rect 40910 20802 40962 20814
rect 40910 20738 40962 20750
rect 41246 20802 41298 20814
rect 41246 20738 41298 20750
rect 41470 20802 41522 20814
rect 41470 20738 41522 20750
rect 42366 20802 42418 20814
rect 42366 20738 42418 20750
rect 42590 20802 42642 20814
rect 46286 20802 46338 20814
rect 43810 20750 43822 20802
rect 43874 20750 43886 20802
rect 42590 20738 42642 20750
rect 46286 20738 46338 20750
rect 46734 20802 46786 20814
rect 47966 20802 48018 20814
rect 47058 20750 47070 20802
rect 47122 20750 47134 20802
rect 46734 20738 46786 20750
rect 47966 20738 48018 20750
rect 49422 20802 49474 20814
rect 53790 20802 53842 20814
rect 54126 20802 54178 20814
rect 50866 20750 50878 20802
rect 50930 20750 50942 20802
rect 53442 20750 53454 20802
rect 53506 20750 53518 20802
rect 54002 20750 54014 20802
rect 54066 20750 54078 20802
rect 49422 20738 49474 20750
rect 53790 20738 53842 20750
rect 54126 20738 54178 20750
rect 54238 20802 54290 20814
rect 55682 20750 55694 20802
rect 55746 20750 55758 20802
rect 57250 20750 57262 20802
rect 57314 20750 57326 20802
rect 54238 20738 54290 20750
rect 2382 20690 2434 20702
rect 2382 20626 2434 20638
rect 2718 20690 2770 20702
rect 2718 20626 2770 20638
rect 24110 20690 24162 20702
rect 24110 20626 24162 20638
rect 24670 20690 24722 20702
rect 24670 20626 24722 20638
rect 25006 20690 25058 20702
rect 25006 20626 25058 20638
rect 25566 20690 25618 20702
rect 25566 20626 25618 20638
rect 27134 20690 27186 20702
rect 27134 20626 27186 20638
rect 28030 20690 28082 20702
rect 28030 20626 28082 20638
rect 28702 20690 28754 20702
rect 28702 20626 28754 20638
rect 35982 20690 36034 20702
rect 35982 20626 36034 20638
rect 36094 20690 36146 20702
rect 36094 20626 36146 20638
rect 36206 20690 36258 20702
rect 44046 20690 44098 20702
rect 48638 20690 48690 20702
rect 50094 20690 50146 20702
rect 43698 20638 43710 20690
rect 43762 20638 43774 20690
rect 46498 20638 46510 20690
rect 46562 20638 46574 20690
rect 48850 20638 48862 20690
rect 48914 20638 48926 20690
rect 50306 20638 50318 20690
rect 50370 20638 50382 20690
rect 57698 20638 57710 20690
rect 57762 20638 57774 20690
rect 36206 20626 36258 20638
rect 44046 20626 44098 20638
rect 48638 20626 48690 20638
rect 50094 20626 50146 20638
rect 3278 20578 3330 20590
rect 3278 20514 3330 20526
rect 23438 20578 23490 20590
rect 23438 20514 23490 20526
rect 23998 20578 24050 20590
rect 23998 20514 24050 20526
rect 27246 20578 27298 20590
rect 27246 20514 27298 20526
rect 27358 20578 27410 20590
rect 27358 20514 27410 20526
rect 27470 20578 27522 20590
rect 27470 20514 27522 20526
rect 27918 20578 27970 20590
rect 27918 20514 27970 20526
rect 28254 20578 28306 20590
rect 28254 20514 28306 20526
rect 30158 20578 30210 20590
rect 34526 20578 34578 20590
rect 37998 20578 38050 20590
rect 31826 20526 31838 20578
rect 31890 20526 31902 20578
rect 35522 20526 35534 20578
rect 35586 20526 35598 20578
rect 30158 20514 30210 20526
rect 34526 20514 34578 20526
rect 37998 20514 38050 20526
rect 39790 20578 39842 20590
rect 39790 20514 39842 20526
rect 41246 20578 41298 20590
rect 41246 20514 41298 20526
rect 42478 20578 42530 20590
rect 42478 20514 42530 20526
rect 42814 20578 42866 20590
rect 42814 20514 42866 20526
rect 44158 20578 44210 20590
rect 44158 20514 44210 20526
rect 44270 20578 44322 20590
rect 48750 20578 48802 20590
rect 46722 20526 46734 20578
rect 46786 20526 46798 20578
rect 47618 20526 47630 20578
rect 47682 20526 47694 20578
rect 44270 20514 44322 20526
rect 48750 20514 48802 20526
rect 49086 20578 49138 20590
rect 49086 20514 49138 20526
rect 50878 20578 50930 20590
rect 50878 20514 50930 20526
rect 51774 20578 51826 20590
rect 51774 20514 51826 20526
rect 52670 20578 52722 20590
rect 52670 20514 52722 20526
rect 55582 20578 55634 20590
rect 55582 20514 55634 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 23102 20242 23154 20254
rect 23102 20178 23154 20190
rect 24782 20242 24834 20254
rect 24782 20178 24834 20190
rect 26462 20242 26514 20254
rect 30606 20242 30658 20254
rect 29026 20190 29038 20242
rect 29090 20190 29102 20242
rect 26462 20178 26514 20190
rect 30606 20178 30658 20190
rect 31838 20242 31890 20254
rect 37326 20242 37378 20254
rect 33954 20190 33966 20242
rect 34018 20190 34030 20242
rect 31838 20178 31890 20190
rect 37326 20178 37378 20190
rect 38222 20242 38274 20254
rect 38222 20178 38274 20190
rect 42926 20242 42978 20254
rect 42926 20178 42978 20190
rect 43934 20242 43986 20254
rect 43934 20178 43986 20190
rect 44158 20242 44210 20254
rect 52334 20242 52386 20254
rect 56366 20242 56418 20254
rect 45490 20190 45502 20242
rect 45554 20190 45566 20242
rect 53330 20190 53342 20242
rect 53394 20190 53406 20242
rect 44158 20178 44210 20190
rect 52334 20178 52386 20190
rect 56366 20178 56418 20190
rect 57486 20242 57538 20254
rect 57486 20178 57538 20190
rect 24334 20130 24386 20142
rect 24334 20066 24386 20078
rect 25566 20130 25618 20142
rect 25566 20066 25618 20078
rect 28142 20130 28194 20142
rect 28142 20066 28194 20078
rect 28366 20130 28418 20142
rect 28366 20066 28418 20078
rect 29934 20130 29986 20142
rect 29934 20066 29986 20078
rect 31054 20130 31106 20142
rect 31054 20066 31106 20078
rect 34862 20130 34914 20142
rect 34862 20066 34914 20078
rect 35422 20130 35474 20142
rect 35422 20066 35474 20078
rect 35870 20130 35922 20142
rect 35870 20066 35922 20078
rect 36878 20130 36930 20142
rect 36878 20066 36930 20078
rect 36990 20130 37042 20142
rect 36990 20066 37042 20078
rect 39006 20130 39058 20142
rect 39006 20066 39058 20078
rect 39454 20130 39506 20142
rect 39454 20066 39506 20078
rect 40350 20130 40402 20142
rect 40350 20066 40402 20078
rect 40798 20130 40850 20142
rect 40798 20066 40850 20078
rect 42030 20130 42082 20142
rect 50766 20130 50818 20142
rect 45378 20078 45390 20130
rect 45442 20078 45454 20130
rect 42030 20066 42082 20078
rect 50766 20066 50818 20078
rect 50878 20130 50930 20142
rect 50878 20066 50930 20078
rect 52110 20130 52162 20142
rect 52110 20066 52162 20078
rect 26686 20018 26738 20030
rect 26686 19954 26738 19966
rect 27134 20018 27186 20030
rect 27134 19954 27186 19966
rect 28478 20018 28530 20030
rect 28478 19954 28530 19966
rect 29374 20018 29426 20030
rect 29374 19954 29426 19966
rect 30718 20018 30770 20030
rect 30718 19954 30770 19966
rect 30830 20018 30882 20030
rect 30830 19954 30882 19966
rect 34302 20018 34354 20030
rect 34302 19954 34354 19966
rect 35086 20018 35138 20030
rect 35086 19954 35138 19966
rect 37102 20018 37154 20030
rect 38558 20018 38610 20030
rect 42366 20018 42418 20030
rect 50542 20018 50594 20030
rect 51886 20018 51938 20030
rect 38210 19966 38222 20018
rect 38274 19966 38286 20018
rect 38770 19966 38782 20018
rect 38834 19966 38846 20018
rect 43138 19966 43150 20018
rect 43202 19966 43214 20018
rect 44370 19966 44382 20018
rect 44434 19966 44446 20018
rect 45490 19966 45502 20018
rect 45554 19966 45566 20018
rect 48178 19966 48190 20018
rect 48242 19966 48254 20018
rect 48626 19966 48638 20018
rect 48690 19966 48702 20018
rect 51202 19966 51214 20018
rect 51266 19966 51278 20018
rect 37102 19954 37154 19966
rect 38558 19954 38610 19966
rect 42366 19954 42418 19966
rect 50542 19954 50594 19966
rect 51886 19954 51938 19966
rect 53006 20018 53058 20030
rect 53006 19954 53058 19966
rect 53790 20018 53842 20030
rect 54786 19966 54798 20018
rect 54850 19966 54862 20018
rect 55234 19966 55246 20018
rect 55298 19966 55310 20018
rect 57698 19966 57710 20018
rect 57762 19966 57774 20018
rect 53790 19954 53842 19966
rect 22430 19906 22482 19918
rect 22430 19842 22482 19854
rect 23550 19906 23602 19918
rect 23550 19842 23602 19854
rect 26574 19906 26626 19918
rect 26574 19842 26626 19854
rect 27694 19906 27746 19918
rect 27694 19842 27746 19854
rect 32510 19906 32562 19918
rect 32510 19842 32562 19854
rect 34974 19906 35026 19918
rect 34974 19842 35026 19854
rect 36318 19906 36370 19918
rect 36318 19842 36370 19854
rect 39902 19906 39954 19918
rect 39902 19842 39954 19854
rect 41470 19906 41522 19918
rect 41470 19842 41522 19854
rect 43822 19906 43874 19918
rect 43822 19842 43874 19854
rect 49422 19906 49474 19918
rect 49422 19842 49474 19854
rect 49870 19906 49922 19918
rect 51998 19906 52050 19918
rect 51314 19854 51326 19906
rect 51378 19854 51390 19906
rect 55346 19854 55358 19906
rect 55410 19854 55422 19906
rect 49870 19842 49922 19854
rect 51998 19842 52050 19854
rect 24222 19794 24274 19806
rect 24222 19730 24274 19742
rect 31726 19794 31778 19806
rect 31726 19730 31778 19742
rect 32062 19794 32114 19806
rect 55570 19742 55582 19794
rect 55634 19742 55646 19794
rect 32062 19730 32114 19742
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 25902 19458 25954 19470
rect 31614 19458 31666 19470
rect 30818 19406 30830 19458
rect 30882 19455 30894 19458
rect 31154 19455 31166 19458
rect 30882 19409 31166 19455
rect 30882 19406 30894 19409
rect 31154 19406 31166 19409
rect 31218 19406 31230 19458
rect 25902 19394 25954 19406
rect 31614 19394 31666 19406
rect 44270 19458 44322 19470
rect 51102 19458 51154 19470
rect 46946 19406 46958 19458
rect 47010 19455 47022 19458
rect 47618 19455 47630 19458
rect 47010 19409 47630 19455
rect 47010 19406 47022 19409
rect 47618 19406 47630 19409
rect 47682 19406 47694 19458
rect 44270 19394 44322 19406
rect 51102 19394 51154 19406
rect 26126 19346 26178 19358
rect 26126 19282 26178 19294
rect 26574 19346 26626 19358
rect 26574 19282 26626 19294
rect 32398 19346 32450 19358
rect 32398 19282 32450 19294
rect 32846 19346 32898 19358
rect 32846 19282 32898 19294
rect 36206 19346 36258 19358
rect 36206 19282 36258 19294
rect 36542 19346 36594 19358
rect 36542 19282 36594 19294
rect 39566 19346 39618 19358
rect 39566 19282 39618 19294
rect 42030 19346 42082 19358
rect 42030 19282 42082 19294
rect 46286 19346 46338 19358
rect 46286 19282 46338 19294
rect 46734 19346 46786 19358
rect 46734 19282 46786 19294
rect 47182 19346 47234 19358
rect 47182 19282 47234 19294
rect 47630 19346 47682 19358
rect 47630 19282 47682 19294
rect 48078 19346 48130 19358
rect 48078 19282 48130 19294
rect 48526 19346 48578 19358
rect 48526 19282 48578 19294
rect 48974 19346 49026 19358
rect 48974 19282 49026 19294
rect 49422 19346 49474 19358
rect 49422 19282 49474 19294
rect 49870 19346 49922 19358
rect 49870 19282 49922 19294
rect 53342 19346 53394 19358
rect 53342 19282 53394 19294
rect 24110 19234 24162 19246
rect 33630 19234 33682 19246
rect 24434 19182 24446 19234
rect 24498 19182 24510 19234
rect 24110 19170 24162 19182
rect 33630 19170 33682 19182
rect 34526 19234 34578 19246
rect 34526 19170 34578 19182
rect 34862 19234 34914 19246
rect 34862 19170 34914 19182
rect 35310 19234 35362 19246
rect 35310 19170 35362 19182
rect 38334 19234 38386 19246
rect 38334 19170 38386 19182
rect 43150 19234 43202 19246
rect 43150 19170 43202 19182
rect 44382 19234 44434 19246
rect 44382 19170 44434 19182
rect 50542 19234 50594 19246
rect 50542 19170 50594 19182
rect 50990 19234 51042 19246
rect 50990 19170 51042 19182
rect 51326 19234 51378 19246
rect 51326 19170 51378 19182
rect 55470 19234 55522 19246
rect 55470 19170 55522 19182
rect 56254 19234 56306 19246
rect 57138 19182 57150 19234
rect 57202 19182 57214 19234
rect 56254 19170 56306 19182
rect 21646 19122 21698 19134
rect 21646 19058 21698 19070
rect 21870 19122 21922 19134
rect 21870 19058 21922 19070
rect 22206 19122 22258 19134
rect 22206 19058 22258 19070
rect 25006 19122 25058 19134
rect 25006 19058 25058 19070
rect 30830 19122 30882 19134
rect 30830 19058 30882 19070
rect 31390 19122 31442 19134
rect 31390 19058 31442 19070
rect 33518 19122 33570 19134
rect 33518 19058 33570 19070
rect 34750 19122 34802 19134
rect 34750 19058 34802 19070
rect 35646 19122 35698 19134
rect 35646 19058 35698 19070
rect 39118 19122 39170 19134
rect 39118 19058 39170 19070
rect 40014 19122 40066 19134
rect 40014 19058 40066 19070
rect 45950 19122 46002 19134
rect 45950 19058 46002 19070
rect 51550 19122 51602 19134
rect 51550 19058 51602 19070
rect 54350 19122 54402 19134
rect 54350 19058 54402 19070
rect 55022 19122 55074 19134
rect 55022 19058 55074 19070
rect 55246 19122 55298 19134
rect 55246 19058 55298 19070
rect 58046 19122 58098 19134
rect 58046 19058 58098 19070
rect 22094 19010 22146 19022
rect 22094 18946 22146 18958
rect 22654 19010 22706 19022
rect 22654 18946 22706 18958
rect 23550 19010 23602 19022
rect 27246 19010 27298 19022
rect 25554 18958 25566 19010
rect 25618 18958 25630 19010
rect 23550 18946 23602 18958
rect 27246 18946 27298 18958
rect 28702 19010 28754 19022
rect 28702 18946 28754 18958
rect 29598 19010 29650 19022
rect 33294 19010 33346 19022
rect 31938 18958 31950 19010
rect 32002 18958 32014 19010
rect 29598 18946 29650 18958
rect 33294 18946 33346 18958
rect 34190 19010 34242 19022
rect 34190 18946 34242 18958
rect 35534 19010 35586 19022
rect 35534 18946 35586 18958
rect 37550 19010 37602 19022
rect 37550 18946 37602 18958
rect 37998 19010 38050 19022
rect 37998 18946 38050 18958
rect 38222 19010 38274 19022
rect 38222 18946 38274 18958
rect 38782 19010 38834 19022
rect 38782 18946 38834 18958
rect 39006 19010 39058 19022
rect 39006 18946 39058 18958
rect 40798 19010 40850 19022
rect 41582 19010 41634 19022
rect 43598 19010 43650 19022
rect 41122 18958 41134 19010
rect 41186 18958 41198 19010
rect 42802 18958 42814 19010
rect 42866 18958 42878 19010
rect 40798 18946 40850 18958
rect 41582 18946 41634 18958
rect 43598 18946 43650 18958
rect 44270 19010 44322 19022
rect 44270 18946 44322 18958
rect 45390 19010 45442 19022
rect 45390 18946 45442 18958
rect 51662 19010 51714 19022
rect 51662 18946 51714 18958
rect 51998 19010 52050 19022
rect 51998 18946 52050 18958
rect 52446 19010 52498 19022
rect 52446 18946 52498 18958
rect 54014 19010 54066 19022
rect 54014 18946 54066 18958
rect 55358 19010 55410 19022
rect 55358 18946 55410 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 24222 18674 24274 18686
rect 24222 18610 24274 18622
rect 24894 18674 24946 18686
rect 24894 18610 24946 18622
rect 27582 18674 27634 18686
rect 27582 18610 27634 18622
rect 28030 18674 28082 18686
rect 28030 18610 28082 18622
rect 31390 18674 31442 18686
rect 31390 18610 31442 18622
rect 33518 18674 33570 18686
rect 33518 18610 33570 18622
rect 37886 18674 37938 18686
rect 37886 18610 37938 18622
rect 39006 18674 39058 18686
rect 39006 18610 39058 18622
rect 39342 18674 39394 18686
rect 39342 18610 39394 18622
rect 40126 18674 40178 18686
rect 40126 18610 40178 18622
rect 42814 18674 42866 18686
rect 42814 18610 42866 18622
rect 43934 18674 43986 18686
rect 43934 18610 43986 18622
rect 44158 18674 44210 18686
rect 44158 18610 44210 18622
rect 47294 18674 47346 18686
rect 47294 18610 47346 18622
rect 48190 18674 48242 18686
rect 48190 18610 48242 18622
rect 48414 18674 48466 18686
rect 48414 18610 48466 18622
rect 16942 18562 16994 18574
rect 16942 18498 16994 18510
rect 23214 18562 23266 18574
rect 23214 18498 23266 18510
rect 23550 18562 23602 18574
rect 23550 18498 23602 18510
rect 24446 18562 24498 18574
rect 24446 18498 24498 18510
rect 25790 18562 25842 18574
rect 25790 18498 25842 18510
rect 25902 18562 25954 18574
rect 25902 18498 25954 18510
rect 26462 18562 26514 18574
rect 26462 18498 26514 18510
rect 27694 18562 27746 18574
rect 27694 18498 27746 18510
rect 31614 18562 31666 18574
rect 31614 18498 31666 18510
rect 35310 18562 35362 18574
rect 35310 18498 35362 18510
rect 35982 18562 36034 18574
rect 35982 18498 36034 18510
rect 36094 18562 36146 18574
rect 36094 18498 36146 18510
rect 38782 18562 38834 18574
rect 38782 18498 38834 18510
rect 40238 18562 40290 18574
rect 40238 18498 40290 18510
rect 42366 18562 42418 18574
rect 42366 18498 42418 18510
rect 44046 18562 44098 18574
rect 44046 18498 44098 18510
rect 44382 18562 44434 18574
rect 44382 18498 44434 18510
rect 46622 18562 46674 18574
rect 46622 18498 46674 18510
rect 47630 18562 47682 18574
rect 47630 18498 47682 18510
rect 48302 18562 48354 18574
rect 57486 18562 57538 18574
rect 51650 18510 51662 18562
rect 51714 18510 51726 18562
rect 53442 18510 53454 18562
rect 53506 18510 53518 18562
rect 54338 18510 54350 18562
rect 54402 18510 54414 18562
rect 56242 18510 56254 18562
rect 56306 18510 56318 18562
rect 48302 18498 48354 18510
rect 57486 18498 57538 18510
rect 57822 18562 57874 18574
rect 57822 18498 57874 18510
rect 18174 18450 18226 18462
rect 19630 18450 19682 18462
rect 21198 18450 21250 18462
rect 22094 18450 22146 18462
rect 16482 18398 16494 18450
rect 16546 18398 16558 18450
rect 18946 18398 18958 18450
rect 19010 18398 19022 18450
rect 20178 18398 20190 18450
rect 20242 18398 20254 18450
rect 21634 18398 21646 18450
rect 21698 18398 21710 18450
rect 18174 18386 18226 18398
rect 19630 18386 19682 18398
rect 21198 18386 21250 18398
rect 22094 18386 22146 18398
rect 26798 18450 26850 18462
rect 26798 18386 26850 18398
rect 27022 18450 27074 18462
rect 27022 18386 27074 18398
rect 27806 18450 27858 18462
rect 27806 18386 27858 18398
rect 29262 18450 29314 18462
rect 29262 18386 29314 18398
rect 29822 18450 29874 18462
rect 29822 18386 29874 18398
rect 30718 18450 30770 18462
rect 30718 18386 30770 18398
rect 32062 18450 32114 18462
rect 32062 18386 32114 18398
rect 34974 18450 35026 18462
rect 34974 18386 35026 18398
rect 35758 18450 35810 18462
rect 35758 18386 35810 18398
rect 36542 18450 36594 18462
rect 36542 18386 36594 18398
rect 36990 18450 37042 18462
rect 36990 18386 37042 18398
rect 39230 18450 39282 18462
rect 39230 18386 39282 18398
rect 40798 18450 40850 18462
rect 40798 18386 40850 18398
rect 41918 18450 41970 18462
rect 41918 18386 41970 18398
rect 42030 18450 42082 18462
rect 42030 18386 42082 18398
rect 43822 18450 43874 18462
rect 43822 18386 43874 18398
rect 44942 18450 44994 18462
rect 44942 18386 44994 18398
rect 46734 18450 46786 18462
rect 46734 18386 46786 18398
rect 48862 18450 48914 18462
rect 48862 18386 48914 18398
rect 49646 18450 49698 18462
rect 53902 18450 53954 18462
rect 49970 18398 49982 18450
rect 50034 18398 50046 18450
rect 50754 18398 50766 18450
rect 50818 18398 50830 18450
rect 51314 18398 51326 18450
rect 51378 18398 51390 18450
rect 52770 18398 52782 18450
rect 52834 18398 52846 18450
rect 53666 18398 53678 18450
rect 53730 18398 53742 18450
rect 54450 18398 54462 18450
rect 54514 18398 54526 18450
rect 55122 18398 55134 18450
rect 55186 18398 55198 18450
rect 55682 18398 55694 18450
rect 55746 18398 55758 18450
rect 56466 18398 56478 18450
rect 56530 18398 56542 18450
rect 49646 18386 49698 18398
rect 53902 18386 53954 18398
rect 22766 18338 22818 18350
rect 26910 18338 26962 18350
rect 16706 18286 16718 18338
rect 16770 18286 16782 18338
rect 24098 18286 24110 18338
rect 24162 18286 24174 18338
rect 22766 18274 22818 18286
rect 26910 18274 26962 18286
rect 28814 18338 28866 18350
rect 28814 18274 28866 18286
rect 30382 18338 30434 18350
rect 30382 18274 30434 18286
rect 31502 18338 31554 18350
rect 31502 18274 31554 18286
rect 32398 18338 32450 18350
rect 32398 18274 32450 18286
rect 32846 18338 32898 18350
rect 32846 18274 32898 18286
rect 33966 18338 34018 18350
rect 37438 18338 37490 18350
rect 34738 18286 34750 18338
rect 34802 18286 34814 18338
rect 33966 18274 34018 18286
rect 37438 18274 37490 18286
rect 39118 18338 39170 18350
rect 39118 18274 39170 18286
rect 42254 18338 42306 18350
rect 42254 18274 42306 18286
rect 45726 18338 45778 18350
rect 45726 18274 45778 18286
rect 56030 18338 56082 18350
rect 56030 18274 56082 18286
rect 25790 18226 25842 18238
rect 40014 18226 40066 18238
rect 29810 18174 29822 18226
rect 29874 18223 29886 18226
rect 30706 18223 30718 18226
rect 29874 18177 30718 18223
rect 29874 18174 29886 18177
rect 30706 18174 30718 18177
rect 30770 18174 30782 18226
rect 32162 18174 32174 18226
rect 32226 18223 32238 18226
rect 32834 18223 32846 18226
rect 32226 18177 32846 18223
rect 32226 18174 32238 18177
rect 32834 18174 32846 18177
rect 32898 18174 32910 18226
rect 25790 18162 25842 18174
rect 40014 18162 40066 18174
rect 45838 18226 45890 18238
rect 45838 18162 45890 18174
rect 46622 18226 46674 18238
rect 49746 18174 49758 18226
rect 49810 18174 49822 18226
rect 46622 18162 46674 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 16606 17890 16658 17902
rect 16606 17826 16658 17838
rect 17502 17890 17554 17902
rect 30606 17890 30658 17902
rect 20850 17838 20862 17890
rect 20914 17838 20926 17890
rect 17502 17826 17554 17838
rect 30606 17826 30658 17838
rect 30830 17890 30882 17902
rect 30830 17826 30882 17838
rect 39006 17890 39058 17902
rect 39006 17826 39058 17838
rect 39902 17890 39954 17902
rect 39902 17826 39954 17838
rect 44382 17890 44434 17902
rect 44382 17826 44434 17838
rect 50990 17890 51042 17902
rect 50990 17826 51042 17838
rect 51326 17890 51378 17902
rect 51326 17826 51378 17838
rect 19854 17778 19906 17790
rect 15138 17726 15150 17778
rect 15202 17726 15214 17778
rect 16258 17726 16270 17778
rect 16322 17726 16334 17778
rect 19854 17714 19906 17726
rect 20526 17778 20578 17790
rect 20526 17714 20578 17726
rect 26126 17778 26178 17790
rect 48302 17778 48354 17790
rect 57934 17778 57986 17790
rect 28018 17726 28030 17778
rect 28082 17726 28094 17778
rect 55906 17726 55918 17778
rect 55970 17726 55982 17778
rect 26126 17714 26178 17726
rect 48302 17714 48354 17726
rect 57934 17714 57986 17726
rect 14366 17666 14418 17678
rect 16830 17666 16882 17678
rect 2818 17614 2830 17666
rect 2882 17614 2894 17666
rect 15250 17614 15262 17666
rect 15314 17614 15326 17666
rect 14366 17602 14418 17614
rect 16830 17602 16882 17614
rect 20302 17666 20354 17678
rect 23886 17666 23938 17678
rect 22642 17614 22654 17666
rect 22706 17614 22718 17666
rect 23202 17614 23214 17666
rect 23266 17614 23278 17666
rect 20302 17602 20354 17614
rect 23886 17602 23938 17614
rect 24110 17666 24162 17678
rect 24110 17602 24162 17614
rect 24558 17666 24610 17678
rect 24558 17602 24610 17614
rect 24894 17666 24946 17678
rect 29822 17666 29874 17678
rect 27234 17614 27246 17666
rect 27298 17614 27310 17666
rect 24894 17602 24946 17614
rect 29822 17602 29874 17614
rect 32398 17666 32450 17678
rect 33518 17666 33570 17678
rect 32610 17614 32622 17666
rect 32674 17614 32686 17666
rect 32398 17602 32450 17614
rect 33518 17602 33570 17614
rect 33854 17666 33906 17678
rect 33854 17602 33906 17614
rect 34414 17666 34466 17678
rect 34414 17602 34466 17614
rect 35086 17666 35138 17678
rect 35086 17602 35138 17614
rect 35310 17666 35362 17678
rect 35310 17602 35362 17614
rect 36206 17666 36258 17678
rect 36878 17666 36930 17678
rect 36530 17614 36542 17666
rect 36594 17614 36606 17666
rect 36206 17602 36258 17614
rect 36878 17602 36930 17614
rect 38894 17666 38946 17678
rect 51214 17666 51266 17678
rect 53454 17666 53506 17678
rect 39218 17614 39230 17666
rect 39282 17614 39294 17666
rect 40226 17614 40238 17666
rect 40290 17614 40302 17666
rect 41234 17614 41246 17666
rect 41298 17614 41310 17666
rect 42130 17614 42142 17666
rect 42194 17614 42206 17666
rect 42690 17614 42702 17666
rect 42754 17614 42766 17666
rect 44146 17614 44158 17666
rect 44210 17614 44222 17666
rect 44706 17614 44718 17666
rect 44770 17614 44782 17666
rect 46050 17614 46062 17666
rect 46114 17614 46126 17666
rect 47394 17614 47406 17666
rect 47458 17614 47470 17666
rect 49634 17614 49646 17666
rect 49698 17614 49710 17666
rect 52546 17614 52558 17666
rect 52610 17614 52622 17666
rect 54898 17614 54910 17666
rect 54962 17614 54974 17666
rect 56802 17614 56814 17666
rect 56866 17614 56878 17666
rect 57250 17614 57262 17666
rect 57314 17614 57326 17666
rect 38894 17602 38946 17614
rect 51214 17602 51266 17614
rect 53454 17602 53506 17614
rect 16046 17554 16098 17566
rect 1922 17502 1934 17554
rect 1986 17502 1998 17554
rect 16046 17490 16098 17502
rect 16270 17554 16322 17566
rect 16270 17490 16322 17502
rect 17838 17554 17890 17566
rect 17838 17490 17890 17502
rect 18398 17554 18450 17566
rect 18398 17490 18450 17502
rect 18622 17554 18674 17566
rect 25342 17554 25394 17566
rect 21634 17502 21646 17554
rect 21698 17502 21710 17554
rect 18622 17490 18674 17502
rect 25342 17490 25394 17502
rect 25566 17554 25618 17566
rect 28478 17554 28530 17566
rect 28242 17502 28254 17554
rect 28306 17502 28318 17554
rect 25566 17490 25618 17502
rect 28478 17490 28530 17502
rect 28590 17554 28642 17566
rect 28590 17490 28642 17502
rect 29486 17554 29538 17566
rect 29486 17490 29538 17502
rect 29710 17554 29762 17566
rect 29710 17490 29762 17502
rect 31166 17554 31218 17566
rect 31166 17490 31218 17502
rect 31390 17554 31442 17566
rect 31390 17490 31442 17502
rect 31950 17554 32002 17566
rect 31950 17490 32002 17502
rect 33742 17554 33794 17566
rect 33742 17490 33794 17502
rect 35198 17554 35250 17566
rect 35198 17490 35250 17502
rect 37662 17554 37714 17566
rect 37662 17490 37714 17502
rect 38558 17554 38610 17566
rect 43934 17554 43986 17566
rect 50878 17554 50930 17566
rect 41906 17502 41918 17554
rect 41970 17502 41982 17554
rect 42578 17502 42590 17554
rect 42642 17502 42654 17554
rect 45714 17502 45726 17554
rect 45778 17502 45790 17554
rect 49746 17502 49758 17554
rect 49810 17502 49822 17554
rect 38558 17490 38610 17502
rect 43934 17490 43986 17502
rect 50878 17490 50930 17502
rect 56702 17554 56754 17566
rect 56702 17490 56754 17502
rect 17614 17442 17666 17454
rect 17614 17378 17666 17390
rect 18510 17442 18562 17454
rect 18510 17378 18562 17390
rect 23998 17442 24050 17454
rect 23998 17378 24050 17390
rect 25230 17442 25282 17454
rect 25230 17378 25282 17390
rect 26686 17442 26738 17454
rect 26686 17378 26738 17390
rect 26798 17442 26850 17454
rect 26798 17378 26850 17390
rect 26910 17442 26962 17454
rect 26910 17378 26962 17390
rect 28814 17442 28866 17454
rect 28814 17378 28866 17390
rect 30494 17442 30546 17454
rect 30494 17378 30546 17390
rect 32174 17442 32226 17454
rect 32174 17378 32226 17390
rect 32286 17442 32338 17454
rect 32286 17378 32338 17390
rect 33406 17442 33458 17454
rect 33406 17378 33458 17390
rect 33630 17442 33682 17454
rect 36318 17442 36370 17454
rect 35746 17390 35758 17442
rect 35810 17390 35822 17442
rect 33630 17378 33682 17390
rect 36318 17378 36370 17390
rect 37550 17442 37602 17454
rect 37550 17378 37602 17390
rect 38670 17442 38722 17454
rect 38670 17378 38722 17390
rect 40014 17442 40066 17454
rect 40014 17378 40066 17390
rect 40686 17442 40738 17454
rect 40686 17378 40738 17390
rect 44718 17442 44770 17454
rect 44718 17378 44770 17390
rect 50318 17442 50370 17454
rect 50318 17378 50370 17390
rect 52334 17442 52386 17454
rect 52334 17378 52386 17390
rect 53790 17442 53842 17454
rect 53790 17378 53842 17390
rect 54238 17442 54290 17454
rect 54238 17378 54290 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 2382 17106 2434 17118
rect 2382 17042 2434 17054
rect 3278 17106 3330 17118
rect 25790 17106 25842 17118
rect 16706 17054 16718 17106
rect 16770 17054 16782 17106
rect 22978 17054 22990 17106
rect 23042 17054 23054 17106
rect 3278 17042 3330 17054
rect 25790 17042 25842 17054
rect 25902 17106 25954 17118
rect 25902 17042 25954 17054
rect 26462 17106 26514 17118
rect 26462 17042 26514 17054
rect 27246 17106 27298 17118
rect 27246 17042 27298 17054
rect 28478 17106 28530 17118
rect 28478 17042 28530 17054
rect 28702 17106 28754 17118
rect 28702 17042 28754 17054
rect 28926 17106 28978 17118
rect 28926 17042 28978 17054
rect 29598 17106 29650 17118
rect 30494 17106 30546 17118
rect 29922 17054 29934 17106
rect 29986 17054 29998 17106
rect 29598 17042 29650 17054
rect 30494 17042 30546 17054
rect 31278 17106 31330 17118
rect 31278 17042 31330 17054
rect 31950 17106 32002 17118
rect 31950 17042 32002 17054
rect 32958 17106 33010 17118
rect 32958 17042 33010 17054
rect 34750 17106 34802 17118
rect 36766 17106 36818 17118
rect 35186 17054 35198 17106
rect 35250 17054 35262 17106
rect 34750 17042 34802 17054
rect 36766 17042 36818 17054
rect 39342 17106 39394 17118
rect 39342 17042 39394 17054
rect 40462 17106 40514 17118
rect 43934 17106 43986 17118
rect 42242 17054 42254 17106
rect 42306 17054 42318 17106
rect 40462 17042 40514 17054
rect 43934 17042 43986 17054
rect 45166 17106 45218 17118
rect 45166 17042 45218 17054
rect 45838 17106 45890 17118
rect 45838 17042 45890 17054
rect 46846 17106 46898 17118
rect 46846 17042 46898 17054
rect 48190 17106 48242 17118
rect 48190 17042 48242 17054
rect 51774 17106 51826 17118
rect 51774 17042 51826 17054
rect 51998 17106 52050 17118
rect 51998 17042 52050 17054
rect 53006 17106 53058 17118
rect 57474 17054 57486 17106
rect 57538 17054 57550 17106
rect 53006 17042 53058 17054
rect 2718 16994 2770 17006
rect 27470 16994 27522 17006
rect 15362 16942 15374 16994
rect 15426 16942 15438 16994
rect 16930 16942 16942 16994
rect 16994 16942 17006 16994
rect 24210 16942 24222 16994
rect 24274 16942 24286 16994
rect 2718 16930 2770 16942
rect 27470 16930 27522 16942
rect 27582 16994 27634 17006
rect 27582 16930 27634 16942
rect 33966 16994 34018 17006
rect 33966 16930 34018 16942
rect 34526 16994 34578 17006
rect 34526 16930 34578 16942
rect 37438 16994 37490 17006
rect 37438 16930 37490 16942
rect 37998 16994 38050 17006
rect 37998 16930 38050 16942
rect 38110 16994 38162 17006
rect 38110 16930 38162 16942
rect 38222 16994 38274 17006
rect 38222 16930 38274 16942
rect 40686 16994 40738 17006
rect 40686 16930 40738 16942
rect 40798 16994 40850 17006
rect 44718 16994 44770 17006
rect 42914 16942 42926 16994
rect 42978 16942 42990 16994
rect 40798 16930 40850 16942
rect 44718 16930 44770 16942
rect 46174 16994 46226 17006
rect 46174 16930 46226 16942
rect 50206 16994 50258 17006
rect 50206 16930 50258 16942
rect 53454 16994 53506 17006
rect 53454 16930 53506 16942
rect 54126 16994 54178 17006
rect 54126 16930 54178 16942
rect 54238 16994 54290 17006
rect 56702 16994 56754 17006
rect 55346 16942 55358 16994
rect 55410 16942 55422 16994
rect 54238 16930 54290 16942
rect 16382 16882 16434 16894
rect 30830 16882 30882 16894
rect 15922 16830 15934 16882
rect 15986 16830 15998 16882
rect 19954 16830 19966 16882
rect 20018 16830 20030 16882
rect 21298 16830 21310 16882
rect 21362 16830 21374 16882
rect 21634 16830 21646 16882
rect 21698 16830 21710 16882
rect 22978 16830 22990 16882
rect 23042 16830 23054 16882
rect 24658 16830 24670 16882
rect 24722 16830 24734 16882
rect 16382 16818 16434 16830
rect 30830 16818 30882 16830
rect 31838 16882 31890 16894
rect 31838 16818 31890 16830
rect 32062 16882 32114 16894
rect 32062 16818 32114 16830
rect 32510 16882 32562 16894
rect 34974 16882 35026 16894
rect 33618 16830 33630 16882
rect 33682 16830 33694 16882
rect 32510 16818 32562 16830
rect 34974 16818 35026 16830
rect 35198 16882 35250 16894
rect 35198 16818 35250 16830
rect 36318 16882 36370 16894
rect 36318 16818 36370 16830
rect 36542 16882 36594 16894
rect 41470 16882 41522 16894
rect 47406 16882 47458 16894
rect 52446 16882 52498 16894
rect 39442 16830 39454 16882
rect 39506 16830 39518 16882
rect 39890 16830 39902 16882
rect 39954 16830 39966 16882
rect 42018 16830 42030 16882
rect 42082 16830 42094 16882
rect 43138 16830 43150 16882
rect 43202 16830 43214 16882
rect 43922 16830 43934 16882
rect 43986 16830 43998 16882
rect 44482 16830 44494 16882
rect 44546 16830 44558 16882
rect 49858 16830 49870 16882
rect 49922 16830 49934 16882
rect 50866 16830 50878 16882
rect 50930 16830 50942 16882
rect 36542 16818 36594 16830
rect 41470 16818 41522 16830
rect 47406 16818 47458 16830
rect 52446 16818 52498 16830
rect 53230 16882 53282 16894
rect 53230 16818 53282 16830
rect 53902 16882 53954 16894
rect 53902 16818 53954 16830
rect 54686 16882 54738 16894
rect 54686 16818 54738 16830
rect 55134 16882 55186 16894
rect 55134 16818 55186 16830
rect 28814 16770 28866 16782
rect 28814 16706 28866 16718
rect 36094 16770 36146 16782
rect 48750 16770 48802 16782
rect 51886 16770 51938 16782
rect 36642 16718 36654 16770
rect 36706 16718 36718 16770
rect 49746 16718 49758 16770
rect 49810 16718 49822 16770
rect 50754 16718 50766 16770
rect 50818 16718 50830 16770
rect 36094 16706 36146 16718
rect 48750 16706 48802 16718
rect 51886 16706 51938 16718
rect 53342 16770 53394 16782
rect 53342 16706 53394 16718
rect 25678 16658 25730 16670
rect 25678 16594 25730 16606
rect 33630 16658 33682 16670
rect 33630 16594 33682 16606
rect 35870 16658 35922 16670
rect 38658 16606 38670 16658
rect 38722 16606 38734 16658
rect 44146 16606 44158 16658
rect 44210 16606 44222 16658
rect 54450 16606 54462 16658
rect 54514 16655 54526 16658
rect 55361 16655 55407 16942
rect 56702 16930 56754 16942
rect 57822 16882 57874 16894
rect 57822 16818 57874 16830
rect 54514 16609 55407 16655
rect 55582 16658 55634 16670
rect 54514 16606 54526 16609
rect 35870 16594 35922 16606
rect 55582 16594 55634 16606
rect 56030 16658 56082 16670
rect 56030 16594 56082 16606
rect 56254 16658 56306 16670
rect 56254 16594 56306 16606
rect 56478 16658 56530 16670
rect 56478 16594 56530 16606
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 14814 16322 14866 16334
rect 36430 16322 36482 16334
rect 28690 16270 28702 16322
rect 28754 16319 28766 16322
rect 28914 16319 28926 16322
rect 28754 16273 28926 16319
rect 28754 16270 28766 16273
rect 28914 16270 28926 16273
rect 28978 16270 28990 16322
rect 33506 16270 33518 16322
rect 33570 16319 33582 16322
rect 34738 16319 34750 16322
rect 33570 16273 34750 16319
rect 33570 16270 33582 16273
rect 34738 16270 34750 16273
rect 34802 16270 34814 16322
rect 14814 16258 14866 16270
rect 36430 16258 36482 16270
rect 36766 16322 36818 16334
rect 44382 16322 44434 16334
rect 43250 16270 43262 16322
rect 43314 16270 43326 16322
rect 36766 16258 36818 16270
rect 44382 16258 44434 16270
rect 47182 16322 47234 16334
rect 47182 16258 47234 16270
rect 48526 16322 48578 16334
rect 48526 16258 48578 16270
rect 50542 16322 50594 16334
rect 50542 16258 50594 16270
rect 16494 16210 16546 16222
rect 16494 16146 16546 16158
rect 19182 16210 19234 16222
rect 19182 16146 19234 16158
rect 19966 16210 20018 16222
rect 19966 16146 20018 16158
rect 21534 16210 21586 16222
rect 21534 16146 21586 16158
rect 23214 16210 23266 16222
rect 23214 16146 23266 16158
rect 25566 16210 25618 16222
rect 25566 16146 25618 16158
rect 26350 16210 26402 16222
rect 26350 16146 26402 16158
rect 28926 16210 28978 16222
rect 28926 16146 28978 16158
rect 29598 16210 29650 16222
rect 29598 16146 29650 16158
rect 29934 16210 29986 16222
rect 29934 16146 29986 16158
rect 33406 16210 33458 16222
rect 33406 16146 33458 16158
rect 34190 16210 34242 16222
rect 34190 16146 34242 16158
rect 34750 16210 34802 16222
rect 34750 16146 34802 16158
rect 35646 16210 35698 16222
rect 45390 16210 45442 16222
rect 41794 16158 41806 16210
rect 41858 16158 41870 16210
rect 44146 16158 44158 16210
rect 44210 16158 44222 16210
rect 35646 16146 35698 16158
rect 45390 16146 45442 16158
rect 47854 16210 47906 16222
rect 47854 16146 47906 16158
rect 51998 16210 52050 16222
rect 51998 16146 52050 16158
rect 52446 16210 52498 16222
rect 52446 16146 52498 16158
rect 53902 16210 53954 16222
rect 55918 16210 55970 16222
rect 55682 16158 55694 16210
rect 55746 16158 55758 16210
rect 53902 16146 53954 16158
rect 55918 16146 55970 16158
rect 16382 16098 16434 16110
rect 16034 16046 16046 16098
rect 16098 16046 16110 16098
rect 16382 16034 16434 16046
rect 17166 16098 17218 16110
rect 17166 16034 17218 16046
rect 24110 16098 24162 16110
rect 31390 16098 31442 16110
rect 24882 16046 24894 16098
rect 24946 16046 24958 16098
rect 24110 16034 24162 16046
rect 31390 16034 31442 16046
rect 32510 16098 32562 16110
rect 47294 16098 47346 16110
rect 38658 16046 38670 16098
rect 38722 16046 38734 16098
rect 39666 16046 39678 16098
rect 39730 16046 39742 16098
rect 40674 16046 40686 16098
rect 40738 16046 40750 16098
rect 42914 16046 42926 16098
rect 42978 16046 42990 16098
rect 43474 16046 43486 16098
rect 43538 16046 43550 16098
rect 46386 16046 46398 16098
rect 46450 16046 46462 16098
rect 32510 16034 32562 16046
rect 47294 16034 47346 16046
rect 48414 16098 48466 16110
rect 48414 16034 48466 16046
rect 49086 16098 49138 16110
rect 49086 16034 49138 16046
rect 49870 16098 49922 16110
rect 49870 16034 49922 16046
rect 50318 16098 50370 16110
rect 50318 16034 50370 16046
rect 56814 16098 56866 16110
rect 56814 16034 56866 16046
rect 14702 15986 14754 15998
rect 14702 15922 14754 15934
rect 18958 15986 19010 15998
rect 28030 15986 28082 15998
rect 24658 15934 24670 15986
rect 24722 15934 24734 15986
rect 18958 15922 19010 15934
rect 28030 15922 28082 15934
rect 28366 15986 28418 15998
rect 28366 15922 28418 15934
rect 32846 15986 32898 15998
rect 32846 15922 32898 15934
rect 33742 15986 33794 15998
rect 33742 15922 33794 15934
rect 36654 15986 36706 15998
rect 36654 15922 36706 15934
rect 37774 15986 37826 15998
rect 37774 15922 37826 15934
rect 38110 15986 38162 15998
rect 41918 15986 41970 15998
rect 40114 15934 40126 15986
rect 40178 15934 40190 15986
rect 40786 15934 40798 15986
rect 40850 15934 40862 15986
rect 38110 15922 38162 15934
rect 41918 15922 41970 15934
rect 42142 15986 42194 15998
rect 42142 15922 42194 15934
rect 42702 15986 42754 15998
rect 42702 15922 42754 15934
rect 44158 15986 44210 15998
rect 47182 15986 47234 15998
rect 46162 15934 46174 15986
rect 46226 15934 46238 15986
rect 44158 15922 44210 15934
rect 47182 15922 47234 15934
rect 48526 15986 48578 15998
rect 48526 15922 48578 15934
rect 49758 15986 49810 15998
rect 49758 15922 49810 15934
rect 50094 15986 50146 15998
rect 50094 15922 50146 15934
rect 51102 15986 51154 15998
rect 51102 15922 51154 15934
rect 55694 15986 55746 15998
rect 55694 15922 55746 15934
rect 57374 15986 57426 15998
rect 57374 15922 57426 15934
rect 57710 15986 57762 15998
rect 57710 15922 57762 15934
rect 14814 15874 14866 15886
rect 14814 15810 14866 15822
rect 17054 15874 17106 15886
rect 20414 15874 20466 15886
rect 19506 15822 19518 15874
rect 19570 15822 19582 15874
rect 17054 15810 17106 15822
rect 20414 15810 20466 15822
rect 21982 15874 22034 15886
rect 21982 15810 22034 15822
rect 23774 15874 23826 15886
rect 23774 15810 23826 15822
rect 26686 15874 26738 15886
rect 26686 15810 26738 15822
rect 27134 15874 27186 15886
rect 27134 15810 27186 15822
rect 31838 15874 31890 15886
rect 31838 15810 31890 15822
rect 31950 15874 32002 15886
rect 31950 15810 32002 15822
rect 32062 15874 32114 15886
rect 32062 15810 32114 15822
rect 32734 15874 32786 15886
rect 32734 15810 32786 15822
rect 35198 15874 35250 15886
rect 42814 15874 42866 15886
rect 39778 15822 39790 15874
rect 39842 15822 39854 15874
rect 35198 15810 35250 15822
rect 42814 15810 42866 15822
rect 51550 15874 51602 15886
rect 51550 15810 51602 15822
rect 53342 15874 53394 15886
rect 54798 15874 54850 15886
rect 54450 15822 54462 15874
rect 54514 15822 54526 15874
rect 56466 15822 56478 15874
rect 56530 15822 56542 15874
rect 53342 15810 53394 15822
rect 54798 15810 54850 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 16830 15538 16882 15550
rect 16034 15486 16046 15538
rect 16098 15486 16110 15538
rect 16830 15474 16882 15486
rect 18398 15538 18450 15550
rect 28254 15538 28306 15550
rect 27906 15486 27918 15538
rect 27970 15486 27982 15538
rect 18398 15474 18450 15486
rect 28254 15474 28306 15486
rect 29598 15538 29650 15550
rect 29598 15474 29650 15486
rect 30046 15538 30098 15550
rect 30046 15474 30098 15486
rect 37774 15538 37826 15550
rect 37774 15474 37826 15486
rect 38222 15538 38274 15550
rect 38222 15474 38274 15486
rect 40350 15538 40402 15550
rect 40350 15474 40402 15486
rect 42366 15538 42418 15550
rect 42366 15474 42418 15486
rect 43710 15538 43762 15550
rect 43710 15474 43762 15486
rect 44270 15538 44322 15550
rect 44270 15474 44322 15486
rect 45502 15538 45554 15550
rect 45502 15474 45554 15486
rect 46958 15538 47010 15550
rect 46958 15474 47010 15486
rect 49422 15538 49474 15550
rect 49422 15474 49474 15486
rect 52894 15538 52946 15550
rect 52894 15474 52946 15486
rect 55022 15538 55074 15550
rect 57810 15486 57822 15538
rect 57874 15486 57886 15538
rect 55022 15474 55074 15486
rect 26574 15426 26626 15438
rect 37326 15426 37378 15438
rect 14466 15374 14478 15426
rect 14530 15374 14542 15426
rect 15922 15374 15934 15426
rect 15986 15374 15998 15426
rect 20514 15374 20526 15426
rect 20578 15374 20590 15426
rect 21410 15374 21422 15426
rect 21474 15374 21486 15426
rect 34850 15374 34862 15426
rect 34914 15374 34926 15426
rect 26574 15362 26626 15374
rect 37326 15362 37378 15374
rect 42814 15426 42866 15438
rect 42814 15362 42866 15374
rect 44606 15426 44658 15438
rect 44606 15362 44658 15374
rect 45726 15426 45778 15438
rect 45726 15362 45778 15374
rect 48414 15426 48466 15438
rect 52670 15426 52722 15438
rect 50978 15374 50990 15426
rect 51042 15374 51054 15426
rect 51426 15374 51438 15426
rect 51490 15374 51502 15426
rect 48414 15362 48466 15374
rect 52670 15362 52722 15374
rect 54126 15426 54178 15438
rect 54126 15362 54178 15374
rect 56702 15426 56754 15438
rect 56702 15362 56754 15374
rect 25566 15314 25618 15326
rect 40798 15314 40850 15326
rect 14690 15262 14702 15314
rect 14754 15262 14766 15314
rect 19170 15262 19182 15314
rect 19234 15262 19246 15314
rect 22642 15262 22654 15314
rect 22706 15262 22718 15314
rect 24546 15262 24558 15314
rect 24610 15262 24622 15314
rect 26226 15262 26238 15314
rect 26290 15262 26302 15314
rect 29138 15262 29150 15314
rect 29202 15262 29214 15314
rect 33618 15262 33630 15314
rect 33682 15262 33694 15314
rect 33954 15262 33966 15314
rect 34018 15262 34030 15314
rect 35074 15262 35086 15314
rect 35138 15262 35150 15314
rect 35970 15262 35982 15314
rect 36034 15262 36046 15314
rect 36418 15262 36430 15314
rect 36482 15262 36494 15314
rect 39330 15262 39342 15314
rect 39394 15262 39406 15314
rect 39554 15262 39566 15314
rect 39618 15262 39630 15314
rect 25566 15250 25618 15262
rect 40798 15250 40850 15262
rect 41470 15314 41522 15326
rect 41470 15250 41522 15262
rect 46174 15314 46226 15326
rect 46174 15250 46226 15262
rect 47182 15314 47234 15326
rect 52558 15314 52610 15326
rect 47506 15262 47518 15314
rect 47570 15262 47582 15314
rect 50194 15262 50206 15314
rect 50258 15262 50270 15314
rect 50530 15262 50542 15314
rect 50594 15262 50606 15314
rect 51762 15262 51774 15314
rect 51826 15262 51838 15314
rect 47182 15250 47234 15262
rect 52558 15250 52610 15262
rect 53230 15314 53282 15326
rect 55806 15314 55858 15326
rect 53666 15262 53678 15314
rect 53730 15262 53742 15314
rect 53890 15262 53902 15314
rect 53954 15262 53966 15314
rect 54786 15262 54798 15314
rect 54850 15262 54862 15314
rect 53230 15250 53282 15262
rect 55806 15250 55858 15262
rect 56366 15314 56418 15326
rect 56366 15250 56418 15262
rect 57486 15314 57538 15326
rect 57486 15250 57538 15262
rect 26462 15202 26514 15214
rect 20402 15150 20414 15202
rect 20466 15150 20478 15202
rect 22530 15150 22542 15202
rect 22594 15150 22606 15202
rect 24434 15150 24446 15202
rect 24498 15150 24510 15202
rect 26462 15138 26514 15150
rect 27358 15202 27410 15214
rect 27358 15138 27410 15150
rect 32286 15202 32338 15214
rect 32286 15138 32338 15150
rect 32734 15202 32786 15214
rect 35758 15202 35810 15214
rect 41918 15202 41970 15214
rect 34962 15150 34974 15202
rect 35026 15150 35038 15202
rect 38882 15150 38894 15202
rect 38946 15150 38958 15202
rect 32734 15138 32786 15150
rect 35758 15138 35810 15150
rect 41918 15138 41970 15150
rect 43262 15202 43314 15214
rect 43262 15138 43314 15150
rect 47070 15202 47122 15214
rect 47070 15138 47122 15150
rect 47966 15202 48018 15214
rect 47966 15138 48018 15150
rect 55694 15202 55746 15214
rect 55694 15138 55746 15150
rect 28814 15090 28866 15102
rect 23762 15038 23774 15090
rect 23826 15038 23838 15090
rect 28814 15026 28866 15038
rect 29150 15090 29202 15102
rect 45390 15090 45442 15102
rect 38770 15038 38782 15090
rect 38834 15038 38846 15090
rect 40226 15038 40238 15090
rect 40290 15087 40302 15090
rect 41010 15087 41022 15090
rect 40290 15041 41022 15087
rect 40290 15038 40302 15041
rect 41010 15038 41022 15041
rect 41074 15038 41086 15090
rect 43138 15038 43150 15090
rect 43202 15087 43214 15090
rect 44146 15087 44158 15090
rect 43202 15041 44158 15087
rect 43202 15038 43214 15041
rect 44146 15038 44158 15041
rect 44210 15038 44222 15090
rect 29150 15026 29202 15038
rect 45390 15026 45442 15038
rect 54238 15090 54290 15102
rect 54238 15026 54290 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 14926 14754 14978 14766
rect 14926 14690 14978 14702
rect 16158 14754 16210 14766
rect 16158 14690 16210 14702
rect 36206 14754 36258 14766
rect 36206 14690 36258 14702
rect 52670 14754 52722 14766
rect 52670 14690 52722 14702
rect 14254 14642 14306 14654
rect 14254 14578 14306 14590
rect 17614 14642 17666 14654
rect 17614 14578 17666 14590
rect 18846 14642 18898 14654
rect 18846 14578 18898 14590
rect 20302 14642 20354 14654
rect 25678 14642 25730 14654
rect 33742 14642 33794 14654
rect 36766 14642 36818 14654
rect 21858 14590 21870 14642
rect 21922 14590 21934 14642
rect 22530 14590 22542 14642
rect 22594 14590 22606 14642
rect 28690 14590 28702 14642
rect 28754 14590 28766 14642
rect 31378 14590 31390 14642
rect 31442 14590 31454 14642
rect 35298 14590 35310 14642
rect 35362 14590 35374 14642
rect 20302 14578 20354 14590
rect 25678 14578 25730 14590
rect 33742 14578 33794 14590
rect 36766 14578 36818 14590
rect 37438 14642 37490 14654
rect 37438 14578 37490 14590
rect 37886 14642 37938 14654
rect 37886 14578 37938 14590
rect 48414 14642 48466 14654
rect 48414 14578 48466 14590
rect 48862 14642 48914 14654
rect 58046 14642 58098 14654
rect 50194 14590 50206 14642
rect 50258 14590 50270 14642
rect 53890 14590 53902 14642
rect 53954 14590 53966 14642
rect 48862 14578 48914 14590
rect 58046 14578 58098 14590
rect 14702 14530 14754 14542
rect 14702 14466 14754 14478
rect 18958 14530 19010 14542
rect 18958 14466 19010 14478
rect 19406 14530 19458 14542
rect 19406 14466 19458 14478
rect 20638 14530 20690 14542
rect 24222 14530 24274 14542
rect 21522 14478 21534 14530
rect 21586 14478 21598 14530
rect 22642 14478 22654 14530
rect 22706 14478 22718 14530
rect 20638 14466 20690 14478
rect 24222 14466 24274 14478
rect 24782 14530 24834 14542
rect 24782 14466 24834 14478
rect 25790 14530 25842 14542
rect 25790 14466 25842 14478
rect 26798 14530 26850 14542
rect 26798 14466 26850 14478
rect 27358 14530 27410 14542
rect 29486 14530 29538 14542
rect 36318 14530 36370 14542
rect 40798 14530 40850 14542
rect 28466 14478 28478 14530
rect 28530 14478 28542 14530
rect 31938 14478 31950 14530
rect 32002 14478 32014 14530
rect 35634 14478 35646 14530
rect 35698 14478 35710 14530
rect 39218 14478 39230 14530
rect 39282 14478 39294 14530
rect 40226 14478 40238 14530
rect 40290 14478 40302 14530
rect 27358 14466 27410 14478
rect 29486 14466 29538 14478
rect 36318 14466 36370 14478
rect 40798 14466 40850 14478
rect 41694 14530 41746 14542
rect 41694 14466 41746 14478
rect 41806 14530 41858 14542
rect 41806 14466 41858 14478
rect 42590 14530 42642 14542
rect 42590 14466 42642 14478
rect 42814 14530 42866 14542
rect 42814 14466 42866 14478
rect 43150 14530 43202 14542
rect 43150 14466 43202 14478
rect 45838 14530 45890 14542
rect 50542 14530 50594 14542
rect 55022 14530 55074 14542
rect 47730 14478 47742 14530
rect 47794 14478 47806 14530
rect 53442 14478 53454 14530
rect 53506 14478 53518 14530
rect 54226 14478 54238 14530
rect 54290 14478 54302 14530
rect 45838 14466 45890 14478
rect 50542 14466 50594 14478
rect 55022 14466 55074 14478
rect 57374 14530 57426 14542
rect 57374 14466 57426 14478
rect 13806 14418 13858 14430
rect 13806 14354 13858 14366
rect 15934 14418 15986 14430
rect 15934 14354 15986 14366
rect 17054 14418 17106 14430
rect 17054 14354 17106 14366
rect 20862 14418 20914 14430
rect 20862 14354 20914 14366
rect 24110 14418 24162 14430
rect 24110 14354 24162 14366
rect 27806 14418 27858 14430
rect 27806 14354 27858 14366
rect 29822 14418 29874 14430
rect 29822 14354 29874 14366
rect 31054 14418 31106 14430
rect 31054 14354 31106 14366
rect 35422 14418 35474 14430
rect 35422 14354 35474 14366
rect 39006 14418 39058 14430
rect 39006 14354 39058 14366
rect 40686 14418 40738 14430
rect 40686 14354 40738 14366
rect 44270 14418 44322 14430
rect 44270 14354 44322 14366
rect 45502 14418 45554 14430
rect 45502 14354 45554 14366
rect 47070 14418 47122 14430
rect 47070 14354 47122 14366
rect 49310 14418 49362 14430
rect 49310 14354 49362 14366
rect 51438 14418 51490 14430
rect 55134 14418 55186 14430
rect 54114 14366 54126 14418
rect 54178 14366 54190 14418
rect 51438 14354 51490 14366
rect 55134 14354 55186 14366
rect 55582 14418 55634 14430
rect 55582 14354 55634 14366
rect 56142 14418 56194 14430
rect 56142 14354 56194 14366
rect 16046 14306 16098 14318
rect 15250 14254 15262 14306
rect 15314 14254 15326 14306
rect 16046 14242 16098 14254
rect 16606 14306 16658 14318
rect 16606 14242 16658 14254
rect 17950 14306 18002 14318
rect 17950 14242 18002 14254
rect 18734 14306 18786 14318
rect 18734 14242 18786 14254
rect 23438 14306 23490 14318
rect 23438 14242 23490 14254
rect 24334 14306 24386 14318
rect 24334 14242 24386 14254
rect 25342 14306 25394 14318
rect 25342 14242 25394 14254
rect 25566 14306 25618 14318
rect 25566 14242 25618 14254
rect 26686 14306 26738 14318
rect 26686 14242 26738 14254
rect 26910 14306 26962 14318
rect 26910 14242 26962 14254
rect 29710 14306 29762 14318
rect 29710 14242 29762 14254
rect 30270 14306 30322 14318
rect 30270 14242 30322 14254
rect 33294 14306 33346 14318
rect 33294 14242 33346 14254
rect 35870 14306 35922 14318
rect 35870 14242 35922 14254
rect 38446 14306 38498 14318
rect 38446 14242 38498 14254
rect 39454 14306 39506 14318
rect 39454 14242 39506 14254
rect 39566 14306 39618 14318
rect 39566 14242 39618 14254
rect 40462 14306 40514 14318
rect 40462 14242 40514 14254
rect 41358 14306 41410 14318
rect 41358 14242 41410 14254
rect 41470 14306 41522 14318
rect 41470 14242 41522 14254
rect 41582 14306 41634 14318
rect 41582 14242 41634 14254
rect 42814 14306 42866 14318
rect 42814 14242 42866 14254
rect 44046 14306 44098 14318
rect 44046 14242 44098 14254
rect 44382 14306 44434 14318
rect 44382 14242 44434 14254
rect 44494 14306 44546 14318
rect 44494 14242 44546 14254
rect 46734 14306 46786 14318
rect 46734 14242 46786 14254
rect 47966 14306 48018 14318
rect 47966 14242 48018 14254
rect 50318 14306 50370 14318
rect 50318 14242 50370 14254
rect 51102 14306 51154 14318
rect 51102 14242 51154 14254
rect 52446 14306 52498 14318
rect 52446 14242 52498 14254
rect 52558 14306 52610 14318
rect 52558 14242 52610 14254
rect 55358 14306 55410 14318
rect 57038 14306 57090 14318
rect 56466 14254 56478 14306
rect 56530 14254 56542 14306
rect 55358 14242 55410 14254
rect 57038 14242 57090 14254
rect 57934 14306 57986 14318
rect 57934 14242 57986 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 13918 13970 13970 13982
rect 13918 13906 13970 13918
rect 15710 13970 15762 13982
rect 15710 13906 15762 13918
rect 16494 13970 16546 13982
rect 19742 13970 19794 13982
rect 18722 13918 18734 13970
rect 18786 13918 18798 13970
rect 16494 13906 16546 13918
rect 19742 13906 19794 13918
rect 20190 13970 20242 13982
rect 20190 13906 20242 13918
rect 22990 13970 23042 13982
rect 22990 13906 23042 13918
rect 24558 13970 24610 13982
rect 24558 13906 24610 13918
rect 26014 13970 26066 13982
rect 26014 13906 26066 13918
rect 26126 13970 26178 13982
rect 26126 13906 26178 13918
rect 26238 13970 26290 13982
rect 26238 13906 26290 13918
rect 31390 13970 31442 13982
rect 31390 13906 31442 13918
rect 35198 13970 35250 13982
rect 35198 13906 35250 13918
rect 37214 13970 37266 13982
rect 37214 13906 37266 13918
rect 40574 13970 40626 13982
rect 40574 13906 40626 13918
rect 42590 13970 42642 13982
rect 42590 13906 42642 13918
rect 43934 13970 43986 13982
rect 43934 13906 43986 13918
rect 44046 13970 44098 13982
rect 44046 13906 44098 13918
rect 44830 13970 44882 13982
rect 44830 13906 44882 13918
rect 45726 13970 45778 13982
rect 48190 13970 48242 13982
rect 46834 13918 46846 13970
rect 46898 13918 46910 13970
rect 45726 13906 45778 13918
rect 48190 13906 48242 13918
rect 50542 13970 50594 13982
rect 50542 13906 50594 13918
rect 51438 13970 51490 13982
rect 51438 13906 51490 13918
rect 52446 13970 52498 13982
rect 52446 13906 52498 13918
rect 55134 13970 55186 13982
rect 55134 13906 55186 13918
rect 55806 13970 55858 13982
rect 55806 13906 55858 13918
rect 56142 13970 56194 13982
rect 56142 13906 56194 13918
rect 57374 13970 57426 13982
rect 57374 13906 57426 13918
rect 15822 13858 15874 13870
rect 15822 13794 15874 13806
rect 16718 13858 16770 13870
rect 16718 13794 16770 13806
rect 22542 13858 22594 13870
rect 31278 13858 31330 13870
rect 24882 13806 24894 13858
rect 24946 13806 24958 13858
rect 28354 13806 28366 13858
rect 28418 13806 28430 13858
rect 22542 13794 22594 13806
rect 31278 13794 31330 13806
rect 36206 13858 36258 13870
rect 36206 13794 36258 13806
rect 38110 13858 38162 13870
rect 39566 13858 39618 13870
rect 39330 13806 39342 13858
rect 39394 13806 39406 13858
rect 38110 13794 38162 13806
rect 39566 13794 39618 13806
rect 39678 13858 39730 13870
rect 39678 13794 39730 13806
rect 40350 13858 40402 13870
rect 40350 13794 40402 13806
rect 41918 13858 41970 13870
rect 49982 13858 50034 13870
rect 53118 13858 53170 13870
rect 46722 13806 46734 13858
rect 46786 13806 46798 13858
rect 50866 13806 50878 13858
rect 50930 13806 50942 13858
rect 41918 13794 41970 13806
rect 49982 13794 50034 13806
rect 53118 13794 53170 13806
rect 53454 13858 53506 13870
rect 53454 13794 53506 13806
rect 54126 13858 54178 13870
rect 54126 13794 54178 13806
rect 54462 13858 54514 13870
rect 54462 13794 54514 13806
rect 55358 13858 55410 13870
rect 55358 13794 55410 13806
rect 14478 13746 14530 13758
rect 14478 13682 14530 13694
rect 14702 13746 14754 13758
rect 15486 13746 15538 13758
rect 14914 13694 14926 13746
rect 14978 13694 14990 13746
rect 14702 13682 14754 13694
rect 15486 13682 15538 13694
rect 16046 13746 16098 13758
rect 16046 13682 16098 13694
rect 16830 13746 16882 13758
rect 16830 13682 16882 13694
rect 19070 13746 19122 13758
rect 22318 13746 22370 13758
rect 21970 13694 21982 13746
rect 22034 13694 22046 13746
rect 19070 13682 19122 13694
rect 22318 13682 22370 13694
rect 25566 13746 25618 13758
rect 25566 13682 25618 13694
rect 27806 13746 27858 13758
rect 30270 13746 30322 13758
rect 28466 13694 28478 13746
rect 28530 13694 28542 13746
rect 29250 13694 29262 13746
rect 29314 13694 29326 13746
rect 27806 13682 27858 13694
rect 30270 13682 30322 13694
rect 35758 13746 35810 13758
rect 35758 13682 35810 13694
rect 36542 13746 36594 13758
rect 38670 13746 38722 13758
rect 38322 13694 38334 13746
rect 38386 13694 38398 13746
rect 36542 13682 36594 13694
rect 38670 13682 38722 13694
rect 39902 13746 39954 13758
rect 39902 13682 39954 13694
rect 40686 13746 40738 13758
rect 40686 13682 40738 13694
rect 41806 13746 41858 13758
rect 41806 13682 41858 13694
rect 42142 13746 42194 13758
rect 42142 13682 42194 13694
rect 43374 13746 43426 13758
rect 46510 13746 46562 13758
rect 48414 13746 48466 13758
rect 43698 13694 43710 13746
rect 43762 13694 43774 13746
rect 47170 13694 47182 13746
rect 47234 13694 47246 13746
rect 43374 13682 43426 13694
rect 46510 13682 46562 13694
rect 48414 13682 48466 13694
rect 49422 13746 49474 13758
rect 51774 13746 51826 13758
rect 49746 13694 49758 13746
rect 49810 13694 49822 13746
rect 49422 13682 49474 13694
rect 51774 13682 51826 13694
rect 52222 13746 52274 13758
rect 52222 13682 52274 13694
rect 52558 13746 52610 13758
rect 52558 13682 52610 13694
rect 55022 13746 55074 13758
rect 55022 13682 55074 13694
rect 19294 13634 19346 13646
rect 19294 13570 19346 13582
rect 20862 13634 20914 13646
rect 20862 13570 20914 13582
rect 23438 13634 23490 13646
rect 23438 13570 23490 13582
rect 28926 13634 28978 13646
rect 32398 13634 32450 13646
rect 42926 13634 42978 13646
rect 29138 13582 29150 13634
rect 29202 13582 29214 13634
rect 39106 13582 39118 13634
rect 39170 13582 39182 13634
rect 28926 13570 28978 13582
rect 32398 13570 32450 13582
rect 42926 13570 42978 13582
rect 44382 13634 44434 13646
rect 44382 13570 44434 13582
rect 45278 13634 45330 13646
rect 45278 13570 45330 13582
rect 48302 13634 48354 13646
rect 56590 13634 56642 13646
rect 49970 13582 49982 13634
rect 50034 13582 50046 13634
rect 48302 13570 48354 13582
rect 56590 13570 56642 13582
rect 57822 13634 57874 13646
rect 57822 13570 57874 13582
rect 14366 13522 14418 13534
rect 31502 13522 31554 13534
rect 19506 13470 19518 13522
rect 19570 13519 19582 13522
rect 20178 13519 20190 13522
rect 19570 13473 20190 13519
rect 19570 13470 19582 13473
rect 20178 13470 20190 13473
rect 20242 13470 20254 13522
rect 14366 13458 14418 13470
rect 31502 13458 31554 13470
rect 37998 13522 38050 13534
rect 47058 13470 47070 13522
rect 47122 13470 47134 13522
rect 37998 13458 38050 13470
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 15262 13186 15314 13198
rect 15262 13122 15314 13134
rect 15934 13186 15986 13198
rect 15934 13122 15986 13134
rect 16382 13186 16434 13198
rect 16382 13122 16434 13134
rect 28254 13186 28306 13198
rect 28254 13122 28306 13134
rect 29934 13186 29986 13198
rect 29934 13122 29986 13134
rect 36094 13186 36146 13198
rect 36094 13122 36146 13134
rect 15038 13074 15090 13086
rect 15038 13010 15090 13022
rect 16494 13074 16546 13086
rect 16494 13010 16546 13022
rect 20862 13074 20914 13086
rect 20862 13010 20914 13022
rect 21534 13074 21586 13086
rect 21534 13010 21586 13022
rect 28590 13074 28642 13086
rect 30494 13074 30546 13086
rect 29586 13022 29598 13074
rect 29650 13022 29662 13074
rect 28590 13010 28642 13022
rect 30494 13010 30546 13022
rect 31614 13074 31666 13086
rect 31614 13010 31666 13022
rect 34862 13074 34914 13086
rect 34862 13010 34914 13022
rect 37550 13074 37602 13086
rect 37550 13010 37602 13022
rect 38334 13074 38386 13086
rect 38334 13010 38386 13022
rect 39230 13074 39282 13086
rect 39230 13010 39282 13022
rect 39454 13074 39506 13086
rect 39454 13010 39506 13022
rect 41246 13074 41298 13086
rect 41246 13010 41298 13022
rect 41582 13074 41634 13086
rect 41582 13010 41634 13022
rect 43486 13074 43538 13086
rect 43486 13010 43538 13022
rect 45502 13074 45554 13086
rect 45502 13010 45554 13022
rect 45950 13074 46002 13086
rect 45950 13010 46002 13022
rect 52670 13074 52722 13086
rect 57262 13074 57314 13086
rect 53778 13022 53790 13074
rect 53842 13022 53854 13074
rect 54898 13022 54910 13074
rect 54962 13022 54974 13074
rect 52670 13010 52722 13022
rect 57262 13010 57314 13022
rect 15486 12962 15538 12974
rect 15486 12898 15538 12910
rect 24670 12962 24722 12974
rect 24670 12898 24722 12910
rect 25118 12962 25170 12974
rect 31950 12962 32002 12974
rect 26002 12910 26014 12962
rect 26066 12910 26078 12962
rect 25118 12898 25170 12910
rect 31950 12898 32002 12910
rect 32958 12962 33010 12974
rect 32958 12898 33010 12910
rect 33182 12962 33234 12974
rect 33182 12898 33234 12910
rect 33966 12962 34018 12974
rect 33966 12898 34018 12910
rect 35086 12962 35138 12974
rect 35086 12898 35138 12910
rect 42702 12962 42754 12974
rect 42702 12898 42754 12910
rect 42926 12962 42978 12974
rect 42926 12898 42978 12910
rect 44158 12962 44210 12974
rect 44158 12898 44210 12910
rect 44382 12962 44434 12974
rect 44382 12898 44434 12910
rect 46510 12962 46562 12974
rect 46510 12898 46562 12910
rect 46734 12962 46786 12974
rect 48626 12910 48638 12962
rect 48690 12910 48702 12962
rect 50306 12910 50318 12962
rect 50370 12910 50382 12962
rect 51874 12910 51886 12962
rect 51938 12910 51950 12962
rect 54226 12910 54238 12962
rect 54290 12910 54302 12962
rect 46734 12898 46786 12910
rect 18958 12850 19010 12862
rect 18958 12786 19010 12798
rect 19854 12850 19906 12862
rect 19854 12786 19906 12798
rect 19966 12850 20018 12862
rect 19966 12786 20018 12798
rect 25454 12850 25506 12862
rect 25454 12786 25506 12798
rect 28814 12850 28866 12862
rect 28814 12786 28866 12798
rect 31502 12850 31554 12862
rect 31502 12786 31554 12798
rect 31838 12850 31890 12862
rect 33854 12850 33906 12862
rect 32610 12798 32622 12850
rect 32674 12798 32686 12850
rect 31838 12786 31890 12798
rect 33854 12786 33906 12798
rect 34750 12850 34802 12862
rect 34750 12786 34802 12798
rect 35310 12850 35362 12862
rect 35310 12786 35362 12798
rect 35870 12850 35922 12862
rect 35870 12786 35922 12798
rect 42366 12850 42418 12862
rect 53454 12850 53506 12862
rect 48850 12798 48862 12850
rect 48914 12798 48926 12850
rect 51426 12798 51438 12850
rect 51490 12798 51502 12850
rect 42366 12786 42418 12798
rect 53454 12786 53506 12798
rect 53790 12850 53842 12862
rect 56130 12798 56142 12850
rect 56194 12798 56206 12850
rect 53790 12786 53842 12798
rect 18510 12738 18562 12750
rect 18510 12674 18562 12686
rect 19070 12738 19122 12750
rect 19070 12674 19122 12686
rect 19294 12738 19346 12750
rect 19294 12674 19346 12686
rect 19630 12738 19682 12750
rect 19630 12674 19682 12686
rect 20526 12738 20578 12750
rect 20526 12674 20578 12686
rect 26350 12738 26402 12750
rect 26350 12674 26402 12686
rect 26462 12738 26514 12750
rect 26462 12674 26514 12686
rect 26574 12738 26626 12750
rect 26574 12674 26626 12686
rect 29710 12738 29762 12750
rect 29710 12674 29762 12686
rect 30942 12738 30994 12750
rect 30942 12674 30994 12686
rect 33630 12738 33682 12750
rect 37886 12738 37938 12750
rect 40350 12738 40402 12750
rect 42814 12738 42866 12750
rect 46622 12738 46674 12750
rect 36418 12686 36430 12738
rect 36482 12686 36494 12738
rect 39778 12686 39790 12738
rect 39842 12686 39854 12738
rect 40674 12686 40686 12738
rect 40738 12686 40750 12738
rect 44706 12686 44718 12738
rect 44770 12686 44782 12738
rect 33630 12674 33682 12686
rect 37886 12674 37938 12686
rect 40350 12674 40402 12686
rect 42814 12674 42866 12686
rect 46622 12674 46674 12686
rect 46958 12738 47010 12750
rect 46958 12674 47010 12686
rect 47518 12738 47570 12750
rect 47518 12674 47570 12686
rect 49646 12738 49698 12750
rect 49646 12674 49698 12686
rect 53678 12738 53730 12750
rect 53678 12674 53730 12686
rect 56814 12738 56866 12750
rect 56814 12674 56866 12686
rect 57710 12738 57762 12750
rect 57710 12674 57762 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 2718 12402 2770 12414
rect 2718 12338 2770 12350
rect 15150 12402 15202 12414
rect 15150 12338 15202 12350
rect 15374 12402 15426 12414
rect 15374 12338 15426 12350
rect 24894 12402 24946 12414
rect 24894 12338 24946 12350
rect 29262 12402 29314 12414
rect 29262 12338 29314 12350
rect 30382 12402 30434 12414
rect 30382 12338 30434 12350
rect 31166 12402 31218 12414
rect 31166 12338 31218 12350
rect 34750 12402 34802 12414
rect 34750 12338 34802 12350
rect 35198 12402 35250 12414
rect 39342 12402 39394 12414
rect 36642 12350 36654 12402
rect 36706 12350 36718 12402
rect 35198 12338 35250 12350
rect 39342 12338 39394 12350
rect 39678 12402 39730 12414
rect 39678 12338 39730 12350
rect 40238 12402 40290 12414
rect 40238 12338 40290 12350
rect 42030 12402 42082 12414
rect 42030 12338 42082 12350
rect 42814 12402 42866 12414
rect 42814 12338 42866 12350
rect 43710 12402 43762 12414
rect 43710 12338 43762 12350
rect 44270 12402 44322 12414
rect 44270 12338 44322 12350
rect 47182 12402 47234 12414
rect 47182 12338 47234 12350
rect 48750 12402 48802 12414
rect 51662 12402 51714 12414
rect 49522 12350 49534 12402
rect 49586 12350 49598 12402
rect 48750 12338 48802 12350
rect 51662 12338 51714 12350
rect 52222 12402 52274 12414
rect 52222 12338 52274 12350
rect 53454 12402 53506 12414
rect 53454 12338 53506 12350
rect 54126 12402 54178 12414
rect 54126 12338 54178 12350
rect 54686 12402 54738 12414
rect 54686 12338 54738 12350
rect 55134 12402 55186 12414
rect 55134 12338 55186 12350
rect 56030 12402 56082 12414
rect 56030 12338 56082 12350
rect 56590 12402 56642 12414
rect 56590 12338 56642 12350
rect 57374 12402 57426 12414
rect 57374 12338 57426 12350
rect 27246 12290 27298 12302
rect 27246 12226 27298 12238
rect 28254 12290 28306 12302
rect 28254 12226 28306 12238
rect 28590 12290 28642 12302
rect 28590 12226 28642 12238
rect 32622 12290 32674 12302
rect 32622 12226 32674 12238
rect 37102 12290 37154 12302
rect 37102 12226 37154 12238
rect 40574 12290 40626 12302
rect 50990 12290 51042 12302
rect 45490 12238 45502 12290
rect 45554 12238 45566 12290
rect 46162 12238 46174 12290
rect 46226 12238 46238 12290
rect 40574 12226 40626 12238
rect 50990 12226 51042 12238
rect 54238 12290 54290 12302
rect 54238 12226 54290 12238
rect 15262 12178 15314 12190
rect 18622 12178 18674 12190
rect 21198 12178 21250 12190
rect 2482 12126 2494 12178
rect 2546 12126 2558 12178
rect 15698 12126 15710 12178
rect 15762 12126 15774 12178
rect 19506 12126 19518 12178
rect 19570 12126 19582 12178
rect 20850 12126 20862 12178
rect 20914 12126 20926 12178
rect 15262 12114 15314 12126
rect 18622 12114 18674 12126
rect 21198 12114 21250 12126
rect 21982 12178 22034 12190
rect 25902 12178 25954 12190
rect 22642 12126 22654 12178
rect 22706 12126 22718 12178
rect 21982 12114 22034 12126
rect 25902 12114 25954 12126
rect 26350 12178 26402 12190
rect 28702 12178 28754 12190
rect 27570 12126 27582 12178
rect 27634 12126 27646 12178
rect 26350 12114 26402 12126
rect 28702 12114 28754 12126
rect 31054 12178 31106 12190
rect 31502 12178 31554 12190
rect 32510 12178 32562 12190
rect 31266 12126 31278 12178
rect 31330 12126 31342 12178
rect 31826 12126 31838 12178
rect 31890 12126 31902 12178
rect 31054 12114 31106 12126
rect 31502 12114 31554 12126
rect 32510 12114 32562 12126
rect 35534 12178 35586 12190
rect 35534 12114 35586 12126
rect 35870 12178 35922 12190
rect 35870 12114 35922 12126
rect 37214 12178 37266 12190
rect 37214 12114 37266 12126
rect 37326 12178 37378 12190
rect 37326 12114 37378 12126
rect 38782 12178 38834 12190
rect 38782 12114 38834 12126
rect 42590 12178 42642 12190
rect 42590 12114 42642 12126
rect 43262 12178 43314 12190
rect 47406 12178 47458 12190
rect 44818 12126 44830 12178
rect 44882 12126 44894 12178
rect 45714 12126 45726 12178
rect 45778 12126 45790 12178
rect 46498 12126 46510 12178
rect 46562 12126 46574 12178
rect 43262 12114 43314 12126
rect 47406 12114 47458 12126
rect 47854 12178 47906 12190
rect 47854 12114 47906 12126
rect 49870 12178 49922 12190
rect 49870 12114 49922 12126
rect 50094 12178 50146 12190
rect 51550 12178 51602 12190
rect 50754 12126 50766 12178
rect 50818 12126 50830 12178
rect 50094 12114 50146 12126
rect 51550 12114 51602 12126
rect 53230 12178 53282 12190
rect 53230 12114 53282 12126
rect 53566 12178 53618 12190
rect 53566 12114 53618 12126
rect 3166 12066 3218 12078
rect 20302 12066 20354 12078
rect 27358 12066 27410 12078
rect 19394 12014 19406 12066
rect 19458 12014 19470 12066
rect 22866 12014 22878 12066
rect 22930 12014 22942 12066
rect 3166 12002 3218 12014
rect 20302 12002 20354 12014
rect 27358 12002 27410 12014
rect 28366 12066 28418 12078
rect 28366 12002 28418 12014
rect 29934 12066 29986 12078
rect 29934 12002 29986 12014
rect 30494 12066 30546 12078
rect 30494 12002 30546 12014
rect 33518 12066 33570 12078
rect 33518 12002 33570 12014
rect 33966 12066 34018 12078
rect 33966 12002 34018 12014
rect 41470 12066 41522 12078
rect 41470 12002 41522 12014
rect 42702 12066 42754 12078
rect 42702 12002 42754 12014
rect 47294 12066 47346 12078
rect 47294 12002 47346 12014
rect 48190 12066 48242 12078
rect 48190 12002 48242 12014
rect 52670 12066 52722 12078
rect 52670 12002 52722 12014
rect 55694 12066 55746 12078
rect 55694 12002 55746 12014
rect 57822 12066 57874 12078
rect 57822 12002 57874 12014
rect 26126 11954 26178 11966
rect 26126 11890 26178 11902
rect 26798 11954 26850 11966
rect 26798 11890 26850 11902
rect 32398 11954 32450 11966
rect 32398 11890 32450 11902
rect 35310 11954 35362 11966
rect 35310 11890 35362 11902
rect 36094 11954 36146 11966
rect 36094 11890 36146 11902
rect 51662 11954 51714 11966
rect 51662 11890 51714 11902
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 31390 11618 31442 11630
rect 42814 11618 42866 11630
rect 22866 11566 22878 11618
rect 22930 11566 22942 11618
rect 25666 11566 25678 11618
rect 25730 11566 25742 11618
rect 28802 11566 28814 11618
rect 28866 11615 28878 11618
rect 29026 11615 29038 11618
rect 28866 11569 29038 11615
rect 28866 11566 28878 11569
rect 29026 11566 29038 11569
rect 29090 11566 29102 11618
rect 32498 11566 32510 11618
rect 32562 11566 32574 11618
rect 39218 11566 39230 11618
rect 39282 11615 39294 11618
rect 39778 11615 39790 11618
rect 39282 11569 39790 11615
rect 39282 11566 39294 11569
rect 39778 11566 39790 11569
rect 39842 11566 39854 11618
rect 31390 11554 31442 11566
rect 42814 11554 42866 11566
rect 43150 11618 43202 11630
rect 43150 11554 43202 11566
rect 44158 11618 44210 11630
rect 44158 11554 44210 11566
rect 44382 11618 44434 11630
rect 44382 11554 44434 11566
rect 44830 11618 44882 11630
rect 44830 11554 44882 11566
rect 46958 11618 47010 11630
rect 47394 11566 47406 11618
rect 47458 11615 47470 11618
rect 48178 11615 48190 11618
rect 47458 11569 48190 11615
rect 47458 11566 47470 11569
rect 48178 11566 48190 11569
rect 48242 11566 48254 11618
rect 54562 11566 54574 11618
rect 54626 11615 54638 11618
rect 55458 11615 55470 11618
rect 54626 11569 55470 11615
rect 54626 11566 54638 11569
rect 55458 11566 55470 11569
rect 55522 11615 55534 11618
rect 55906 11615 55918 11618
rect 55522 11569 55918 11615
rect 55522 11566 55534 11569
rect 55906 11566 55918 11569
rect 55970 11566 55982 11618
rect 56354 11566 56366 11618
rect 56418 11615 56430 11618
rect 56802 11615 56814 11618
rect 56418 11569 56814 11615
rect 56418 11566 56430 11569
rect 56802 11566 56814 11569
rect 56866 11566 56878 11618
rect 46958 11554 47010 11566
rect 14254 11506 14306 11518
rect 14254 11442 14306 11454
rect 18286 11506 18338 11518
rect 18286 11442 18338 11454
rect 20526 11506 20578 11518
rect 20526 11442 20578 11454
rect 21870 11506 21922 11518
rect 28814 11506 28866 11518
rect 23202 11454 23214 11506
rect 23266 11454 23278 11506
rect 21870 11442 21922 11454
rect 28814 11442 28866 11454
rect 32062 11506 32114 11518
rect 32062 11442 32114 11454
rect 34190 11506 34242 11518
rect 34190 11442 34242 11454
rect 36206 11506 36258 11518
rect 36206 11442 36258 11454
rect 36766 11506 36818 11518
rect 36766 11442 36818 11454
rect 38782 11506 38834 11518
rect 38782 11442 38834 11454
rect 39118 11506 39170 11518
rect 39118 11442 39170 11454
rect 39790 11506 39842 11518
rect 39790 11442 39842 11454
rect 40126 11506 40178 11518
rect 40126 11442 40178 11454
rect 40574 11506 40626 11518
rect 40574 11442 40626 11454
rect 41582 11506 41634 11518
rect 41582 11442 41634 11454
rect 43262 11506 43314 11518
rect 43262 11442 43314 11454
rect 48302 11506 48354 11518
rect 48302 11442 48354 11454
rect 49198 11506 49250 11518
rect 49198 11442 49250 11454
rect 51102 11506 51154 11518
rect 51102 11442 51154 11454
rect 51662 11506 51714 11518
rect 51662 11442 51714 11454
rect 55134 11506 55186 11518
rect 55134 11442 55186 11454
rect 55582 11506 55634 11518
rect 55582 11442 55634 11454
rect 55918 11506 55970 11518
rect 55918 11442 55970 11454
rect 56814 11506 56866 11518
rect 56814 11442 56866 11454
rect 57374 11506 57426 11518
rect 57374 11442 57426 11454
rect 15150 11394 15202 11406
rect 2818 11342 2830 11394
rect 2882 11342 2894 11394
rect 14914 11342 14926 11394
rect 14978 11342 14990 11394
rect 15150 11330 15202 11342
rect 15710 11394 15762 11406
rect 15710 11330 15762 11342
rect 19742 11394 19794 11406
rect 19742 11330 19794 11342
rect 19854 11394 19906 11406
rect 23998 11394 24050 11406
rect 27918 11394 27970 11406
rect 23090 11342 23102 11394
rect 23154 11342 23166 11394
rect 24994 11342 25006 11394
rect 25058 11342 25070 11394
rect 25218 11342 25230 11394
rect 25282 11342 25294 11394
rect 26338 11342 26350 11394
rect 26402 11342 26414 11394
rect 19854 11330 19906 11342
rect 23998 11330 24050 11342
rect 27918 11330 27970 11342
rect 28254 11394 28306 11406
rect 30606 11394 30658 11406
rect 29586 11342 29598 11394
rect 29650 11342 29662 11394
rect 28254 11330 28306 11342
rect 30606 11330 30658 11342
rect 31054 11394 31106 11406
rect 31054 11330 31106 11342
rect 31950 11394 32002 11406
rect 33630 11394 33682 11406
rect 32610 11342 32622 11394
rect 32674 11342 32686 11394
rect 31950 11330 32002 11342
rect 33630 11330 33682 11342
rect 42926 11394 42978 11406
rect 42926 11330 42978 11342
rect 43934 11394 43986 11406
rect 43934 11330 43986 11342
rect 45614 11394 45666 11406
rect 45614 11330 45666 11342
rect 45950 11394 46002 11406
rect 50430 11394 50482 11406
rect 46162 11342 46174 11394
rect 46226 11342 46238 11394
rect 46386 11342 46398 11394
rect 46450 11391 46462 11394
rect 46722 11391 46734 11394
rect 46450 11345 46734 11391
rect 46450 11342 46462 11345
rect 46722 11342 46734 11345
rect 46786 11342 46798 11394
rect 49970 11342 49982 11394
rect 50034 11342 50046 11394
rect 45950 11330 46002 11342
rect 50430 11330 50482 11342
rect 50654 11394 50706 11406
rect 50654 11330 50706 11342
rect 53566 11394 53618 11406
rect 53566 11330 53618 11342
rect 53678 11394 53730 11406
rect 53678 11330 53730 11342
rect 53790 11394 53842 11406
rect 53790 11330 53842 11342
rect 54014 11394 54066 11406
rect 54014 11330 54066 11342
rect 15934 11282 15986 11294
rect 1922 11230 1934 11282
rect 1986 11230 1998 11282
rect 15934 11218 15986 11230
rect 16046 11282 16098 11294
rect 16046 11218 16098 11230
rect 19630 11282 19682 11294
rect 19630 11218 19682 11230
rect 27582 11282 27634 11294
rect 27582 11218 27634 11230
rect 29934 11282 29986 11294
rect 35982 11282 36034 11294
rect 32162 11230 32174 11282
rect 32226 11230 32238 11282
rect 35858 11230 35870 11282
rect 35922 11230 35934 11282
rect 29934 11218 29986 11230
rect 35982 11218 36034 11230
rect 37550 11282 37602 11294
rect 37550 11218 37602 11230
rect 37886 11282 37938 11294
rect 37886 11218 37938 11230
rect 46846 11282 46898 11294
rect 46846 11218 46898 11230
rect 48750 11282 48802 11294
rect 48750 11218 48802 11230
rect 50318 11282 50370 11294
rect 50318 11218 50370 11230
rect 52446 11282 52498 11294
rect 52446 11218 52498 11230
rect 18174 11170 18226 11182
rect 24110 11170 24162 11182
rect 19170 11118 19182 11170
rect 19234 11118 19246 11170
rect 18174 11106 18226 11118
rect 24110 11106 24162 11118
rect 24334 11170 24386 11182
rect 24334 11106 24386 11118
rect 26686 11170 26738 11182
rect 26686 11106 26738 11118
rect 28030 11170 28082 11182
rect 28030 11106 28082 11118
rect 29822 11170 29874 11182
rect 29822 11106 29874 11118
rect 31278 11170 31330 11182
rect 31278 11106 31330 11118
rect 33182 11170 33234 11182
rect 33182 11106 33234 11118
rect 36094 11170 36146 11182
rect 36094 11106 36146 11118
rect 36318 11170 36370 11182
rect 36318 11106 36370 11118
rect 41134 11170 41186 11182
rect 41134 11106 41186 11118
rect 42030 11170 42082 11182
rect 42030 11106 42082 11118
rect 45726 11170 45778 11182
rect 45726 11106 45778 11118
rect 45838 11170 45890 11182
rect 45838 11106 45890 11118
rect 47406 11170 47458 11182
rect 47406 11106 47458 11118
rect 47854 11170 47906 11182
rect 47854 11106 47906 11118
rect 49646 11170 49698 11182
rect 49646 11106 49698 11118
rect 52558 11170 52610 11182
rect 52558 11106 52610 11118
rect 53902 11170 53954 11182
rect 53902 11106 53954 11118
rect 54574 11170 54626 11182
rect 54574 11106 54626 11118
rect 56366 11170 56418 11182
rect 56366 11106 56418 11118
rect 57710 11170 57762 11182
rect 57710 11106 57762 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 2382 10834 2434 10846
rect 2382 10770 2434 10782
rect 3278 10834 3330 10846
rect 3278 10770 3330 10782
rect 14814 10834 14866 10846
rect 14814 10770 14866 10782
rect 16606 10834 16658 10846
rect 16606 10770 16658 10782
rect 17950 10834 18002 10846
rect 17950 10770 18002 10782
rect 24894 10834 24946 10846
rect 24894 10770 24946 10782
rect 28366 10834 28418 10846
rect 28366 10770 28418 10782
rect 37102 10834 37154 10846
rect 37102 10770 37154 10782
rect 37438 10834 37490 10846
rect 37438 10770 37490 10782
rect 39342 10834 39394 10846
rect 39342 10770 39394 10782
rect 41582 10834 41634 10846
rect 41582 10770 41634 10782
rect 42478 10834 42530 10846
rect 42478 10770 42530 10782
rect 42926 10834 42978 10846
rect 42926 10770 42978 10782
rect 43262 10834 43314 10846
rect 43262 10770 43314 10782
rect 43822 10834 43874 10846
rect 43822 10770 43874 10782
rect 44494 10834 44546 10846
rect 44494 10770 44546 10782
rect 45054 10834 45106 10846
rect 45054 10770 45106 10782
rect 46062 10834 46114 10846
rect 46062 10770 46114 10782
rect 47182 10834 47234 10846
rect 47182 10770 47234 10782
rect 47742 10834 47794 10846
rect 47742 10770 47794 10782
rect 48078 10834 48130 10846
rect 48078 10770 48130 10782
rect 48638 10834 48690 10846
rect 48638 10770 48690 10782
rect 49534 10834 49586 10846
rect 49534 10770 49586 10782
rect 50318 10834 50370 10846
rect 50318 10770 50370 10782
rect 51214 10834 51266 10846
rect 51214 10770 51266 10782
rect 51774 10834 51826 10846
rect 51774 10770 51826 10782
rect 53566 10834 53618 10846
rect 53566 10770 53618 10782
rect 54126 10834 54178 10846
rect 54126 10770 54178 10782
rect 54574 10834 54626 10846
rect 54574 10770 54626 10782
rect 55134 10834 55186 10846
rect 55134 10770 55186 10782
rect 55694 10834 55746 10846
rect 55694 10770 55746 10782
rect 56478 10834 56530 10846
rect 56478 10770 56530 10782
rect 57374 10834 57426 10846
rect 57374 10770 57426 10782
rect 57822 10834 57874 10846
rect 57822 10770 57874 10782
rect 2718 10722 2770 10734
rect 2718 10658 2770 10670
rect 15934 10722 15986 10734
rect 15934 10658 15986 10670
rect 16830 10722 16882 10734
rect 16830 10658 16882 10670
rect 18062 10722 18114 10734
rect 18062 10658 18114 10670
rect 19182 10722 19234 10734
rect 19182 10658 19234 10670
rect 19518 10722 19570 10734
rect 19518 10658 19570 10670
rect 23998 10722 24050 10734
rect 23998 10658 24050 10670
rect 30494 10722 30546 10734
rect 35758 10722 35810 10734
rect 32050 10670 32062 10722
rect 32114 10670 32126 10722
rect 30494 10658 30546 10670
rect 35758 10658 35810 10670
rect 36094 10722 36146 10734
rect 36094 10658 36146 10670
rect 37662 10722 37714 10734
rect 37662 10658 37714 10670
rect 38670 10722 38722 10734
rect 38670 10658 38722 10670
rect 44942 10722 44994 10734
rect 44942 10658 44994 10670
rect 50206 10722 50258 10734
rect 50206 10658 50258 10670
rect 50542 10722 50594 10734
rect 50542 10658 50594 10670
rect 51102 10722 51154 10734
rect 51102 10658 51154 10670
rect 52782 10722 52834 10734
rect 52782 10658 52834 10670
rect 52894 10722 52946 10734
rect 52894 10658 52946 10670
rect 53342 10722 53394 10734
rect 53342 10658 53394 10670
rect 53678 10722 53730 10734
rect 53678 10658 53730 10670
rect 16158 10610 16210 10622
rect 15586 10558 15598 10610
rect 15650 10558 15662 10610
rect 16158 10546 16210 10558
rect 16942 10610 16994 10622
rect 16942 10546 16994 10558
rect 17726 10610 17778 10622
rect 17726 10546 17778 10558
rect 18286 10610 18338 10622
rect 18286 10546 18338 10558
rect 19630 10610 19682 10622
rect 19630 10546 19682 10558
rect 22542 10610 22594 10622
rect 27582 10610 27634 10622
rect 31390 10610 31442 10622
rect 24322 10558 24334 10610
rect 24386 10558 24398 10610
rect 25890 10558 25902 10610
rect 25954 10558 25966 10610
rect 26114 10558 26126 10610
rect 26178 10558 26190 10610
rect 29138 10558 29150 10610
rect 29202 10558 29214 10610
rect 29362 10558 29374 10610
rect 29426 10558 29438 10610
rect 31154 10558 31166 10610
rect 31218 10558 31230 10610
rect 22542 10546 22594 10558
rect 27582 10546 27634 10558
rect 31390 10546 31442 10558
rect 32398 10610 32450 10622
rect 32398 10546 32450 10558
rect 34302 10610 34354 10622
rect 34302 10546 34354 10558
rect 34638 10610 34690 10622
rect 34638 10546 34690 10558
rect 34750 10610 34802 10622
rect 34750 10546 34802 10558
rect 37774 10610 37826 10622
rect 39454 10610 39506 10622
rect 38434 10558 38446 10610
rect 38498 10558 38510 10610
rect 37774 10546 37826 10558
rect 39454 10546 39506 10558
rect 40014 10610 40066 10622
rect 40014 10546 40066 10558
rect 40238 10610 40290 10622
rect 40238 10546 40290 10558
rect 50094 10610 50146 10622
rect 50094 10546 50146 10558
rect 15038 10498 15090 10510
rect 15038 10434 15090 10446
rect 16046 10498 16098 10510
rect 16046 10434 16098 10446
rect 19294 10498 19346 10510
rect 25678 10498 25730 10510
rect 22866 10446 22878 10498
rect 22930 10446 22942 10498
rect 19294 10434 19346 10446
rect 25678 10434 25730 10446
rect 27806 10498 27858 10510
rect 32846 10498 32898 10510
rect 28914 10446 28926 10498
rect 28978 10446 28990 10498
rect 27806 10434 27858 10446
rect 32846 10434 32898 10446
rect 33742 10498 33794 10510
rect 33742 10434 33794 10446
rect 34414 10498 34466 10510
rect 34414 10434 34466 10446
rect 36542 10498 36594 10510
rect 36542 10434 36594 10446
rect 41918 10498 41970 10510
rect 41918 10434 41970 10446
rect 45726 10498 45778 10510
rect 45726 10434 45778 10446
rect 46734 10498 46786 10510
rect 46734 10434 46786 10446
rect 56030 10498 56082 10510
rect 56030 10434 56082 10446
rect 14702 10386 14754 10398
rect 39342 10386 39394 10398
rect 45054 10386 45106 10398
rect 22978 10334 22990 10386
rect 23042 10334 23054 10386
rect 27234 10334 27246 10386
rect 27298 10334 27310 10386
rect 36306 10334 36318 10386
rect 36370 10383 36382 10386
rect 36866 10383 36878 10386
rect 36370 10337 36878 10383
rect 36370 10334 36382 10337
rect 36866 10334 36878 10337
rect 36930 10334 36942 10386
rect 40562 10334 40574 10386
rect 40626 10334 40638 10386
rect 14702 10322 14754 10334
rect 39342 10322 39394 10334
rect 45054 10322 45106 10334
rect 51214 10386 51266 10398
rect 51214 10322 51266 10334
rect 52782 10386 52834 10398
rect 57362 10334 57374 10386
rect 57426 10383 57438 10386
rect 57922 10383 57934 10386
rect 57426 10337 57934 10383
rect 57426 10334 57438 10337
rect 57922 10334 57934 10337
rect 57986 10334 57998 10386
rect 52782 10322 52834 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 17502 10050 17554 10062
rect 17502 9986 17554 9998
rect 17838 10050 17890 10062
rect 17838 9986 17890 9998
rect 26350 10050 26402 10062
rect 33182 10050 33234 10062
rect 32162 9998 32174 10050
rect 32226 10047 32238 10050
rect 32386 10047 32398 10050
rect 32226 10001 32398 10047
rect 32226 9998 32238 10001
rect 32386 9998 32398 10001
rect 32450 10047 32462 10050
rect 32834 10047 32846 10050
rect 32450 10001 32846 10047
rect 32450 9998 32462 10001
rect 32834 9998 32846 10001
rect 32898 9998 32910 10050
rect 26350 9986 26402 9998
rect 33182 9986 33234 9998
rect 33406 10050 33458 10062
rect 33406 9986 33458 9998
rect 33966 10050 34018 10062
rect 33966 9986 34018 9998
rect 44718 10050 44770 10062
rect 51550 10050 51602 10062
rect 48066 9998 48078 10050
rect 48130 10047 48142 10050
rect 48514 10047 48526 10050
rect 48130 10001 48526 10047
rect 48130 9998 48142 10001
rect 48514 9998 48526 10001
rect 48578 9998 48590 10050
rect 44718 9986 44770 9998
rect 51550 9986 51602 9998
rect 15598 9938 15650 9950
rect 21534 9938 21586 9950
rect 14578 9886 14590 9938
rect 14642 9886 14654 9938
rect 16482 9886 16494 9938
rect 16546 9886 16558 9938
rect 15598 9874 15650 9886
rect 21534 9874 21586 9886
rect 23102 9938 23154 9950
rect 23102 9874 23154 9886
rect 28814 9938 28866 9950
rect 28814 9874 28866 9886
rect 34750 9938 34802 9950
rect 34750 9874 34802 9886
rect 34862 9938 34914 9950
rect 34862 9874 34914 9886
rect 35534 9938 35586 9950
rect 35534 9874 35586 9886
rect 35758 9938 35810 9950
rect 35758 9874 35810 9886
rect 37886 9938 37938 9950
rect 41918 9938 41970 9950
rect 38322 9886 38334 9938
rect 38386 9886 38398 9938
rect 37886 9874 37938 9886
rect 41918 9874 41970 9886
rect 45390 9938 45442 9950
rect 45390 9874 45442 9886
rect 46174 9938 46226 9950
rect 46174 9874 46226 9886
rect 46510 9938 46562 9950
rect 46510 9874 46562 9886
rect 48526 9938 48578 9950
rect 48526 9874 48578 9886
rect 49086 9938 49138 9950
rect 49086 9874 49138 9886
rect 49646 9938 49698 9950
rect 52558 9938 52610 9950
rect 50306 9886 50318 9938
rect 50370 9886 50382 9938
rect 49646 9874 49698 9886
rect 52558 9874 52610 9886
rect 53790 9938 53842 9950
rect 53790 9874 53842 9886
rect 54686 9938 54738 9950
rect 54686 9874 54738 9886
rect 55246 9938 55298 9950
rect 55246 9874 55298 9886
rect 55582 9938 55634 9950
rect 55582 9874 55634 9886
rect 57038 9938 57090 9950
rect 57038 9874 57090 9886
rect 57374 9938 57426 9950
rect 57374 9874 57426 9886
rect 24110 9826 24162 9838
rect 14690 9774 14702 9826
rect 14754 9774 14766 9826
rect 16258 9774 16270 9826
rect 16322 9774 16334 9826
rect 24110 9762 24162 9774
rect 25230 9826 25282 9838
rect 29486 9826 29538 9838
rect 26002 9774 26014 9826
rect 26066 9774 26078 9826
rect 25230 9762 25282 9774
rect 29486 9762 29538 9774
rect 29822 9826 29874 9838
rect 29822 9762 29874 9774
rect 30046 9826 30098 9838
rect 30046 9762 30098 9774
rect 33854 9826 33906 9838
rect 33854 9762 33906 9774
rect 36766 9826 36818 9838
rect 40014 9826 40066 9838
rect 42142 9826 42194 9838
rect 38546 9774 38558 9826
rect 38610 9774 38622 9826
rect 40674 9774 40686 9826
rect 40738 9774 40750 9826
rect 41458 9774 41470 9826
rect 41522 9774 41534 9826
rect 36766 9762 36818 9774
rect 40014 9762 40066 9774
rect 42142 9762 42194 9774
rect 42814 9826 42866 9838
rect 53342 9826 53394 9838
rect 47506 9774 47518 9826
rect 47570 9774 47582 9826
rect 50194 9774 50206 9826
rect 50258 9774 50270 9826
rect 42814 9762 42866 9774
rect 53342 9762 53394 9774
rect 58046 9826 58098 9838
rect 58046 9762 58098 9774
rect 2382 9714 2434 9726
rect 2382 9650 2434 9662
rect 2718 9714 2770 9726
rect 2718 9650 2770 9662
rect 3278 9714 3330 9726
rect 3278 9650 3330 9662
rect 13806 9714 13858 9726
rect 13806 9650 13858 9662
rect 17614 9714 17666 9726
rect 17614 9650 17666 9662
rect 22990 9714 23042 9726
rect 22990 9650 23042 9662
rect 23214 9714 23266 9726
rect 23214 9650 23266 9662
rect 25790 9714 25842 9726
rect 25790 9650 25842 9662
rect 36094 9714 36146 9726
rect 36094 9650 36146 9662
rect 36318 9714 36370 9726
rect 36318 9650 36370 9662
rect 39902 9714 39954 9726
rect 42702 9714 42754 9726
rect 40226 9662 40238 9714
rect 40290 9662 40302 9714
rect 42466 9662 42478 9714
rect 42530 9662 42542 9714
rect 39902 9650 39954 9662
rect 42702 9650 42754 9662
rect 43822 9714 43874 9726
rect 43822 9650 43874 9662
rect 51326 9714 51378 9726
rect 51326 9650 51378 9662
rect 52110 9714 52162 9726
rect 52110 9650 52162 9662
rect 54350 9714 54402 9726
rect 54350 9650 54402 9662
rect 23774 9602 23826 9614
rect 23774 9538 23826 9550
rect 24894 9602 24946 9614
rect 24894 9538 24946 9550
rect 26238 9602 26290 9614
rect 26238 9538 26290 9550
rect 26686 9602 26738 9614
rect 26686 9538 26738 9550
rect 27134 9602 27186 9614
rect 27134 9538 27186 9550
rect 29822 9602 29874 9614
rect 29822 9538 29874 9550
rect 30606 9602 30658 9614
rect 30606 9538 30658 9550
rect 32510 9602 32562 9614
rect 32510 9538 32562 9550
rect 33070 9602 33122 9614
rect 33070 9538 33122 9550
rect 35422 9602 35474 9614
rect 35422 9538 35474 9550
rect 39342 9602 39394 9614
rect 39342 9538 39394 9550
rect 43486 9602 43538 9614
rect 43486 9538 43538 9550
rect 44494 9602 44546 9614
rect 44494 9538 44546 9550
rect 44606 9602 44658 9614
rect 44606 9538 44658 9550
rect 47294 9602 47346 9614
rect 47294 9538 47346 9550
rect 48190 9602 48242 9614
rect 48190 9538 48242 9550
rect 51438 9602 51490 9614
rect 51438 9538 51490 9550
rect 56030 9602 56082 9614
rect 56030 9538 56082 9550
rect 56478 9602 56530 9614
rect 56478 9538 56530 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 21982 9266 22034 9278
rect 21982 9202 22034 9214
rect 25006 9266 25058 9278
rect 25006 9202 25058 9214
rect 25678 9266 25730 9278
rect 25678 9202 25730 9214
rect 27470 9266 27522 9278
rect 27470 9202 27522 9214
rect 29038 9266 29090 9278
rect 32846 9266 32898 9278
rect 31602 9214 31614 9266
rect 31666 9214 31678 9266
rect 29038 9202 29090 9214
rect 32846 9202 32898 9214
rect 35982 9266 36034 9278
rect 35982 9202 36034 9214
rect 36206 9266 36258 9278
rect 36206 9202 36258 9214
rect 37214 9266 37266 9278
rect 37214 9202 37266 9214
rect 38446 9266 38498 9278
rect 38446 9202 38498 9214
rect 39230 9266 39282 9278
rect 39230 9202 39282 9214
rect 40350 9266 40402 9278
rect 40350 9202 40402 9214
rect 40910 9266 40962 9278
rect 46062 9266 46114 9278
rect 41682 9214 41694 9266
rect 41746 9214 41758 9266
rect 40910 9202 40962 9214
rect 46062 9202 46114 9214
rect 46510 9266 46562 9278
rect 48638 9266 48690 9278
rect 47282 9214 47294 9266
rect 47346 9214 47358 9266
rect 46510 9202 46562 9214
rect 48638 9202 48690 9214
rect 51886 9266 51938 9278
rect 51886 9202 51938 9214
rect 55582 9266 55634 9278
rect 55582 9202 55634 9214
rect 56030 9266 56082 9278
rect 56030 9202 56082 9214
rect 56478 9266 56530 9278
rect 56478 9202 56530 9214
rect 57374 9266 57426 9278
rect 57374 9202 57426 9214
rect 58046 9266 58098 9278
rect 58046 9202 58098 9214
rect 12686 9154 12738 9166
rect 12686 9090 12738 9102
rect 13022 9154 13074 9166
rect 13022 9090 13074 9102
rect 26686 9154 26738 9166
rect 26686 9090 26738 9102
rect 26910 9154 26962 9166
rect 34974 9154 35026 9166
rect 29810 9102 29822 9154
rect 29874 9102 29886 9154
rect 31378 9102 31390 9154
rect 31442 9102 31454 9154
rect 26910 9090 26962 9102
rect 34974 9090 35026 9102
rect 35198 9154 35250 9166
rect 35198 9090 35250 9102
rect 35534 9154 35586 9166
rect 35534 9090 35586 9102
rect 39342 9154 39394 9166
rect 39342 9090 39394 9102
rect 39678 9154 39730 9166
rect 39678 9090 39730 9102
rect 42478 9154 42530 9166
rect 47742 9154 47794 9166
rect 42914 9102 42926 9154
rect 42978 9102 42990 9154
rect 43362 9102 43374 9154
rect 43426 9102 43438 9154
rect 42478 9090 42530 9102
rect 47742 9090 47794 9102
rect 33742 9042 33794 9054
rect 19618 8990 19630 9042
rect 19682 8990 19694 9042
rect 21074 8990 21086 9042
rect 21138 8990 21150 9042
rect 25890 8990 25902 9042
rect 25954 8990 25966 9042
rect 26114 8990 26126 9042
rect 26178 8990 26190 9042
rect 30146 8990 30158 9042
rect 30210 8990 30222 9042
rect 33742 8978 33794 8990
rect 33966 9042 34018 9054
rect 33966 8978 34018 8990
rect 34190 9042 34242 9054
rect 36318 9042 36370 9054
rect 34402 8990 34414 9042
rect 34466 8990 34478 9042
rect 34190 8978 34242 8990
rect 36318 8978 36370 8990
rect 38222 9042 38274 9054
rect 38222 8978 38274 8990
rect 38334 9042 38386 9054
rect 38334 8978 38386 8990
rect 38782 9042 38834 9054
rect 38782 8978 38834 8990
rect 39454 9042 39506 9054
rect 39454 8978 39506 8990
rect 42030 9042 42082 9054
rect 44718 9042 44770 9054
rect 47854 9042 47906 9054
rect 43586 8990 43598 9042
rect 43650 8990 43662 9042
rect 45042 8990 45054 9042
rect 45106 8990 45118 9042
rect 42030 8978 42082 8990
rect 44718 8978 44770 8990
rect 47854 8978 47906 8990
rect 47966 9042 48018 9054
rect 50766 9042 50818 9054
rect 50306 8990 50318 9042
rect 50370 8990 50382 9042
rect 47966 8978 48018 8990
rect 50766 8978 50818 8990
rect 51438 9042 51490 9054
rect 55022 9042 55074 9054
rect 52882 8990 52894 9042
rect 52946 8990 52958 9042
rect 54450 8990 54462 9042
rect 54514 8990 54526 9042
rect 51438 8978 51490 8990
rect 55022 8978 55074 8990
rect 22542 8930 22594 8942
rect 20626 8878 20638 8930
rect 20690 8878 20702 8930
rect 22542 8866 22594 8878
rect 22990 8930 23042 8942
rect 32174 8930 32226 8942
rect 25778 8878 25790 8930
rect 25842 8878 25854 8930
rect 26898 8878 26910 8930
rect 26962 8878 26974 8930
rect 22990 8866 23042 8878
rect 32174 8866 32226 8878
rect 35422 8930 35474 8942
rect 35422 8866 35474 8878
rect 36766 8930 36818 8942
rect 36766 8866 36818 8878
rect 45614 8930 45666 8942
rect 45614 8866 45666 8878
rect 49870 8930 49922 8942
rect 53566 8930 53618 8942
rect 52658 8878 52670 8930
rect 52722 8878 52734 8930
rect 49870 8866 49922 8878
rect 53566 8866 53618 8878
rect 55134 8930 55186 8942
rect 55134 8866 55186 8878
rect 33630 8818 33682 8830
rect 19506 8766 19518 8818
rect 19570 8766 19582 8818
rect 33630 8754 33682 8766
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 21982 8482 22034 8494
rect 36542 8482 36594 8494
rect 16482 8430 16494 8482
rect 16546 8430 16558 8482
rect 25666 8430 25678 8482
rect 25730 8479 25742 8482
rect 25890 8479 25902 8482
rect 25730 8433 25902 8479
rect 25730 8430 25742 8433
rect 25890 8430 25902 8433
rect 25954 8430 25966 8482
rect 21982 8418 22034 8430
rect 36542 8418 36594 8430
rect 42926 8482 42978 8494
rect 42926 8418 42978 8430
rect 43598 8482 43650 8494
rect 43598 8418 43650 8430
rect 19630 8370 19682 8382
rect 17154 8318 17166 8370
rect 17218 8318 17230 8370
rect 19630 8306 19682 8318
rect 20414 8370 20466 8382
rect 20414 8306 20466 8318
rect 22766 8370 22818 8382
rect 22766 8306 22818 8318
rect 23550 8370 23602 8382
rect 23550 8306 23602 8318
rect 24446 8370 24498 8382
rect 24446 8306 24498 8318
rect 25342 8370 25394 8382
rect 31166 8370 31218 8382
rect 27010 8318 27022 8370
rect 27074 8318 27086 8370
rect 30482 8318 30494 8370
rect 30546 8318 30558 8370
rect 25342 8306 25394 8318
rect 31166 8306 31218 8318
rect 33294 8370 33346 8382
rect 33294 8306 33346 8318
rect 34638 8370 34690 8382
rect 34638 8306 34690 8318
rect 36430 8370 36482 8382
rect 36430 8306 36482 8318
rect 39230 8370 39282 8382
rect 39230 8306 39282 8318
rect 42142 8370 42194 8382
rect 42142 8306 42194 8318
rect 43150 8370 43202 8382
rect 48526 8370 48578 8382
rect 48066 8318 48078 8370
rect 48130 8318 48142 8370
rect 43150 8306 43202 8318
rect 48526 8306 48578 8318
rect 48974 8370 49026 8382
rect 48974 8306 49026 8318
rect 49534 8370 49586 8382
rect 49534 8306 49586 8318
rect 49870 8370 49922 8382
rect 56366 8370 56418 8382
rect 53778 8318 53790 8370
rect 53842 8318 53854 8370
rect 49870 8306 49922 8318
rect 56366 8306 56418 8318
rect 57486 8370 57538 8382
rect 57486 8306 57538 8318
rect 58046 8370 58098 8382
rect 58046 8306 58098 8318
rect 18510 8258 18562 8270
rect 20638 8258 20690 8270
rect 17266 8206 17278 8258
rect 17330 8206 17342 8258
rect 18610 8206 18622 8258
rect 18674 8206 18686 8258
rect 18510 8194 18562 8206
rect 20638 8194 20690 8206
rect 25006 8258 25058 8270
rect 25006 8194 25058 8206
rect 25118 8258 25170 8270
rect 25118 8194 25170 8206
rect 25566 8258 25618 8270
rect 25566 8194 25618 8206
rect 25902 8258 25954 8270
rect 25902 8194 25954 8206
rect 26574 8258 26626 8270
rect 28030 8258 28082 8270
rect 37550 8258 37602 8270
rect 26898 8206 26910 8258
rect 26962 8206 26974 8258
rect 30034 8206 30046 8258
rect 30098 8206 30110 8258
rect 34178 8206 34190 8258
rect 34242 8206 34254 8258
rect 34962 8206 34974 8258
rect 35026 8206 35038 8258
rect 26574 8194 26626 8206
rect 28030 8194 28082 8206
rect 37550 8194 37602 8206
rect 39006 8258 39058 8270
rect 39006 8194 39058 8206
rect 40910 8258 40962 8270
rect 40910 8194 40962 8206
rect 41134 8258 41186 8270
rect 41134 8194 41186 8206
rect 41358 8258 41410 8270
rect 41358 8194 41410 8206
rect 42702 8258 42754 8270
rect 42702 8194 42754 8206
rect 44046 8258 44098 8270
rect 44046 8194 44098 8206
rect 45502 8258 45554 8270
rect 47742 8258 47794 8270
rect 45826 8206 45838 8258
rect 45890 8206 45902 8258
rect 45502 8194 45554 8206
rect 47742 8194 47794 8206
rect 51998 8258 52050 8270
rect 51998 8194 52050 8206
rect 52446 8258 52498 8270
rect 54574 8258 54626 8270
rect 53666 8206 53678 8258
rect 53730 8206 53742 8258
rect 52446 8194 52498 8206
rect 54574 8194 54626 8206
rect 55134 8258 55186 8270
rect 55134 8194 55186 8206
rect 18062 8146 18114 8158
rect 22206 8146 22258 8158
rect 18274 8094 18286 8146
rect 18338 8094 18350 8146
rect 18062 8082 18114 8094
rect 22206 8082 22258 8094
rect 23774 8146 23826 8158
rect 23774 8082 23826 8094
rect 27694 8146 27746 8158
rect 27694 8082 27746 8094
rect 27806 8146 27858 8158
rect 27806 8082 27858 8094
rect 29598 8146 29650 8158
rect 29598 8082 29650 8094
rect 33070 8146 33122 8158
rect 38782 8146 38834 8158
rect 34626 8094 34638 8146
rect 34690 8094 34702 8146
rect 35074 8094 35086 8146
rect 35138 8094 35150 8146
rect 33070 8082 33122 8094
rect 38782 8082 38834 8094
rect 39342 8146 39394 8158
rect 39342 8082 39394 8094
rect 41582 8146 41634 8158
rect 41582 8082 41634 8094
rect 46734 8146 46786 8158
rect 46734 8082 46786 8094
rect 50990 8146 51042 8158
rect 50990 8082 51042 8094
rect 51662 8146 51714 8158
rect 51662 8082 51714 8094
rect 52558 8146 52610 8158
rect 52558 8082 52610 8094
rect 18846 8034 18898 8046
rect 27134 8034 27186 8046
rect 20066 7982 20078 8034
rect 20130 7982 20142 8034
rect 21634 7982 21646 8034
rect 21698 7982 21710 8034
rect 23202 7982 23214 8034
rect 23266 7982 23278 8034
rect 18846 7970 18898 7982
rect 27134 7970 27186 7982
rect 28478 8034 28530 8046
rect 28478 7970 28530 7982
rect 33182 8034 33234 8046
rect 33182 7970 33234 7982
rect 35982 8034 36034 8046
rect 39902 8034 39954 8046
rect 37874 7982 37886 8034
rect 37938 7982 37950 8034
rect 35982 7970 36034 7982
rect 39902 7970 39954 7982
rect 44382 8034 44434 8046
rect 44382 7970 44434 7982
rect 45614 8034 45666 8046
rect 45614 7970 45666 7982
rect 46958 8034 47010 8046
rect 46958 7970 47010 7982
rect 47070 8034 47122 8046
rect 47070 7970 47122 7982
rect 47182 8034 47234 8046
rect 47182 7970 47234 7982
rect 47966 8034 48018 8046
rect 47966 7970 48018 7982
rect 50318 8034 50370 8046
rect 50318 7970 50370 7982
rect 51774 8034 51826 8046
rect 51774 7970 51826 7982
rect 52782 8034 52834 8046
rect 52782 7970 52834 7982
rect 55246 8034 55298 8046
rect 55246 7970 55298 7982
rect 55470 8034 55522 8046
rect 55470 7970 55522 7982
rect 55806 8034 55858 8046
rect 55806 7970 55858 7982
rect 56926 8034 56978 8046
rect 56926 7970 56978 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 20414 7698 20466 7710
rect 20414 7634 20466 7646
rect 31614 7698 31666 7710
rect 31614 7634 31666 7646
rect 36990 7698 37042 7710
rect 36990 7634 37042 7646
rect 37886 7698 37938 7710
rect 37886 7634 37938 7646
rect 38334 7698 38386 7710
rect 38334 7634 38386 7646
rect 42478 7698 42530 7710
rect 42478 7634 42530 7646
rect 42702 7698 42754 7710
rect 42702 7634 42754 7646
rect 42814 7698 42866 7710
rect 42814 7634 42866 7646
rect 43822 7698 43874 7710
rect 43822 7634 43874 7646
rect 44382 7698 44434 7710
rect 44382 7634 44434 7646
rect 45054 7698 45106 7710
rect 45054 7634 45106 7646
rect 47518 7698 47570 7710
rect 47518 7634 47570 7646
rect 48190 7698 48242 7710
rect 48190 7634 48242 7646
rect 50654 7698 50706 7710
rect 50654 7634 50706 7646
rect 51662 7698 51714 7710
rect 51662 7634 51714 7646
rect 54350 7698 54402 7710
rect 54350 7634 54402 7646
rect 56814 7698 56866 7710
rect 56814 7634 56866 7646
rect 57598 7698 57650 7710
rect 57598 7634 57650 7646
rect 58046 7698 58098 7710
rect 58046 7634 58098 7646
rect 17726 7586 17778 7598
rect 17726 7522 17778 7534
rect 18062 7586 18114 7598
rect 18062 7522 18114 7534
rect 18286 7586 18338 7598
rect 18286 7522 18338 7534
rect 20078 7586 20130 7598
rect 20078 7522 20130 7534
rect 20302 7586 20354 7598
rect 20302 7522 20354 7534
rect 24894 7586 24946 7598
rect 24894 7522 24946 7534
rect 28478 7586 28530 7598
rect 28478 7522 28530 7534
rect 29374 7586 29426 7598
rect 29374 7522 29426 7534
rect 36206 7586 36258 7598
rect 36206 7522 36258 7534
rect 36542 7586 36594 7598
rect 36542 7522 36594 7534
rect 43486 7586 43538 7598
rect 43486 7522 43538 7534
rect 45502 7586 45554 7598
rect 45502 7522 45554 7534
rect 45726 7586 45778 7598
rect 45726 7522 45778 7534
rect 48414 7586 48466 7598
rect 48414 7522 48466 7534
rect 49646 7586 49698 7598
rect 49646 7522 49698 7534
rect 49758 7586 49810 7598
rect 52770 7534 52782 7586
rect 52834 7534 52846 7586
rect 49758 7522 49810 7534
rect 20750 7474 20802 7486
rect 23886 7474 23938 7486
rect 25678 7474 25730 7486
rect 22082 7422 22094 7474
rect 22146 7422 22158 7474
rect 23426 7422 23438 7474
rect 23490 7422 23502 7474
rect 24546 7422 24558 7474
rect 24610 7422 24622 7474
rect 20750 7410 20802 7422
rect 23886 7410 23938 7422
rect 25678 7410 25730 7422
rect 26574 7474 26626 7486
rect 31726 7474 31778 7486
rect 27010 7422 27022 7474
rect 27074 7422 27086 7474
rect 28130 7422 28142 7474
rect 28194 7422 28206 7474
rect 29026 7422 29038 7474
rect 29090 7422 29102 7474
rect 26574 7410 26626 7422
rect 31726 7410 31778 7422
rect 31950 7474 32002 7486
rect 35198 7474 35250 7486
rect 42926 7474 42978 7486
rect 32162 7422 32174 7474
rect 32226 7422 32238 7474
rect 35634 7422 35646 7474
rect 35698 7422 35710 7474
rect 31950 7410 32002 7422
rect 35198 7410 35250 7422
rect 42926 7410 42978 7422
rect 46174 7474 46226 7486
rect 46174 7410 46226 7422
rect 46622 7474 46674 7486
rect 46622 7410 46674 7422
rect 46846 7474 46898 7486
rect 46846 7410 46898 7422
rect 47854 7474 47906 7486
rect 53218 7422 53230 7474
rect 53282 7422 53294 7474
rect 53554 7422 53566 7474
rect 53618 7422 53630 7474
rect 56130 7422 56142 7474
rect 56194 7422 56206 7474
rect 47854 7410 47906 7422
rect 17838 7362 17890 7374
rect 17838 7298 17890 7310
rect 21422 7362 21474 7374
rect 22990 7362 23042 7374
rect 22306 7310 22318 7362
rect 22370 7310 22382 7362
rect 21422 7298 21474 7310
rect 22990 7298 23042 7310
rect 25790 7362 25842 7374
rect 25790 7298 25842 7310
rect 27470 7362 27522 7374
rect 29822 7362 29874 7374
rect 28242 7310 28254 7362
rect 28306 7310 28318 7362
rect 27470 7298 27522 7310
rect 29822 7298 29874 7310
rect 30942 7362 30994 7374
rect 30942 7298 30994 7310
rect 31838 7362 31890 7374
rect 31838 7298 31890 7310
rect 37438 7362 37490 7374
rect 37438 7298 37490 7310
rect 45950 7362 46002 7374
rect 45950 7298 46002 7310
rect 47070 7362 47122 7374
rect 47070 7298 47122 7310
rect 50206 7362 50258 7374
rect 50206 7298 50258 7310
rect 51102 7362 51154 7374
rect 51102 7298 51154 7310
rect 51998 7362 52050 7374
rect 52770 7310 52782 7362
rect 52834 7310 52846 7362
rect 55346 7310 55358 7362
rect 55410 7310 55422 7362
rect 51998 7298 52050 7310
rect 24558 7250 24610 7262
rect 24558 7186 24610 7198
rect 29038 7250 29090 7262
rect 29038 7186 29090 7198
rect 35086 7250 35138 7262
rect 35086 7186 35138 7198
rect 35422 7250 35474 7262
rect 35422 7186 35474 7198
rect 48526 7250 48578 7262
rect 48526 7186 48578 7198
rect 49646 7250 49698 7262
rect 49646 7186 49698 7198
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 41918 6914 41970 6926
rect 19170 6862 19182 6914
rect 19234 6862 19246 6914
rect 51314 6862 51326 6914
rect 51378 6862 51390 6914
rect 41918 6850 41970 6862
rect 20974 6802 21026 6814
rect 20974 6738 21026 6750
rect 21646 6802 21698 6814
rect 21646 6738 21698 6750
rect 28702 6802 28754 6814
rect 28702 6738 28754 6750
rect 33294 6802 33346 6814
rect 33294 6738 33346 6750
rect 42702 6802 42754 6814
rect 57822 6802 57874 6814
rect 49186 6750 49198 6802
rect 49250 6750 49262 6802
rect 42702 6738 42754 6750
rect 57822 6738 57874 6750
rect 19294 6690 19346 6702
rect 22878 6690 22930 6702
rect 19618 6638 19630 6690
rect 19682 6638 19694 6690
rect 19294 6626 19346 6638
rect 22878 6626 22930 6638
rect 23214 6690 23266 6702
rect 23214 6626 23266 6638
rect 23438 6690 23490 6702
rect 23438 6626 23490 6638
rect 23998 6690 24050 6702
rect 23998 6626 24050 6638
rect 24222 6690 24274 6702
rect 24222 6626 24274 6638
rect 24670 6690 24722 6702
rect 24670 6626 24722 6638
rect 27470 6690 27522 6702
rect 27470 6626 27522 6638
rect 28030 6690 28082 6702
rect 28030 6626 28082 6638
rect 30830 6690 30882 6702
rect 30830 6626 30882 6638
rect 31390 6690 31442 6702
rect 31390 6626 31442 6638
rect 31614 6690 31666 6702
rect 31614 6626 31666 6638
rect 32174 6690 32226 6702
rect 33070 6690 33122 6702
rect 32834 6638 32846 6690
rect 32898 6638 32910 6690
rect 32174 6626 32226 6638
rect 33070 6626 33122 6638
rect 34638 6690 34690 6702
rect 34638 6626 34690 6638
rect 35310 6690 35362 6702
rect 35310 6626 35362 6638
rect 35758 6690 35810 6702
rect 35758 6626 35810 6638
rect 36542 6690 36594 6702
rect 36542 6626 36594 6638
rect 38222 6690 38274 6702
rect 43598 6690 43650 6702
rect 38770 6638 38782 6690
rect 38834 6638 38846 6690
rect 38222 6626 38274 6638
rect 43598 6626 43650 6638
rect 45390 6690 45442 6702
rect 45390 6626 45442 6638
rect 46174 6690 46226 6702
rect 47966 6690 48018 6702
rect 46610 6638 46622 6690
rect 46674 6638 46686 6690
rect 46174 6626 46226 6638
rect 47966 6626 48018 6638
rect 48190 6690 48242 6702
rect 52558 6690 52610 6702
rect 49298 6638 49310 6690
rect 49362 6638 49374 6690
rect 50642 6638 50654 6690
rect 50706 6638 50718 6690
rect 48190 6626 48242 6638
rect 52558 6626 52610 6638
rect 53454 6690 53506 6702
rect 53454 6626 53506 6638
rect 53790 6690 53842 6702
rect 53790 6626 53842 6638
rect 54238 6690 54290 6702
rect 54238 6626 54290 6638
rect 54798 6690 54850 6702
rect 54798 6626 54850 6638
rect 55918 6690 55970 6702
rect 55918 6626 55970 6638
rect 56814 6690 56866 6702
rect 56814 6626 56866 6638
rect 2718 6578 2770 6590
rect 2718 6514 2770 6526
rect 27134 6578 27186 6590
rect 27134 6514 27186 6526
rect 28142 6578 28194 6590
rect 28142 6514 28194 6526
rect 30718 6578 30770 6590
rect 30718 6514 30770 6526
rect 31726 6578 31778 6590
rect 46062 6578 46114 6590
rect 36194 6526 36206 6578
rect 36258 6526 36270 6578
rect 31726 6514 31778 6526
rect 46062 6514 46114 6526
rect 48526 6578 48578 6590
rect 48526 6514 48578 6526
rect 55358 6578 55410 6590
rect 55358 6514 55410 6526
rect 56254 6578 56306 6590
rect 56254 6514 56306 6526
rect 2382 6466 2434 6478
rect 2382 6402 2434 6414
rect 3166 6466 3218 6478
rect 3166 6402 3218 6414
rect 22990 6466 23042 6478
rect 22990 6402 23042 6414
rect 24110 6466 24162 6478
rect 24110 6402 24162 6414
rect 29486 6466 29538 6478
rect 29486 6402 29538 6414
rect 30494 6466 30546 6478
rect 30494 6402 30546 6414
rect 32398 6466 32450 6478
rect 32398 6402 32450 6414
rect 32958 6466 33010 6478
rect 32958 6402 33010 6414
rect 33854 6466 33906 6478
rect 33854 6402 33906 6414
rect 35086 6466 35138 6478
rect 35086 6402 35138 6414
rect 35198 6466 35250 6478
rect 35198 6402 35250 6414
rect 37438 6466 37490 6478
rect 43038 6466 43090 6478
rect 41122 6414 41134 6466
rect 41186 6414 41198 6466
rect 37438 6402 37490 6414
rect 43038 6402 43090 6414
rect 44046 6466 44098 6478
rect 48078 6466 48130 6478
rect 44370 6414 44382 6466
rect 44434 6414 44446 6466
rect 44046 6402 44098 6414
rect 48078 6402 48130 6414
rect 51998 6466 52050 6478
rect 51998 6402 52050 6414
rect 57150 6466 57202 6478
rect 57150 6402 57202 6414
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 20638 6130 20690 6142
rect 20638 6066 20690 6078
rect 24558 6130 24610 6142
rect 24558 6066 24610 6078
rect 27582 6130 27634 6142
rect 42702 6130 42754 6142
rect 32498 6078 32510 6130
rect 32562 6078 32574 6130
rect 27582 6066 27634 6078
rect 42702 6066 42754 6078
rect 44494 6130 44546 6142
rect 44494 6066 44546 6078
rect 45278 6130 45330 6142
rect 45278 6066 45330 6078
rect 45390 6130 45442 6142
rect 45390 6066 45442 6078
rect 45950 6130 46002 6142
rect 45950 6066 46002 6078
rect 46510 6130 46562 6142
rect 46510 6066 46562 6078
rect 47182 6130 47234 6142
rect 47182 6066 47234 6078
rect 48078 6130 48130 6142
rect 48078 6066 48130 6078
rect 48414 6130 48466 6142
rect 48414 6066 48466 6078
rect 49758 6130 49810 6142
rect 49758 6066 49810 6078
rect 51326 6130 51378 6142
rect 51326 6066 51378 6078
rect 52446 6130 52498 6142
rect 52446 6066 52498 6078
rect 53342 6130 53394 6142
rect 53342 6066 53394 6078
rect 53790 6130 53842 6142
rect 53790 6066 53842 6078
rect 54462 6130 54514 6142
rect 54462 6066 54514 6078
rect 55918 6130 55970 6142
rect 55918 6066 55970 6078
rect 56366 6130 56418 6142
rect 56366 6066 56418 6078
rect 57934 6130 57986 6142
rect 57934 6066 57986 6078
rect 20414 6018 20466 6030
rect 20414 5954 20466 5966
rect 24334 6018 24386 6030
rect 24334 5954 24386 5966
rect 27246 6018 27298 6030
rect 40126 6018 40178 6030
rect 31154 5966 31166 6018
rect 31218 5966 31230 6018
rect 32610 5966 32622 6018
rect 32674 5966 32686 6018
rect 33618 5966 33630 6018
rect 33682 5966 33694 6018
rect 27246 5954 27298 5966
rect 40126 5954 40178 5966
rect 40910 6018 40962 6030
rect 40910 5954 40962 5966
rect 42814 6018 42866 6030
rect 43822 6018 43874 6030
rect 43474 5966 43486 6018
rect 43538 5966 43550 6018
rect 42814 5954 42866 5966
rect 43822 5954 43874 5966
rect 44382 6018 44434 6030
rect 44382 5954 44434 5966
rect 45502 6018 45554 6030
rect 45502 5954 45554 5966
rect 49870 6018 49922 6030
rect 49870 5954 49922 5966
rect 53006 6018 53058 6030
rect 53006 5954 53058 5966
rect 54910 6018 54962 6030
rect 54910 5954 54962 5966
rect 28366 5906 28418 5918
rect 2818 5854 2830 5906
rect 2882 5854 2894 5906
rect 22082 5854 22094 5906
rect 22146 5854 22158 5906
rect 28366 5842 28418 5854
rect 33966 5906 34018 5918
rect 33966 5842 34018 5854
rect 35758 5906 35810 5918
rect 35758 5842 35810 5854
rect 36206 5906 36258 5918
rect 36206 5842 36258 5854
rect 37214 5906 37266 5918
rect 57374 5906 57426 5918
rect 37874 5854 37886 5906
rect 37938 5854 37950 5906
rect 49522 5854 49534 5906
rect 49586 5854 49598 5906
rect 37214 5842 37266 5854
rect 57374 5842 57426 5854
rect 28142 5794 28194 5806
rect 34190 5794 34242 5806
rect 1922 5742 1934 5794
rect 1986 5742 1998 5794
rect 30706 5742 30718 5794
rect 30770 5742 30782 5794
rect 28142 5730 28194 5742
rect 34190 5730 34242 5742
rect 34638 5794 34690 5806
rect 34638 5730 34690 5742
rect 35310 5794 35362 5806
rect 35310 5730 35362 5742
rect 35982 5794 36034 5806
rect 35982 5730 36034 5742
rect 36654 5794 36706 5806
rect 36654 5730 36706 5742
rect 50318 5794 50370 5806
rect 50318 5730 50370 5742
rect 50878 5794 50930 5806
rect 50878 5730 50930 5742
rect 51774 5794 51826 5806
rect 51774 5730 51826 5742
rect 55246 5794 55298 5806
rect 55246 5730 55298 5742
rect 56814 5794 56866 5806
rect 56814 5730 56866 5742
rect 20750 5682 20802 5694
rect 20750 5618 20802 5630
rect 22094 5682 22146 5694
rect 22094 5618 22146 5630
rect 22430 5682 22482 5694
rect 22430 5618 22482 5630
rect 24670 5682 24722 5694
rect 24670 5618 24722 5630
rect 28702 5682 28754 5694
rect 28702 5618 28754 5630
rect 42590 5682 42642 5694
rect 50866 5630 50878 5682
rect 50930 5679 50942 5682
rect 51762 5679 51774 5682
rect 50930 5633 51774 5679
rect 50930 5630 50942 5633
rect 51762 5630 51774 5633
rect 51826 5630 51838 5682
rect 53890 5630 53902 5682
rect 53954 5679 53966 5682
rect 55234 5679 55246 5682
rect 53954 5633 55246 5679
rect 53954 5630 53966 5633
rect 55234 5630 55246 5633
rect 55298 5630 55310 5682
rect 56018 5630 56030 5682
rect 56082 5679 56094 5682
rect 56802 5679 56814 5682
rect 56082 5633 56814 5679
rect 56082 5630 56094 5633
rect 56802 5630 56814 5633
rect 56866 5630 56878 5682
rect 42590 5618 42642 5630
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 22094 5346 22146 5358
rect 22094 5282 22146 5294
rect 31502 5346 31554 5358
rect 47842 5294 47854 5346
rect 47906 5343 47918 5346
rect 49186 5343 49198 5346
rect 47906 5297 49198 5343
rect 47906 5294 47918 5297
rect 49186 5294 49198 5297
rect 49250 5294 49262 5346
rect 31502 5282 31554 5294
rect 21646 5234 21698 5246
rect 33742 5234 33794 5246
rect 28018 5182 28030 5234
rect 28082 5182 28094 5234
rect 31154 5182 31166 5234
rect 31218 5182 31230 5234
rect 21646 5170 21698 5182
rect 33742 5170 33794 5182
rect 36542 5234 36594 5246
rect 36542 5170 36594 5182
rect 43822 5234 43874 5246
rect 43822 5170 43874 5182
rect 45390 5234 45442 5246
rect 45390 5170 45442 5182
rect 46398 5234 46450 5246
rect 46398 5170 46450 5182
rect 46734 5234 46786 5246
rect 46734 5170 46786 5182
rect 47854 5234 47906 5246
rect 47854 5170 47906 5182
rect 48302 5234 48354 5246
rect 48302 5170 48354 5182
rect 48750 5234 48802 5246
rect 48750 5170 48802 5182
rect 49198 5234 49250 5246
rect 49198 5170 49250 5182
rect 50430 5234 50482 5246
rect 50430 5170 50482 5182
rect 50990 5234 51042 5246
rect 50990 5170 51042 5182
rect 51662 5234 51714 5246
rect 51662 5170 51714 5182
rect 52110 5234 52162 5246
rect 52110 5170 52162 5182
rect 52446 5234 52498 5246
rect 52446 5170 52498 5182
rect 53902 5234 53954 5246
rect 53902 5170 53954 5182
rect 54350 5234 54402 5246
rect 54350 5170 54402 5182
rect 54798 5234 54850 5246
rect 54798 5170 54850 5182
rect 55246 5234 55298 5246
rect 55246 5170 55298 5182
rect 55582 5234 55634 5246
rect 55582 5170 55634 5182
rect 20526 5122 20578 5134
rect 20526 5058 20578 5070
rect 20638 5122 20690 5134
rect 20638 5058 20690 5070
rect 21870 5122 21922 5134
rect 21870 5058 21922 5070
rect 24110 5122 24162 5134
rect 24110 5058 24162 5070
rect 24222 5122 24274 5134
rect 24222 5058 24274 5070
rect 24894 5122 24946 5134
rect 37774 5122 37826 5134
rect 28354 5070 28366 5122
rect 28418 5070 28430 5122
rect 32498 5070 32510 5122
rect 32562 5070 32574 5122
rect 32946 5070 32958 5122
rect 33010 5070 33022 5122
rect 24894 5058 24946 5070
rect 37774 5058 37826 5070
rect 38222 5122 38274 5134
rect 41918 5122 41970 5134
rect 38882 5070 38894 5122
rect 38946 5070 38958 5122
rect 38222 5058 38274 5070
rect 41918 5058 41970 5070
rect 49646 5122 49698 5134
rect 49646 5058 49698 5070
rect 20750 5010 20802 5022
rect 20750 4946 20802 4958
rect 23774 5010 23826 5022
rect 23774 4946 23826 4958
rect 23998 5010 24050 5022
rect 23998 4946 24050 4958
rect 25118 5010 25170 5022
rect 25118 4946 25170 4958
rect 25454 5010 25506 5022
rect 25454 4946 25506 4958
rect 28814 5010 28866 5022
rect 28814 4946 28866 4958
rect 31278 5010 31330 5022
rect 37662 5010 37714 5022
rect 32386 4958 32398 5010
rect 32450 4958 32462 5010
rect 34626 4958 34638 5010
rect 34690 4958 34702 5010
rect 31278 4946 31330 4958
rect 37662 4946 37714 4958
rect 47518 5010 47570 5022
rect 47518 4946 47570 4958
rect 22542 4898 22594 4910
rect 22542 4834 22594 4846
rect 23886 4898 23938 4910
rect 23886 4834 23938 4846
rect 25342 4898 25394 4910
rect 37438 4898 37490 4910
rect 32946 4846 32958 4898
rect 33010 4846 33022 4898
rect 41122 4846 41134 4898
rect 41186 4846 41198 4898
rect 25342 4834 25394 4846
rect 37438 4834 37490 4846
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 3278 4562 3330 4574
rect 3278 4498 3330 4510
rect 33518 4562 33570 4574
rect 37998 4562 38050 4574
rect 37426 4510 37438 4562
rect 37490 4510 37502 4562
rect 33518 4498 33570 4510
rect 37998 4498 38050 4510
rect 38446 4562 38498 4574
rect 46846 4562 46898 4574
rect 38770 4510 38782 4562
rect 38834 4510 38846 4562
rect 38446 4498 38498 4510
rect 46846 4498 46898 4510
rect 47294 4562 47346 4574
rect 47294 4498 47346 4510
rect 47742 4562 47794 4574
rect 47742 4498 47794 4510
rect 54350 4562 54402 4574
rect 54350 4498 54402 4510
rect 2382 4450 2434 4462
rect 2382 4386 2434 4398
rect 2718 4450 2770 4462
rect 2718 4386 2770 4398
rect 26350 4450 26402 4462
rect 26350 4386 26402 4398
rect 30606 4450 30658 4462
rect 30606 4386 30658 4398
rect 39342 4450 39394 4462
rect 39342 4386 39394 4398
rect 39454 4450 39506 4462
rect 39454 4386 39506 4398
rect 48526 4450 48578 4462
rect 48526 4386 48578 4398
rect 57486 4450 57538 4462
rect 57486 4386 57538 4398
rect 22430 4338 22482 4350
rect 26686 4338 26738 4350
rect 30270 4338 30322 4350
rect 21970 4286 21982 4338
rect 22034 4286 22046 4338
rect 23090 4286 23102 4338
rect 23154 4286 23166 4338
rect 28466 4286 28478 4338
rect 28530 4286 28542 4338
rect 29362 4286 29374 4338
rect 29426 4286 29438 4338
rect 22430 4274 22482 4286
rect 26686 4274 26738 4286
rect 30270 4274 30322 4286
rect 31838 4338 31890 4350
rect 34526 4338 34578 4350
rect 40014 4338 40066 4350
rect 56702 4338 56754 4350
rect 32386 4286 32398 4338
rect 32450 4286 32462 4338
rect 34962 4286 34974 4338
rect 35026 4286 35038 4338
rect 48290 4286 48302 4338
rect 48354 4286 48366 4338
rect 54898 4286 54910 4338
rect 54962 4286 54974 4338
rect 57698 4286 57710 4338
rect 57762 4286 57774 4338
rect 31838 4274 31890 4286
rect 34526 4274 34578 4286
rect 40014 4274 40066 4286
rect 56702 4274 56754 4286
rect 23874 4174 23886 4226
rect 23938 4174 23950 4226
rect 28578 4174 28590 4226
rect 28642 4174 28654 4226
rect 28914 4174 28926 4226
rect 28978 4174 28990 4226
rect 32610 4174 32622 4226
rect 32674 4174 32686 4226
rect 55794 4174 55806 4226
rect 55858 4174 55870 4226
rect 39454 4114 39506 4126
rect 39454 4050 39506 4062
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 19294 3666 19346 3678
rect 30270 3666 30322 3678
rect 6962 3614 6974 3666
rect 7026 3614 7038 3666
rect 27570 3614 27582 3666
rect 27634 3614 27646 3666
rect 29362 3614 29374 3666
rect 29426 3614 29438 3666
rect 19294 3602 19346 3614
rect 30270 3602 30322 3614
rect 33182 3666 33234 3678
rect 35646 3666 35698 3678
rect 34514 3614 34526 3666
rect 34578 3614 34590 3666
rect 33182 3602 33234 3614
rect 35646 3602 35698 3614
rect 37102 3666 37154 3678
rect 37102 3602 37154 3614
rect 37550 3666 37602 3678
rect 37550 3602 37602 3614
rect 37998 3666 38050 3678
rect 37998 3602 38050 3614
rect 38446 3666 38498 3678
rect 38446 3602 38498 3614
rect 47966 3666 48018 3678
rect 51314 3614 51326 3666
rect 51378 3614 51390 3666
rect 55234 3614 55246 3666
rect 55298 3614 55310 3666
rect 47966 3602 48018 3614
rect 26798 3554 26850 3566
rect 40910 3554 40962 3566
rect 2818 3502 2830 3554
rect 2882 3502 2894 3554
rect 12226 3502 12238 3554
rect 12290 3502 12302 3554
rect 18722 3502 18734 3554
rect 18786 3502 18798 3554
rect 23650 3502 23662 3554
rect 23714 3502 23726 3554
rect 28466 3502 28478 3554
rect 28530 3502 28542 3554
rect 29810 3502 29822 3554
rect 29874 3502 29886 3554
rect 33842 3502 33854 3554
rect 33906 3502 33918 3554
rect 40002 3502 40014 3554
rect 40066 3502 40078 3554
rect 26798 3490 26850 3502
rect 40910 3490 40962 3502
rect 44270 3554 44322 3566
rect 45154 3502 45166 3554
rect 45218 3502 45230 3554
rect 50642 3502 50654 3554
rect 50706 3502 50718 3554
rect 55906 3502 55918 3554
rect 55970 3502 55982 3554
rect 44270 3490 44322 3502
rect 5070 3442 5122 3454
rect 1922 3390 1934 3442
rect 1986 3390 1998 3442
rect 5842 3390 5854 3442
rect 5906 3390 5918 3442
rect 11106 3390 11118 3442
rect 11170 3390 11182 3442
rect 17602 3390 17614 3442
rect 17666 3390 17678 3442
rect 22530 3390 22542 3442
rect 22594 3390 22606 3442
rect 39106 3390 39118 3442
rect 39170 3390 39182 3442
rect 5070 3378 5122 3390
rect 44930 3278 44942 3330
rect 44994 3278 45006 3330
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 6750 56590 6802 56642
rect 7646 56590 7698 56642
rect 40350 56590 40402 56642
rect 41134 56590 41186 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 4622 56254 4674 56306
rect 16382 56254 16434 56306
rect 27470 56254 27522 56306
rect 31278 56254 31330 56306
rect 33630 56254 33682 56306
rect 38334 56254 38386 56306
rect 38782 56254 38834 56306
rect 39454 56254 39506 56306
rect 42814 56254 42866 56306
rect 2270 56142 2322 56194
rect 14142 56142 14194 56194
rect 22654 56142 22706 56194
rect 26126 56142 26178 56194
rect 26574 56142 26626 56194
rect 30270 56142 30322 56194
rect 35198 56142 35250 56194
rect 41134 56142 41186 56194
rect 43598 56142 43650 56194
rect 55806 56142 55858 56194
rect 7198 56030 7250 56082
rect 12798 56030 12850 56082
rect 17502 56030 17554 56082
rect 18510 56030 18562 56082
rect 22542 56030 22594 56082
rect 24446 56030 24498 56082
rect 25678 56030 25730 56082
rect 27918 56030 27970 56082
rect 28254 56030 28306 56082
rect 28478 56030 28530 56082
rect 34414 56030 34466 56082
rect 36094 56030 36146 56082
rect 39790 56030 39842 56082
rect 42254 56030 42306 56082
rect 46622 56030 46674 56082
rect 52782 56030 52834 56082
rect 54686 56030 54738 56082
rect 3054 55918 3106 55970
rect 4174 55918 4226 55970
rect 5070 55918 5122 55970
rect 6078 55918 6130 55970
rect 6526 55918 6578 55970
rect 7646 55918 7698 55970
rect 8990 55918 9042 55970
rect 9774 55918 9826 55970
rect 10222 55918 10274 55970
rect 10670 55918 10722 55970
rect 11118 55918 11170 55970
rect 12126 55918 12178 55970
rect 13694 55918 13746 55970
rect 14590 55918 14642 55970
rect 15038 55918 15090 55970
rect 15486 55918 15538 55970
rect 15934 55918 15986 55970
rect 16830 55918 16882 55970
rect 17950 55918 18002 55970
rect 19070 55918 19122 55970
rect 20190 55918 20242 55970
rect 20750 55918 20802 55970
rect 21310 55918 21362 55970
rect 22094 55918 22146 55970
rect 23550 55918 23602 55970
rect 25342 55918 25394 55970
rect 28366 55918 28418 55970
rect 29262 55918 29314 55970
rect 31614 55918 31666 55970
rect 32174 55918 32226 55970
rect 33182 55918 33234 55970
rect 33966 55918 34018 55970
rect 36990 55918 37042 55970
rect 37550 55918 37602 55970
rect 37998 55918 38050 55970
rect 40238 55918 40290 55970
rect 43150 55918 43202 55970
rect 46174 55918 46226 55970
rect 47294 55918 47346 55970
rect 53454 55918 53506 55970
rect 14366 55806 14418 55858
rect 15038 55806 15090 55858
rect 15822 55806 15874 55858
rect 16382 55806 16434 55858
rect 20190 55806 20242 55858
rect 20862 55806 20914 55858
rect 22654 55806 22706 55858
rect 30942 55806 30994 55858
rect 31614 55806 31666 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 20302 55470 20354 55522
rect 21086 55470 21138 55522
rect 30382 55470 30434 55522
rect 30942 55470 30994 55522
rect 53902 55470 53954 55522
rect 54686 55470 54738 55522
rect 1934 55358 1986 55410
rect 5854 55358 5906 55410
rect 12910 55358 12962 55410
rect 19854 55358 19906 55410
rect 20302 55358 20354 55410
rect 25790 55358 25842 55410
rect 28478 55358 28530 55410
rect 30606 55358 30658 55410
rect 32958 55358 33010 55410
rect 36542 55358 36594 55410
rect 37886 55358 37938 55410
rect 38894 55358 38946 55410
rect 44606 55358 44658 55410
rect 45838 55358 45890 55410
rect 56030 55358 56082 55410
rect 2830 55246 2882 55298
rect 7534 55246 7586 55298
rect 15038 55246 15090 55298
rect 15150 55246 15202 55298
rect 15262 55246 15314 55298
rect 19182 55246 19234 55298
rect 22094 55246 22146 55298
rect 24222 55246 24274 55298
rect 24894 55246 24946 55298
rect 25230 55246 25282 55298
rect 28030 55246 28082 55298
rect 28254 55246 28306 55298
rect 29934 55246 29986 55298
rect 34302 55246 34354 55298
rect 39342 55246 39394 55298
rect 40014 55246 40066 55298
rect 43150 55246 43202 55298
rect 43374 55246 43426 55298
rect 44046 55246 44098 55298
rect 44494 55246 44546 55298
rect 45726 55246 45778 55298
rect 54910 55246 54962 55298
rect 5070 55134 5122 55186
rect 7198 55134 7250 55186
rect 9438 55134 9490 55186
rect 12126 55134 12178 55186
rect 12574 55134 12626 55186
rect 14702 55134 14754 55186
rect 16270 55134 16322 55186
rect 16606 55134 16658 55186
rect 17166 55134 17218 55186
rect 17278 55134 17330 55186
rect 18174 55134 18226 55186
rect 23102 55134 23154 55186
rect 26238 55134 26290 55186
rect 30158 55134 30210 55186
rect 31166 55134 31218 55186
rect 35758 55134 35810 55186
rect 36094 55134 36146 55186
rect 38558 55134 38610 55186
rect 41134 55134 41186 55186
rect 42478 55134 42530 55186
rect 46622 55134 46674 55186
rect 47182 55134 47234 55186
rect 47518 55134 47570 55186
rect 3726 55022 3778 55074
rect 4174 55022 4226 55074
rect 4622 55022 4674 55074
rect 6302 55022 6354 55074
rect 6750 55022 6802 55074
rect 8094 55022 8146 55074
rect 8542 55022 8594 55074
rect 8878 55022 8930 55074
rect 9774 55022 9826 55074
rect 10670 55022 10722 55074
rect 11006 55022 11058 55074
rect 11678 55022 11730 55074
rect 13694 55022 13746 55074
rect 14142 55022 14194 55074
rect 15150 55022 15202 55074
rect 17502 55022 17554 55074
rect 18286 55022 18338 55074
rect 18398 55022 18450 55074
rect 19406 55022 19458 55074
rect 20862 55022 20914 55074
rect 22318 55022 22370 55074
rect 23214 55022 23266 55074
rect 23326 55022 23378 55074
rect 23998 55022 24050 55074
rect 25006 55022 25058 55074
rect 25678 55022 25730 55074
rect 26686 55022 26738 55074
rect 27134 55022 27186 55074
rect 28926 55022 28978 55074
rect 29710 55022 29762 55074
rect 30046 55022 30098 55074
rect 31390 55022 31442 55074
rect 31614 55022 31666 55074
rect 31726 55022 31778 55074
rect 32174 55022 32226 55074
rect 32622 55022 32674 55074
rect 33406 55022 33458 55074
rect 33966 55022 34018 55074
rect 34862 55022 34914 55074
rect 35198 55022 35250 55074
rect 37438 55022 37490 55074
rect 38782 55022 38834 55074
rect 39790 55022 39842 55074
rect 39902 55022 39954 55074
rect 40462 55022 40514 55074
rect 41246 55022 41298 55074
rect 41470 55022 41522 55074
rect 41918 55022 41970 55074
rect 44718 55022 44770 55074
rect 53902 55022 53954 55074
rect 54350 55022 54402 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 5182 54686 5234 54738
rect 7422 54686 7474 54738
rect 8654 54686 8706 54738
rect 13918 54686 13970 54738
rect 19070 54686 19122 54738
rect 20414 54686 20466 54738
rect 20526 54686 20578 54738
rect 22094 54686 22146 54738
rect 23550 54686 23602 54738
rect 23662 54686 23714 54738
rect 25790 54686 25842 54738
rect 26350 54686 26402 54738
rect 30718 54686 30770 54738
rect 30942 54686 30994 54738
rect 36206 54686 36258 54738
rect 36990 54686 37042 54738
rect 40798 54686 40850 54738
rect 45838 54686 45890 54738
rect 9886 54574 9938 54626
rect 10334 54574 10386 54626
rect 10446 54574 10498 54626
rect 12462 54574 12514 54626
rect 12798 54574 12850 54626
rect 14814 54574 14866 54626
rect 24446 54574 24498 54626
rect 24558 54574 24610 54626
rect 26574 54574 26626 54626
rect 26910 54574 26962 54626
rect 27694 54574 27746 54626
rect 27918 54574 27970 54626
rect 34414 54574 34466 54626
rect 37774 54574 37826 54626
rect 42926 54574 42978 54626
rect 43598 54574 43650 54626
rect 43710 54574 43762 54626
rect 44158 54574 44210 54626
rect 8430 54462 8482 54514
rect 9102 54462 9154 54514
rect 10222 54462 10274 54514
rect 11006 54462 11058 54514
rect 12238 54462 12290 54514
rect 13134 54462 13186 54514
rect 14926 54462 14978 54514
rect 15598 54462 15650 54514
rect 15934 54462 15986 54514
rect 16158 54462 16210 54514
rect 16494 54462 16546 54514
rect 16606 54462 16658 54514
rect 17726 54462 17778 54514
rect 18174 54462 18226 54514
rect 20638 54462 20690 54514
rect 20750 54462 20802 54514
rect 21086 54462 21138 54514
rect 21646 54462 21698 54514
rect 21870 54462 21922 54514
rect 24782 54462 24834 54514
rect 26798 54462 26850 54514
rect 28030 54462 28082 54514
rect 28702 54462 28754 54514
rect 29150 54462 29202 54514
rect 30606 54462 30658 54514
rect 31166 54462 31218 54514
rect 32622 54462 32674 54514
rect 35646 54462 35698 54514
rect 36878 54462 36930 54514
rect 38446 54462 38498 54514
rect 38782 54462 38834 54514
rect 39342 54462 39394 54514
rect 40126 54462 40178 54514
rect 40350 54462 40402 54514
rect 42030 54462 42082 54514
rect 46174 54462 46226 54514
rect 2046 54350 2098 54402
rect 2494 54350 2546 54402
rect 2942 54350 2994 54402
rect 3390 54350 3442 54402
rect 3838 54350 3890 54402
rect 4174 54350 4226 54402
rect 4734 54350 4786 54402
rect 5630 54350 5682 54402
rect 6078 54350 6130 54402
rect 6526 54350 6578 54402
rect 6974 54350 7026 54402
rect 7982 54350 8034 54402
rect 8542 54350 8594 54402
rect 12686 54350 12738 54402
rect 16382 54350 16434 54402
rect 19742 54350 19794 54402
rect 21758 54350 21810 54402
rect 22766 54350 22818 54402
rect 26686 54350 26738 54402
rect 29934 54350 29986 54402
rect 31278 54350 31330 54402
rect 31838 54350 31890 54402
rect 31950 54350 32002 54402
rect 33518 54350 33570 54402
rect 34190 54350 34242 54402
rect 37662 54350 37714 54402
rect 39902 54350 39954 54402
rect 42142 54350 42194 54402
rect 4062 54238 4114 54290
rect 4622 54238 4674 54290
rect 14254 54238 14306 54290
rect 17950 54238 18002 54290
rect 18398 54238 18450 54290
rect 18622 54238 18674 54290
rect 18846 54238 18898 54290
rect 23438 54238 23490 54290
rect 36990 54238 37042 54290
rect 43598 54238 43650 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 9438 53902 9490 53954
rect 20526 53902 20578 53954
rect 22206 53902 22258 53954
rect 28254 53902 28306 53954
rect 28478 53902 28530 53954
rect 28926 53902 28978 53954
rect 30494 53902 30546 53954
rect 34190 53902 34242 53954
rect 39454 53902 39506 53954
rect 39566 53902 39618 53954
rect 42702 53902 42754 53954
rect 42926 53902 42978 53954
rect 5070 53790 5122 53842
rect 9102 53790 9154 53842
rect 25454 53790 25506 53842
rect 28030 53790 28082 53842
rect 30830 53790 30882 53842
rect 32062 53790 32114 53842
rect 33406 53790 33458 53842
rect 33966 53790 34018 53842
rect 37550 53790 37602 53842
rect 39790 53790 39842 53842
rect 5742 53678 5794 53730
rect 6974 53678 7026 53730
rect 9886 53678 9938 53730
rect 10670 53678 10722 53730
rect 14702 53678 14754 53730
rect 15038 53678 15090 53730
rect 15598 53678 15650 53730
rect 16046 53678 16098 53730
rect 16942 53678 16994 53730
rect 17614 53678 17666 53730
rect 17838 53678 17890 53730
rect 18062 53678 18114 53730
rect 18174 53678 18226 53730
rect 19966 53678 20018 53730
rect 20190 53678 20242 53730
rect 21646 53678 21698 53730
rect 22654 53678 22706 53730
rect 24110 53678 24162 53730
rect 29822 53678 29874 53730
rect 30158 53678 30210 53730
rect 31838 53678 31890 53730
rect 33630 53678 33682 53730
rect 34638 53678 34690 53730
rect 35870 53678 35922 53730
rect 37662 53678 37714 53730
rect 37998 53678 38050 53730
rect 41134 53678 41186 53730
rect 43150 53678 43202 53730
rect 43598 53678 43650 53730
rect 1822 53566 1874 53618
rect 6750 53566 6802 53618
rect 7646 53566 7698 53618
rect 7758 53566 7810 53618
rect 9326 53566 9378 53618
rect 10110 53566 10162 53618
rect 10222 53566 10274 53618
rect 13806 53566 13858 53618
rect 16606 53566 16658 53618
rect 18846 53566 18898 53618
rect 23998 53566 24050 53618
rect 25006 53566 25058 53618
rect 26574 53566 26626 53618
rect 27022 53566 27074 53618
rect 27358 53566 27410 53618
rect 30382 53566 30434 53618
rect 32734 53566 32786 53618
rect 33966 53566 34018 53618
rect 39902 53566 39954 53618
rect 40910 53566 40962 53618
rect 41358 53566 41410 53618
rect 42590 53566 42642 53618
rect 45838 53566 45890 53618
rect 2270 53454 2322 53506
rect 2718 53454 2770 53506
rect 3166 53454 3218 53506
rect 3614 53454 3666 53506
rect 4062 53454 4114 53506
rect 4510 53454 4562 53506
rect 6302 53454 6354 53506
rect 7982 53454 8034 53506
rect 8654 53454 8706 53506
rect 11118 53454 11170 53506
rect 11230 53454 11282 53506
rect 11342 53454 11394 53506
rect 11902 53454 11954 53506
rect 12574 53454 12626 53506
rect 13022 53454 13074 53506
rect 14142 53454 14194 53506
rect 14814 53454 14866 53506
rect 16718 53454 16770 53506
rect 18958 53454 19010 53506
rect 19182 53454 19234 53506
rect 21870 53454 21922 53506
rect 22094 53454 22146 53506
rect 22766 53454 22818 53506
rect 22990 53454 23042 53506
rect 24558 53454 24610 53506
rect 26126 53454 26178 53506
rect 35086 53454 35138 53506
rect 35646 53454 35698 53506
rect 35758 53454 35810 53506
rect 36094 53454 36146 53506
rect 36766 53454 36818 53506
rect 40350 53454 40402 53506
rect 41022 53454 41074 53506
rect 41918 53454 41970 53506
rect 44046 53454 44098 53506
rect 45950 53454 46002 53506
rect 46062 53454 46114 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 3502 53118 3554 53170
rect 4286 53118 4338 53170
rect 5630 53118 5682 53170
rect 6190 53118 6242 53170
rect 6526 53118 6578 53170
rect 9774 53118 9826 53170
rect 10670 53118 10722 53170
rect 10894 53118 10946 53170
rect 17614 53118 17666 53170
rect 18398 53118 18450 53170
rect 20526 53118 20578 53170
rect 22542 53118 22594 53170
rect 23550 53118 23602 53170
rect 26798 53118 26850 53170
rect 31166 53118 31218 53170
rect 33742 53118 33794 53170
rect 36766 53118 36818 53170
rect 37550 53118 37602 53170
rect 39118 53118 39170 53170
rect 39566 53118 39618 53170
rect 40014 53118 40066 53170
rect 43038 53118 43090 53170
rect 7310 53006 7362 53058
rect 12686 53006 12738 53058
rect 13694 53006 13746 53058
rect 21422 53006 21474 53058
rect 26014 53006 26066 53058
rect 26126 53006 26178 53058
rect 27918 53006 27970 53058
rect 35646 53006 35698 53058
rect 35758 53006 35810 53058
rect 36542 53006 36594 53058
rect 38222 53006 38274 53058
rect 40798 53006 40850 53058
rect 42478 53006 42530 53058
rect 43598 53006 43650 53058
rect 43710 53006 43762 53058
rect 7198 52894 7250 52946
rect 8094 52894 8146 52946
rect 11006 52894 11058 52946
rect 11902 52894 11954 52946
rect 12574 52894 12626 52946
rect 13134 52894 13186 52946
rect 13358 52894 13410 52946
rect 14702 52894 14754 52946
rect 21198 52894 21250 52946
rect 21982 52894 22034 52946
rect 22206 52894 22258 52946
rect 26686 52894 26738 52946
rect 26910 52894 26962 52946
rect 27358 52894 27410 52946
rect 27806 52894 27858 52946
rect 30942 52894 30994 52946
rect 33966 52894 34018 52946
rect 35982 52894 36034 52946
rect 36430 52894 36482 52946
rect 37438 52894 37490 52946
rect 37774 52894 37826 52946
rect 41582 52894 41634 52946
rect 41806 52894 41858 52946
rect 42142 52894 42194 52946
rect 42254 52894 42306 52946
rect 43934 52894 43986 52946
rect 44830 52894 44882 52946
rect 45950 52894 46002 52946
rect 2158 52782 2210 52834
rect 2606 52782 2658 52834
rect 2942 52782 2994 52834
rect 3950 52782 4002 52834
rect 4846 52782 4898 52834
rect 5294 52782 5346 52834
rect 8654 52782 8706 52834
rect 9102 52782 9154 52834
rect 10334 52782 10386 52834
rect 14366 52782 14418 52834
rect 15262 52782 15314 52834
rect 15598 52782 15650 52834
rect 16158 52782 16210 52834
rect 16494 52782 16546 52834
rect 16942 52782 16994 52834
rect 18958 52782 19010 52834
rect 19406 52782 19458 52834
rect 20190 52782 20242 52834
rect 23102 52782 23154 52834
rect 24446 52782 24498 52834
rect 24782 52782 24834 52834
rect 28478 52782 28530 52834
rect 28926 52782 28978 52834
rect 29374 52782 29426 52834
rect 29822 52782 29874 52834
rect 30270 52782 30322 52834
rect 31614 52782 31666 52834
rect 32062 52782 32114 52834
rect 32622 52782 32674 52834
rect 34526 52782 34578 52834
rect 35198 52782 35250 52834
rect 38670 52782 38722 52834
rect 42366 52782 42418 52834
rect 44494 52782 44546 52834
rect 2046 52670 2098 52722
rect 3726 52670 3778 52722
rect 4174 52670 4226 52722
rect 7310 52670 7362 52722
rect 18286 52670 18338 52722
rect 19182 52670 19234 52722
rect 26014 52670 26066 52722
rect 27918 52670 27970 52722
rect 28702 52670 28754 52722
rect 29150 52670 29202 52722
rect 29822 52670 29874 52722
rect 33630 52670 33682 52722
rect 46174 52670 46226 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 12014 52334 12066 52386
rect 18286 52334 18338 52386
rect 18510 52334 18562 52386
rect 19406 52334 19458 52386
rect 20078 52334 20130 52386
rect 25230 52334 25282 52386
rect 27470 52334 27522 52386
rect 33070 52334 33122 52386
rect 44718 52334 44770 52386
rect 4510 52222 4562 52274
rect 5854 52222 5906 52274
rect 12910 52222 12962 52274
rect 17502 52222 17554 52274
rect 19182 52222 19234 52274
rect 23550 52222 23602 52274
rect 27134 52222 27186 52274
rect 29822 52222 29874 52274
rect 34414 52222 34466 52274
rect 35534 52222 35586 52274
rect 37550 52222 37602 52274
rect 40014 52222 40066 52274
rect 40910 52222 40962 52274
rect 41582 52222 41634 52274
rect 42478 52222 42530 52274
rect 3278 52110 3330 52162
rect 5070 52110 5122 52162
rect 6974 52110 7026 52162
rect 7198 52110 7250 52162
rect 8206 52110 8258 52162
rect 8878 52110 8930 52162
rect 9998 52110 10050 52162
rect 11454 52110 11506 52162
rect 11902 52110 11954 52162
rect 12798 52110 12850 52162
rect 14478 52110 14530 52162
rect 18174 52110 18226 52162
rect 19630 52110 19682 52162
rect 20526 52110 20578 52162
rect 20862 52110 20914 52162
rect 22542 52110 22594 52162
rect 24110 52110 24162 52162
rect 26350 52110 26402 52162
rect 27246 52110 27298 52162
rect 30046 52110 30098 52162
rect 32510 52110 32562 52162
rect 35870 52110 35922 52162
rect 36318 52110 36370 52162
rect 36766 52110 36818 52162
rect 40462 52110 40514 52162
rect 42814 52110 42866 52162
rect 44382 52110 44434 52162
rect 45390 52110 45442 52162
rect 54910 52110 54962 52162
rect 56030 52110 56082 52162
rect 7422 51998 7474 52050
rect 8318 51998 8370 52050
rect 8766 51998 8818 52050
rect 11118 51998 11170 52050
rect 12574 51998 12626 52050
rect 14030 51998 14082 52050
rect 15038 51998 15090 52050
rect 15374 51998 15426 52050
rect 16270 51998 16322 52050
rect 16494 51998 16546 52050
rect 20638 51998 20690 52050
rect 22318 51998 22370 52050
rect 22878 51998 22930 52050
rect 23662 51998 23714 52050
rect 24670 51998 24722 52050
rect 24894 51998 24946 52050
rect 25566 51998 25618 52050
rect 26126 51998 26178 52050
rect 28478 51998 28530 52050
rect 30718 51998 30770 52050
rect 31838 51998 31890 52050
rect 32062 51998 32114 52050
rect 32958 51998 33010 52050
rect 33742 51998 33794 52050
rect 38446 51998 38498 52050
rect 43262 51998 43314 52050
rect 1934 51886 1986 51938
rect 2382 51886 2434 51938
rect 2830 51886 2882 51938
rect 3726 51886 3778 51938
rect 4174 51886 4226 51938
rect 9102 51886 9154 51938
rect 11230 51886 11282 51938
rect 12350 51886 12402 51938
rect 13694 51886 13746 51938
rect 13806 51886 13858 51938
rect 13918 51886 13970 51938
rect 16382 51886 16434 51938
rect 16718 51886 16770 51938
rect 18174 51886 18226 51938
rect 21758 51886 21810 51938
rect 22766 51886 22818 51938
rect 23326 51886 23378 51938
rect 23550 51886 23602 51938
rect 25118 51886 25170 51938
rect 28814 51886 28866 51938
rect 31278 51886 31330 51938
rect 31950 51886 32002 51938
rect 33070 51886 33122 51938
rect 33854 51886 33906 51938
rect 34078 51886 34130 51938
rect 37662 51886 37714 51938
rect 38558 51886 38610 51938
rect 38782 51886 38834 51938
rect 39230 51886 39282 51938
rect 39566 51886 39618 51938
rect 44606 51886 44658 51938
rect 45838 51886 45890 51938
rect 45950 51886 46002 51938
rect 46062 51886 46114 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 1822 51550 1874 51602
rect 2718 51550 2770 51602
rect 5742 51550 5794 51602
rect 6526 51550 6578 51602
rect 6862 51550 6914 51602
rect 8542 51550 8594 51602
rect 8990 51550 9042 51602
rect 9886 51550 9938 51602
rect 14926 51550 14978 51602
rect 17726 51550 17778 51602
rect 17950 51550 18002 51602
rect 19294 51550 19346 51602
rect 20190 51550 20242 51602
rect 20526 51550 20578 51602
rect 21310 51550 21362 51602
rect 22542 51550 22594 51602
rect 23774 51550 23826 51602
rect 24558 51550 24610 51602
rect 31054 51550 31106 51602
rect 34750 51550 34802 51602
rect 35982 51550 36034 51602
rect 39790 51550 39842 51602
rect 40350 51550 40402 51602
rect 41694 51550 41746 51602
rect 48750 51550 48802 51602
rect 4846 51438 4898 51490
rect 5406 51438 5458 51490
rect 7870 51438 7922 51490
rect 7982 51438 8034 51490
rect 8094 51438 8146 51490
rect 12238 51438 12290 51490
rect 16382 51438 16434 51490
rect 16494 51438 16546 51490
rect 23438 51438 23490 51490
rect 23662 51438 23714 51490
rect 24782 51438 24834 51490
rect 25566 51438 25618 51490
rect 26238 51438 26290 51490
rect 28478 51438 28530 51490
rect 30382 51438 30434 51490
rect 31726 51438 31778 51490
rect 33854 51438 33906 51490
rect 36766 51438 36818 51490
rect 38110 51438 38162 51490
rect 38894 51438 38946 51490
rect 43598 51438 43650 51490
rect 44942 51438 44994 51490
rect 4622 51326 4674 51378
rect 9998 51326 10050 51378
rect 10222 51326 10274 51378
rect 10446 51326 10498 51378
rect 11006 51326 11058 51378
rect 11342 51326 11394 51378
rect 11678 51326 11730 51378
rect 12126 51326 12178 51378
rect 12462 51326 12514 51378
rect 12798 51326 12850 51378
rect 13694 51326 13746 51378
rect 15150 51326 15202 51378
rect 16158 51326 16210 51378
rect 16942 51326 16994 51378
rect 17614 51326 17666 51378
rect 18174 51326 18226 51378
rect 18958 51326 19010 51378
rect 19406 51326 19458 51378
rect 19518 51326 19570 51378
rect 22094 51326 22146 51378
rect 22430 51326 22482 51378
rect 22766 51326 22818 51378
rect 23886 51326 23938 51378
rect 23998 51326 24050 51378
rect 24894 51326 24946 51378
rect 26574 51326 26626 51378
rect 27918 51326 27970 51378
rect 28366 51326 28418 51378
rect 30046 51326 30098 51378
rect 31614 51326 31666 51378
rect 33742 51326 33794 51378
rect 34862 51326 34914 51378
rect 35646 51326 35698 51378
rect 38782 51326 38834 51378
rect 39678 51326 39730 51378
rect 42142 51326 42194 51378
rect 42926 51326 42978 51378
rect 44494 51326 44546 51378
rect 44830 51326 44882 51378
rect 45950 51326 46002 51378
rect 48414 51326 48466 51378
rect 2270 51214 2322 51266
rect 3166 51214 3218 51266
rect 3614 51214 3666 51266
rect 4062 51214 4114 51266
rect 10110 51214 10162 51266
rect 10670 51214 10722 51266
rect 10894 51214 10946 51266
rect 11454 51214 11506 51266
rect 13918 51214 13970 51266
rect 14366 51214 14418 51266
rect 16494 51214 16546 51266
rect 21870 51214 21922 51266
rect 22654 51214 22706 51266
rect 27022 51214 27074 51266
rect 28254 51214 28306 51266
rect 29374 51214 29426 51266
rect 35422 51214 35474 51266
rect 37326 51214 37378 51266
rect 38222 51214 38274 51266
rect 40798 51214 40850 51266
rect 42814 51214 42866 51266
rect 45726 51214 45778 51266
rect 47854 51214 47906 51266
rect 3502 51102 3554 51154
rect 4062 51102 4114 51154
rect 26574 51102 26626 51154
rect 32398 51102 32450 51154
rect 32734 51102 32786 51154
rect 36542 51102 36594 51154
rect 36878 51102 36930 51154
rect 37886 51102 37938 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 5854 50766 5906 50818
rect 9662 50766 9714 50818
rect 9998 50766 10050 50818
rect 12462 50766 12514 50818
rect 26574 50766 26626 50818
rect 27246 50766 27298 50818
rect 27918 50766 27970 50818
rect 34190 50766 34242 50818
rect 34526 50766 34578 50818
rect 6638 50654 6690 50706
rect 8206 50654 8258 50706
rect 11006 50654 11058 50706
rect 14254 50654 14306 50706
rect 15710 50654 15762 50706
rect 16046 50654 16098 50706
rect 24446 50654 24498 50706
rect 29934 50654 29986 50706
rect 36094 50654 36146 50706
rect 37438 50654 37490 50706
rect 38110 50654 38162 50706
rect 44158 50654 44210 50706
rect 46062 50654 46114 50706
rect 46510 50654 46562 50706
rect 3054 50542 3106 50594
rect 4398 50542 4450 50594
rect 4622 50542 4674 50594
rect 4846 50542 4898 50594
rect 9998 50542 10050 50594
rect 11342 50542 11394 50594
rect 11566 50542 11618 50594
rect 12014 50542 12066 50594
rect 12238 50542 12290 50594
rect 13694 50542 13746 50594
rect 13918 50542 13970 50594
rect 16158 50542 16210 50594
rect 17726 50542 17778 50594
rect 19182 50542 19234 50594
rect 20078 50542 20130 50594
rect 22318 50542 22370 50594
rect 25790 50542 25842 50594
rect 26238 50542 26290 50594
rect 27470 50542 27522 50594
rect 29822 50542 29874 50594
rect 32398 50542 32450 50594
rect 32734 50542 32786 50594
rect 34526 50542 34578 50594
rect 35534 50542 35586 50594
rect 36206 50542 36258 50594
rect 39566 50542 39618 50594
rect 41582 50542 41634 50594
rect 42254 50542 42306 50594
rect 42478 50542 42530 50594
rect 45838 50542 45890 50594
rect 1934 50430 1986 50482
rect 5966 50430 6018 50482
rect 9102 50430 9154 50482
rect 14142 50430 14194 50482
rect 14254 50430 14306 50482
rect 15262 50430 15314 50482
rect 17390 50430 17442 50482
rect 18286 50430 18338 50482
rect 22878 50430 22930 50482
rect 23774 50430 23826 50482
rect 23886 50430 23938 50482
rect 24894 50430 24946 50482
rect 27806 50430 27858 50482
rect 28030 50430 28082 50482
rect 28478 50430 28530 50482
rect 30718 50430 30770 50482
rect 31166 50430 31218 50482
rect 32062 50430 32114 50482
rect 33406 50430 33458 50482
rect 35086 50430 35138 50482
rect 36542 50430 36594 50482
rect 38334 50430 38386 50482
rect 40238 50430 40290 50482
rect 3950 50318 4002 50370
rect 4510 50318 4562 50370
rect 5854 50318 5906 50370
rect 7086 50318 7138 50370
rect 7870 50318 7922 50370
rect 8654 50318 8706 50370
rect 18622 50318 18674 50370
rect 19518 50318 19570 50370
rect 20190 50318 20242 50370
rect 20414 50318 20466 50370
rect 20862 50318 20914 50370
rect 21982 50318 22034 50370
rect 23214 50318 23266 50370
rect 24110 50318 24162 50370
rect 26462 50318 26514 50370
rect 32510 50318 32562 50370
rect 40798 50318 40850 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 1934 49982 1986 50034
rect 2382 49982 2434 50034
rect 4062 49982 4114 50034
rect 5854 49982 5906 50034
rect 11006 49982 11058 50034
rect 12350 49982 12402 50034
rect 13246 49982 13298 50034
rect 16046 49982 16098 50034
rect 16718 49982 16770 50034
rect 19854 49982 19906 50034
rect 19966 49982 20018 50034
rect 21758 49982 21810 50034
rect 22318 49982 22370 50034
rect 23326 49982 23378 50034
rect 26014 49982 26066 50034
rect 27246 49982 27298 50034
rect 28030 49982 28082 50034
rect 28366 49982 28418 50034
rect 29374 49982 29426 50034
rect 31278 49982 31330 50034
rect 31950 49982 32002 50034
rect 32622 49982 32674 50034
rect 36542 49982 36594 50034
rect 37886 49982 37938 50034
rect 39118 49982 39170 50034
rect 39566 49982 39618 50034
rect 40574 49982 40626 50034
rect 41918 49982 41970 50034
rect 42142 49982 42194 50034
rect 45054 49982 45106 50034
rect 3166 49870 3218 49922
rect 11902 49870 11954 49922
rect 15934 49870 15986 49922
rect 16942 49870 16994 49922
rect 23214 49870 23266 49922
rect 24222 49870 24274 49922
rect 24334 49870 24386 49922
rect 24894 49870 24946 49922
rect 27806 49870 27858 49922
rect 32062 49870 32114 49922
rect 41806 49870 41858 49922
rect 42478 49870 42530 49922
rect 2830 49758 2882 49810
rect 3726 49758 3778 49810
rect 4062 49758 4114 49810
rect 4286 49758 4338 49810
rect 6862 49758 6914 49810
rect 7086 49758 7138 49810
rect 7534 49758 7586 49810
rect 8094 49758 8146 49810
rect 8654 49758 8706 49810
rect 11566 49758 11618 49810
rect 12910 49758 12962 49810
rect 15486 49758 15538 49810
rect 15710 49758 15762 49810
rect 16382 49758 16434 49810
rect 20078 49758 20130 49810
rect 21534 49758 21586 49810
rect 22654 49758 22706 49810
rect 24558 49758 24610 49810
rect 28254 49758 28306 49810
rect 36766 49758 36818 49810
rect 40126 49758 40178 49810
rect 40350 49758 40402 49810
rect 44718 49758 44770 49810
rect 45166 49758 45218 49810
rect 45390 49758 45442 49810
rect 5070 49646 5122 49698
rect 5406 49646 5458 49698
rect 9998 49646 10050 49698
rect 10446 49646 10498 49698
rect 10670 49646 10722 49698
rect 14030 49646 14082 49698
rect 14478 49646 14530 49698
rect 14926 49646 14978 49698
rect 17614 49646 17666 49698
rect 18398 49646 18450 49698
rect 18846 49646 18898 49698
rect 19630 49646 19682 49698
rect 20862 49646 20914 49698
rect 25566 49646 25618 49698
rect 26686 49646 26738 49698
rect 28366 49646 28418 49698
rect 28926 49646 28978 49698
rect 29822 49646 29874 49698
rect 30270 49646 30322 49698
rect 30718 49646 30770 49698
rect 31838 49646 31890 49698
rect 33518 49646 33570 49698
rect 33966 49646 34018 49698
rect 34750 49646 34802 49698
rect 35198 49646 35250 49698
rect 35646 49646 35698 49698
rect 37326 49646 37378 49698
rect 38222 49646 38274 49698
rect 38670 49646 38722 49698
rect 40238 49646 40290 49698
rect 43486 49646 43538 49698
rect 6974 49534 7026 49586
rect 14590 49534 14642 49586
rect 14926 49534 14978 49586
rect 17054 49534 17106 49586
rect 19406 49534 19458 49586
rect 23326 49534 23378 49586
rect 26910 49534 26962 49586
rect 30270 49534 30322 49586
rect 31054 49534 31106 49586
rect 43598 49534 43650 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 4846 49198 4898 49250
rect 11566 49198 11618 49250
rect 13918 49198 13970 49250
rect 14254 49198 14306 49250
rect 21422 49198 21474 49250
rect 22206 49198 22258 49250
rect 23214 49198 23266 49250
rect 25342 49198 25394 49250
rect 25902 49198 25954 49250
rect 32398 49198 32450 49250
rect 40686 49198 40738 49250
rect 3726 49086 3778 49138
rect 5966 49086 6018 49138
rect 7982 49086 8034 49138
rect 8990 49086 9042 49138
rect 12910 49086 12962 49138
rect 16942 49086 16994 49138
rect 18622 49086 18674 49138
rect 19854 49086 19906 49138
rect 24110 49086 24162 49138
rect 24558 49086 24610 49138
rect 25118 49086 25170 49138
rect 25902 49086 25954 49138
rect 27694 49086 27746 49138
rect 28254 49086 28306 49138
rect 33630 49086 33682 49138
rect 33854 49086 33906 49138
rect 36318 49086 36370 49138
rect 46622 49086 46674 49138
rect 2718 48974 2770 49026
rect 6526 48974 6578 49026
rect 6974 48974 7026 49026
rect 7646 48974 7698 49026
rect 9438 48974 9490 49026
rect 13806 48974 13858 49026
rect 14142 48974 14194 49026
rect 16158 48974 16210 49026
rect 17390 48974 17442 49026
rect 18286 48974 18338 49026
rect 18846 48974 18898 49026
rect 19070 48974 19122 49026
rect 19742 48974 19794 49026
rect 23326 48974 23378 49026
rect 23550 48974 23602 49026
rect 30158 48974 30210 49026
rect 30606 48974 30658 49026
rect 33070 48974 33122 49026
rect 34190 48974 34242 49026
rect 37774 48974 37826 49026
rect 38222 48974 38274 49026
rect 40238 48974 40290 49026
rect 40462 48974 40514 49026
rect 43710 48974 43762 49026
rect 43934 48974 43986 49026
rect 46510 48974 46562 49026
rect 1822 48862 1874 48914
rect 4062 48862 4114 48914
rect 4734 48862 4786 48914
rect 4846 48862 4898 48914
rect 7982 48862 8034 48914
rect 9774 48862 9826 48914
rect 10558 48862 10610 48914
rect 10894 48862 10946 48914
rect 11566 48862 11618 48914
rect 11678 48862 11730 48914
rect 16270 48862 16322 48914
rect 16942 48862 16994 48914
rect 19966 48862 20018 48914
rect 26910 48862 26962 48914
rect 27246 48862 27298 48914
rect 29822 48862 29874 48914
rect 31502 48862 31554 48914
rect 32286 48862 32338 48914
rect 33182 48862 33234 48914
rect 37550 48862 37602 48914
rect 41134 48862 41186 48914
rect 41694 48862 41746 48914
rect 42702 48862 42754 48914
rect 42814 48862 42866 48914
rect 43486 48862 43538 48914
rect 45502 48862 45554 48914
rect 45614 48862 45666 48914
rect 47406 48862 47458 48914
rect 2158 48750 2210 48802
rect 3054 48750 3106 48802
rect 3614 48750 3666 48802
rect 3838 48750 3890 48802
rect 12238 48750 12290 48802
rect 15150 48750 15202 48802
rect 15486 48750 15538 48802
rect 18622 48750 18674 48802
rect 20190 48750 20242 48802
rect 20750 48750 20802 48802
rect 21646 48750 21698 48802
rect 22094 48750 22146 48802
rect 22542 48750 22594 48802
rect 23214 48750 23266 48802
rect 25454 48750 25506 48802
rect 26350 48750 26402 48802
rect 28814 48750 28866 48802
rect 30942 48750 30994 48802
rect 32398 48750 32450 48802
rect 35086 48750 35138 48802
rect 35534 48750 35586 48802
rect 36878 48750 36930 48802
rect 37886 48750 37938 48802
rect 37998 48750 38050 48802
rect 38670 48750 38722 48802
rect 41582 48750 41634 48802
rect 43038 48750 43090 48802
rect 43710 48750 43762 48802
rect 45838 48750 45890 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 4846 48414 4898 48466
rect 7758 48414 7810 48466
rect 11678 48414 11730 48466
rect 15262 48414 15314 48466
rect 25566 48414 25618 48466
rect 27134 48414 27186 48466
rect 29038 48414 29090 48466
rect 31838 48414 31890 48466
rect 32734 48414 32786 48466
rect 34862 48414 34914 48466
rect 35870 48414 35922 48466
rect 38894 48414 38946 48466
rect 42142 48414 42194 48466
rect 3166 48302 3218 48354
rect 4174 48302 4226 48354
rect 6414 48302 6466 48354
rect 6862 48302 6914 48354
rect 7422 48302 7474 48354
rect 8654 48302 8706 48354
rect 9998 48302 10050 48354
rect 10334 48302 10386 48354
rect 12910 48302 12962 48354
rect 13246 48302 13298 48354
rect 14926 48302 14978 48354
rect 15934 48302 15986 48354
rect 16606 48302 16658 48354
rect 16830 48302 16882 48354
rect 18174 48302 18226 48354
rect 19854 48302 19906 48354
rect 20078 48302 20130 48354
rect 23662 48302 23714 48354
rect 24782 48302 24834 48354
rect 32286 48302 32338 48354
rect 32846 48302 32898 48354
rect 33854 48302 33906 48354
rect 33966 48302 34018 48354
rect 36990 48302 37042 48354
rect 37774 48302 37826 48354
rect 38558 48302 38610 48354
rect 39790 48302 39842 48354
rect 44270 48302 44322 48354
rect 44494 48302 44546 48354
rect 45390 48302 45442 48354
rect 2830 48190 2882 48242
rect 5070 48190 5122 48242
rect 5406 48190 5458 48242
rect 6302 48190 6354 48242
rect 6638 48190 6690 48242
rect 8990 48190 9042 48242
rect 10894 48190 10946 48242
rect 11118 48190 11170 48242
rect 11678 48190 11730 48242
rect 12686 48190 12738 48242
rect 13806 48190 13858 48242
rect 14814 48190 14866 48242
rect 15822 48190 15874 48242
rect 17726 48190 17778 48242
rect 18398 48190 18450 48242
rect 18846 48190 18898 48242
rect 19294 48190 19346 48242
rect 22990 48190 23042 48242
rect 23214 48190 23266 48242
rect 23550 48190 23602 48242
rect 23886 48190 23938 48242
rect 26686 48190 26738 48242
rect 27358 48190 27410 48242
rect 29710 48190 29762 48242
rect 29934 48190 29986 48242
rect 30382 48190 30434 48242
rect 32622 48190 32674 48242
rect 33630 48190 33682 48242
rect 36430 48190 36482 48242
rect 36878 48190 36930 48242
rect 37886 48190 37938 48242
rect 38110 48190 38162 48242
rect 40014 48190 40066 48242
rect 41582 48190 41634 48242
rect 43374 48190 43426 48242
rect 1934 48078 1986 48130
rect 2382 48078 2434 48130
rect 4286 48078 4338 48130
rect 4958 48078 5010 48130
rect 12126 48078 12178 48130
rect 13134 48078 13186 48130
rect 16942 48078 16994 48130
rect 20190 48078 20242 48130
rect 20638 48078 20690 48130
rect 21310 48078 21362 48130
rect 21870 48078 21922 48130
rect 22318 48078 22370 48130
rect 23774 48078 23826 48130
rect 24558 48078 24610 48130
rect 24894 48078 24946 48130
rect 26014 48078 26066 48130
rect 27246 48078 27298 48130
rect 27918 48078 27970 48130
rect 28590 48078 28642 48130
rect 29822 48078 29874 48130
rect 30718 48078 30770 48130
rect 31166 48078 31218 48130
rect 35310 48078 35362 48130
rect 37550 48078 37602 48130
rect 40350 48078 40402 48130
rect 43486 48078 43538 48130
rect 43710 48078 43762 48130
rect 45278 48078 45330 48130
rect 3950 47966 4002 48018
rect 11342 47966 11394 48018
rect 28702 47966 28754 48018
rect 29486 47966 29538 48018
rect 34414 47966 34466 48018
rect 35422 47966 35474 48018
rect 36206 47966 36258 48018
rect 36654 47966 36706 48018
rect 41806 47966 41858 48018
rect 44606 47966 44658 48018
rect 45166 47966 45218 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 5742 47630 5794 47682
rect 6302 47630 6354 47682
rect 14030 47630 14082 47682
rect 14142 47630 14194 47682
rect 14366 47630 14418 47682
rect 17614 47630 17666 47682
rect 20302 47630 20354 47682
rect 20526 47630 20578 47682
rect 22542 47630 22594 47682
rect 24446 47630 24498 47682
rect 30942 47630 30994 47682
rect 37438 47630 37490 47682
rect 3054 47518 3106 47570
rect 4510 47518 4562 47570
rect 5630 47518 5682 47570
rect 6190 47518 6242 47570
rect 8318 47518 8370 47570
rect 9214 47518 9266 47570
rect 9998 47518 10050 47570
rect 12014 47518 12066 47570
rect 12798 47518 12850 47570
rect 16270 47518 16322 47570
rect 18958 47518 19010 47570
rect 23326 47518 23378 47570
rect 25454 47518 25506 47570
rect 27134 47518 27186 47570
rect 28478 47518 28530 47570
rect 30270 47518 30322 47570
rect 31950 47518 32002 47570
rect 37886 47518 37938 47570
rect 39006 47518 39058 47570
rect 45614 47518 45666 47570
rect 2046 47406 2098 47458
rect 3166 47406 3218 47458
rect 8766 47406 8818 47458
rect 9438 47406 9490 47458
rect 11118 47406 11170 47458
rect 14478 47406 14530 47458
rect 15262 47406 15314 47458
rect 16494 47406 16546 47458
rect 17054 47406 17106 47458
rect 17166 47406 17218 47458
rect 17502 47406 17554 47458
rect 19630 47406 19682 47458
rect 19854 47406 19906 47458
rect 19966 47406 20018 47458
rect 21982 47406 22034 47458
rect 22766 47406 22818 47458
rect 23102 47406 23154 47458
rect 23438 47406 23490 47458
rect 24110 47406 24162 47458
rect 24446 47406 24498 47458
rect 26574 47406 26626 47458
rect 27022 47406 27074 47458
rect 28142 47406 28194 47458
rect 30158 47406 30210 47458
rect 32846 47406 32898 47458
rect 33742 47406 33794 47458
rect 33854 47406 33906 47458
rect 34302 47406 34354 47458
rect 34974 47406 35026 47458
rect 35198 47406 35250 47458
rect 35422 47406 35474 47458
rect 35534 47406 35586 47458
rect 38110 47406 38162 47458
rect 38334 47406 38386 47458
rect 41022 47406 41074 47458
rect 41470 47406 41522 47458
rect 43486 47406 43538 47458
rect 43934 47406 43986 47458
rect 46062 47406 46114 47458
rect 6974 47294 7026 47346
rect 8990 47294 9042 47346
rect 10334 47294 10386 47346
rect 10894 47294 10946 47346
rect 12574 47294 12626 47346
rect 21646 47294 21698 47346
rect 26014 47294 26066 47346
rect 27582 47294 27634 47346
rect 28702 47294 28754 47346
rect 33182 47294 33234 47346
rect 34078 47294 34130 47346
rect 38558 47294 38610 47346
rect 39678 47294 39730 47346
rect 41918 47294 41970 47346
rect 43374 47294 43426 47346
rect 2382 47182 2434 47234
rect 3054 47182 3106 47234
rect 5070 47182 5122 47234
rect 6638 47182 6690 47234
rect 7870 47182 7922 47234
rect 12798 47182 12850 47234
rect 14926 47182 14978 47234
rect 15150 47182 15202 47234
rect 19742 47182 19794 47234
rect 23214 47182 23266 47234
rect 25118 47182 25170 47234
rect 28478 47182 28530 47234
rect 31502 47182 31554 47234
rect 36094 47182 36146 47234
rect 36430 47182 36482 47234
rect 45502 47182 45554 47234
rect 45726 47182 45778 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 1934 46846 1986 46898
rect 2830 46846 2882 46898
rect 3166 46846 3218 46898
rect 5406 46846 5458 46898
rect 8094 46846 8146 46898
rect 8878 46846 8930 46898
rect 9662 46846 9714 46898
rect 9774 46846 9826 46898
rect 10670 46846 10722 46898
rect 13918 46846 13970 46898
rect 16382 46846 16434 46898
rect 16494 46846 16546 46898
rect 18510 46846 18562 46898
rect 19070 46846 19122 46898
rect 19854 46846 19906 46898
rect 21086 46846 21138 46898
rect 22542 46846 22594 46898
rect 23102 46846 23154 46898
rect 26126 46846 26178 46898
rect 27582 46846 27634 46898
rect 30718 46846 30770 46898
rect 32510 46846 32562 46898
rect 33630 46846 33682 46898
rect 34414 46846 34466 46898
rect 36542 46846 36594 46898
rect 39230 46846 39282 46898
rect 40462 46846 40514 46898
rect 4286 46734 4338 46786
rect 6526 46734 6578 46786
rect 7982 46734 8034 46786
rect 8766 46734 8818 46786
rect 10222 46734 10274 46786
rect 28030 46734 28082 46786
rect 29934 46734 29986 46786
rect 30270 46734 30322 46786
rect 37662 46734 37714 46786
rect 37998 46734 38050 46786
rect 43710 46734 43762 46786
rect 2270 46622 2322 46674
rect 3838 46622 3890 46674
rect 3950 46622 4002 46674
rect 6414 46622 6466 46674
rect 9102 46622 9154 46674
rect 9998 46622 10050 46674
rect 11230 46622 11282 46674
rect 12126 46622 12178 46674
rect 13470 46622 13522 46674
rect 13694 46622 13746 46674
rect 16606 46622 16658 46674
rect 16942 46622 16994 46674
rect 18062 46622 18114 46674
rect 18398 46622 18450 46674
rect 18622 46622 18674 46674
rect 19630 46622 19682 46674
rect 20078 46622 20130 46674
rect 20414 46622 20466 46674
rect 23438 46622 23490 46674
rect 24334 46622 24386 46674
rect 26910 46622 26962 46674
rect 27134 46622 27186 46674
rect 28142 46622 28194 46674
rect 28590 46622 28642 46674
rect 29486 46622 29538 46674
rect 30046 46622 30098 46674
rect 31278 46622 31330 46674
rect 37214 46622 37266 46674
rect 37438 46622 37490 46674
rect 37886 46622 37938 46674
rect 40014 46622 40066 46674
rect 40350 46622 40402 46674
rect 40574 46622 40626 46674
rect 44158 46622 44210 46674
rect 44606 46622 44658 46674
rect 56142 46622 56194 46674
rect 5070 46510 5122 46562
rect 5854 46510 5906 46562
rect 7534 46510 7586 46562
rect 11566 46510 11618 46562
rect 12462 46510 12514 46562
rect 12910 46510 12962 46562
rect 14478 46510 14530 46562
rect 14926 46510 14978 46562
rect 15374 46510 15426 46562
rect 15822 46510 15874 46562
rect 19742 46510 19794 46562
rect 21422 46510 21474 46562
rect 22206 46510 22258 46562
rect 23886 46510 23938 46562
rect 24782 46510 24834 46562
rect 25678 46510 25730 46562
rect 26686 46510 26738 46562
rect 31726 46510 31778 46562
rect 32062 46510 32114 46562
rect 33966 46510 34018 46562
rect 34862 46510 34914 46562
rect 35310 46510 35362 46562
rect 35758 46510 35810 46562
rect 55358 46510 55410 46562
rect 4174 46398 4226 46450
rect 5182 46398 5234 46450
rect 5742 46398 5794 46450
rect 6526 46398 6578 46450
rect 8094 46398 8146 46450
rect 10446 46398 10498 46450
rect 11006 46398 11058 46450
rect 11454 46398 11506 46450
rect 12910 46398 12962 46450
rect 14030 46398 14082 46450
rect 28366 46398 28418 46450
rect 29710 46398 29762 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 3614 46062 3666 46114
rect 17054 46062 17106 46114
rect 1934 45950 1986 46002
rect 2606 45950 2658 46002
rect 4510 45950 4562 46002
rect 9886 45950 9938 46002
rect 15150 45950 15202 46002
rect 3390 45838 3442 45890
rect 3838 45838 3890 45890
rect 4398 45838 4450 45890
rect 4622 45838 4674 45890
rect 4958 45838 5010 45890
rect 6302 45838 6354 45890
rect 6862 45838 6914 45890
rect 7982 45838 8034 45890
rect 8430 45838 8482 45890
rect 8990 45838 9042 45890
rect 9550 45838 9602 45890
rect 11006 45838 11058 45890
rect 11342 45838 11394 45890
rect 12686 45838 12738 45890
rect 13694 45838 13746 45890
rect 13918 45838 13970 45890
rect 16158 45838 16210 45890
rect 17054 45838 17106 45890
rect 2494 45726 2546 45778
rect 2718 45726 2770 45778
rect 10110 45726 10162 45778
rect 11230 45726 11282 45778
rect 14030 45726 14082 45778
rect 16718 45726 16770 45778
rect 17166 45726 17218 45778
rect 18398 46062 18450 46114
rect 20414 46062 20466 46114
rect 21870 46062 21922 46114
rect 22206 46062 22258 46114
rect 30270 46062 30322 46114
rect 30718 46062 30770 46114
rect 17950 45950 18002 46002
rect 18398 45950 18450 46002
rect 21870 45950 21922 46002
rect 27582 45950 27634 46002
rect 29486 45950 29538 46002
rect 30270 45950 30322 46002
rect 32958 45950 33010 46002
rect 39006 45950 39058 46002
rect 39678 45950 39730 46002
rect 44270 45950 44322 46002
rect 23438 45838 23490 45890
rect 25454 45838 25506 45890
rect 31390 45838 31442 45890
rect 31614 45838 31666 45890
rect 31838 45838 31890 45890
rect 34190 45838 34242 45890
rect 34526 45838 34578 45890
rect 36430 45838 36482 45890
rect 36766 45838 36818 45890
rect 39454 45838 39506 45890
rect 40126 45838 40178 45890
rect 44046 45838 44098 45890
rect 57374 45838 57426 45890
rect 18846 45726 18898 45778
rect 19518 45726 19570 45778
rect 19854 45726 19906 45778
rect 20526 45726 20578 45778
rect 20750 45726 20802 45778
rect 22430 45726 22482 45778
rect 23998 45726 24050 45778
rect 26014 45726 26066 45778
rect 33518 45726 33570 45778
rect 33630 45726 33682 45778
rect 34862 45726 34914 45778
rect 35310 45726 35362 45778
rect 39902 45726 39954 45778
rect 44382 45726 44434 45778
rect 57150 45726 57202 45778
rect 3726 45614 3778 45666
rect 5854 45614 5906 45666
rect 6750 45614 6802 45666
rect 6974 45614 7026 45666
rect 7422 45614 7474 45666
rect 12126 45614 12178 45666
rect 12798 45614 12850 45666
rect 13022 45614 13074 45666
rect 14478 45614 14530 45666
rect 15710 45614 15762 45666
rect 15934 45614 15986 45666
rect 16046 45614 16098 45666
rect 17502 45614 17554 45666
rect 22766 45614 22818 45666
rect 27022 45614 27074 45666
rect 28254 45614 28306 45666
rect 28702 45614 28754 45666
rect 30718 45614 30770 45666
rect 31726 45614 31778 45666
rect 32286 45614 32338 45666
rect 33854 45614 33906 45666
rect 34526 45614 34578 45666
rect 36542 45614 36594 45666
rect 37550 45614 37602 45666
rect 38334 45614 38386 45666
rect 56702 45614 56754 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 5294 45278 5346 45330
rect 13582 45278 13634 45330
rect 13694 45278 13746 45330
rect 14030 45278 14082 45330
rect 14254 45278 14306 45330
rect 20638 45278 20690 45330
rect 21534 45278 21586 45330
rect 23102 45278 23154 45330
rect 23662 45278 23714 45330
rect 28926 45278 28978 45330
rect 38110 45278 38162 45330
rect 38894 45278 38946 45330
rect 40126 45278 40178 45330
rect 4286 45166 4338 45218
rect 6974 45166 7026 45218
rect 8206 45166 8258 45218
rect 8878 45166 8930 45218
rect 9774 45166 9826 45218
rect 11454 45166 11506 45218
rect 15150 45166 15202 45218
rect 18846 45166 18898 45218
rect 18958 45166 19010 45218
rect 19742 45166 19794 45218
rect 21870 45166 21922 45218
rect 22766 45166 22818 45218
rect 27358 45166 27410 45218
rect 28030 45166 28082 45218
rect 31054 45166 31106 45218
rect 34302 45166 34354 45218
rect 37214 45166 37266 45218
rect 40014 45166 40066 45218
rect 43038 45166 43090 45218
rect 44494 45166 44546 45218
rect 2830 45054 2882 45106
rect 3950 45054 4002 45106
rect 5630 45054 5682 45106
rect 6862 45054 6914 45106
rect 7086 45054 7138 45106
rect 7534 45054 7586 45106
rect 8430 45054 8482 45106
rect 8654 45054 8706 45106
rect 10110 45054 10162 45106
rect 10894 45054 10946 45106
rect 11678 45054 11730 45106
rect 12014 45054 12066 45106
rect 13022 45054 13074 45106
rect 13358 45054 13410 45106
rect 14366 45054 14418 45106
rect 16942 45054 16994 45106
rect 19630 45054 19682 45106
rect 20750 45054 20802 45106
rect 21310 45054 21362 45106
rect 21758 45054 21810 45106
rect 24446 45054 24498 45106
rect 25790 45054 25842 45106
rect 25902 45054 25954 45106
rect 26126 45054 26178 45106
rect 26238 45054 26290 45106
rect 26686 45054 26738 45106
rect 27134 45054 27186 45106
rect 27918 45054 27970 45106
rect 28142 45054 28194 45106
rect 28590 45054 28642 45106
rect 29598 45054 29650 45106
rect 29934 45054 29986 45106
rect 32622 45054 32674 45106
rect 33630 45054 33682 45106
rect 34414 45054 34466 45106
rect 34526 45054 34578 45106
rect 34974 45054 35026 45106
rect 35534 45054 35586 45106
rect 35758 45054 35810 45106
rect 36654 45054 36706 45106
rect 36990 45054 37042 45106
rect 39566 45054 39618 45106
rect 39790 45054 39842 45106
rect 42702 45054 42754 45106
rect 43934 45054 43986 45106
rect 44158 45054 44210 45106
rect 1934 44942 1986 44994
rect 4174 44942 4226 44994
rect 4846 44942 4898 44994
rect 6302 44942 6354 44994
rect 8990 44942 9042 44994
rect 10334 44942 10386 44994
rect 11902 44942 11954 44994
rect 12574 44942 12626 44994
rect 15598 44942 15650 44994
rect 16046 44942 16098 44994
rect 16494 44942 16546 44994
rect 17950 44942 18002 44994
rect 21646 44942 21698 44994
rect 24222 44942 24274 44994
rect 26910 44942 26962 44994
rect 30494 44942 30546 44994
rect 31390 44942 31442 44994
rect 37662 44942 37714 44994
rect 39006 44942 39058 44994
rect 40462 44942 40514 44994
rect 44382 44942 44434 44994
rect 6078 44830 6130 44882
rect 6302 44830 6354 44882
rect 15262 44830 15314 44882
rect 15934 44830 15986 44882
rect 16494 44830 16546 44882
rect 17166 44830 17218 44882
rect 18958 44830 19010 44882
rect 24782 44830 24834 44882
rect 31278 44830 31330 44882
rect 32734 44830 32786 44882
rect 35982 44830 36034 44882
rect 36094 44830 36146 44882
rect 37326 44830 37378 44882
rect 38670 44830 38722 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 6302 44494 6354 44546
rect 10782 44494 10834 44546
rect 11566 44494 11618 44546
rect 12462 44494 12514 44546
rect 12910 44494 12962 44546
rect 15262 44494 15314 44546
rect 17390 44494 17442 44546
rect 20190 44494 20242 44546
rect 25790 44494 25842 44546
rect 26350 44494 26402 44546
rect 30718 44494 30770 44546
rect 31390 44494 31442 44546
rect 32958 44494 33010 44546
rect 38110 44494 38162 44546
rect 38334 44494 38386 44546
rect 39006 44494 39058 44546
rect 45502 44494 45554 44546
rect 2046 44382 2098 44434
rect 2494 44382 2546 44434
rect 6862 44382 6914 44434
rect 10782 44382 10834 44434
rect 18286 44382 18338 44434
rect 18846 44382 18898 44434
rect 25342 44382 25394 44434
rect 25902 44382 25954 44434
rect 26350 44382 26402 44434
rect 27134 44382 27186 44434
rect 31166 44382 31218 44434
rect 35646 44382 35698 44434
rect 40126 44382 40178 44434
rect 42366 44382 42418 44434
rect 43486 44382 43538 44434
rect 2942 44270 2994 44322
rect 6974 44270 7026 44322
rect 7534 44270 7586 44322
rect 8430 44270 8482 44322
rect 9214 44270 9266 44322
rect 9662 44270 9714 44322
rect 9774 44270 9826 44322
rect 12014 44270 12066 44322
rect 12238 44270 12290 44322
rect 15374 44270 15426 44322
rect 15598 44270 15650 44322
rect 18734 44270 18786 44322
rect 19294 44270 19346 44322
rect 21870 44270 21922 44322
rect 23214 44270 23266 44322
rect 23326 44270 23378 44322
rect 24110 44270 24162 44322
rect 28030 44270 28082 44322
rect 28590 44270 28642 44322
rect 29934 44270 29986 44322
rect 31950 44270 32002 44322
rect 32622 44270 32674 44322
rect 36206 44270 36258 44322
rect 36766 44270 36818 44322
rect 38558 44270 38610 44322
rect 39678 44270 39730 44322
rect 41022 44270 41074 44322
rect 41806 44270 41858 44322
rect 42814 44270 42866 44322
rect 43150 44270 43202 44322
rect 44046 44270 44098 44322
rect 44158 44270 44210 44322
rect 44270 44270 44322 44322
rect 44718 44270 44770 44322
rect 45502 44270 45554 44322
rect 4174 44158 4226 44210
rect 5742 44158 5794 44210
rect 6190 44158 6242 44210
rect 8094 44158 8146 44210
rect 9438 44158 9490 44210
rect 11790 44158 11842 44210
rect 13694 44158 13746 44210
rect 15710 44158 15762 44210
rect 16606 44158 16658 44210
rect 16718 44158 16770 44210
rect 17502 44158 17554 44210
rect 19854 44158 19906 44210
rect 20078 44158 20130 44210
rect 21982 44158 22034 44210
rect 22094 44158 22146 44210
rect 23102 44158 23154 44210
rect 23662 44158 23714 44210
rect 26686 44158 26738 44210
rect 27694 44158 27746 44210
rect 29598 44158 29650 44210
rect 32062 44158 32114 44210
rect 35534 44158 35586 44210
rect 35758 44158 35810 44210
rect 37886 44158 37938 44210
rect 45838 44158 45890 44210
rect 3278 44046 3330 44098
rect 3838 44046 3890 44098
rect 5070 44046 5122 44098
rect 5966 44046 6018 44098
rect 11342 44046 11394 44098
rect 14142 44046 14194 44098
rect 14590 44046 14642 44098
rect 16382 44046 16434 44098
rect 17390 44046 17442 44098
rect 18958 44046 19010 44098
rect 20638 44046 20690 44098
rect 22542 44046 22594 44098
rect 24558 44046 24610 44098
rect 28590 44046 28642 44098
rect 29710 44046 29762 44098
rect 30270 44046 30322 44098
rect 30718 44046 30770 44098
rect 33518 44046 33570 44098
rect 43374 44046 43426 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 4510 43710 4562 43762
rect 7870 43710 7922 43762
rect 9774 43710 9826 43762
rect 10782 43710 10834 43762
rect 12574 43710 12626 43762
rect 27582 43710 27634 43762
rect 28030 43710 28082 43762
rect 28254 43710 28306 43762
rect 29710 43710 29762 43762
rect 37214 43710 37266 43762
rect 37998 43710 38050 43762
rect 43934 43710 43986 43762
rect 46062 43710 46114 43762
rect 2830 43598 2882 43650
rect 3614 43598 3666 43650
rect 7646 43598 7698 43650
rect 7982 43598 8034 43650
rect 8542 43598 8594 43650
rect 13582 43598 13634 43650
rect 13694 43598 13746 43650
rect 15150 43598 15202 43650
rect 16718 43598 16770 43650
rect 18846 43598 18898 43650
rect 19966 43598 20018 43650
rect 20190 43598 20242 43650
rect 20638 43598 20690 43650
rect 22094 43598 22146 43650
rect 23438 43598 23490 43650
rect 24222 43598 24274 43650
rect 26350 43598 26402 43650
rect 27246 43598 27298 43650
rect 27358 43598 27410 43650
rect 28142 43598 28194 43650
rect 29374 43598 29426 43650
rect 39454 43598 39506 43650
rect 39902 43598 39954 43650
rect 40798 43598 40850 43650
rect 42590 43598 42642 43650
rect 43710 43598 43762 43650
rect 44046 43598 44098 43650
rect 46174 43598 46226 43650
rect 3278 43486 3330 43538
rect 4174 43486 4226 43538
rect 7422 43486 7474 43538
rect 11118 43486 11170 43538
rect 11902 43486 11954 43538
rect 12350 43486 12402 43538
rect 12462 43486 12514 43538
rect 13358 43486 13410 43538
rect 14030 43486 14082 43538
rect 14590 43486 14642 43538
rect 15038 43486 15090 43538
rect 15262 43486 15314 43538
rect 16382 43486 16434 43538
rect 16494 43486 16546 43538
rect 16942 43486 16994 43538
rect 17726 43486 17778 43538
rect 19406 43486 19458 43538
rect 19742 43486 19794 43538
rect 21534 43486 21586 43538
rect 22542 43486 22594 43538
rect 22990 43486 23042 43538
rect 23998 43486 24050 43538
rect 28702 43486 28754 43538
rect 34302 43486 34354 43538
rect 34526 43486 34578 43538
rect 34638 43486 34690 43538
rect 35086 43486 35138 43538
rect 35646 43486 35698 43538
rect 37662 43486 37714 43538
rect 38670 43486 38722 43538
rect 39230 43486 39282 43538
rect 41806 43486 41858 43538
rect 42366 43486 42418 43538
rect 42702 43486 42754 43538
rect 44158 43486 44210 43538
rect 44830 43486 44882 43538
rect 45054 43486 45106 43538
rect 45950 43486 46002 43538
rect 1934 43374 1986 43426
rect 2382 43374 2434 43426
rect 5182 43374 5234 43426
rect 5518 43374 5570 43426
rect 6078 43374 6130 43426
rect 6526 43374 6578 43426
rect 6974 43374 7026 43426
rect 8990 43374 9042 43426
rect 10222 43374 10274 43426
rect 12126 43374 12178 43426
rect 14142 43374 14194 43426
rect 15822 43374 15874 43426
rect 17054 43374 17106 43426
rect 18062 43374 18114 43426
rect 20078 43374 20130 43426
rect 21086 43374 21138 43426
rect 25006 43374 25058 43426
rect 25902 43374 25954 43426
rect 30158 43374 30210 43426
rect 30606 43374 30658 43426
rect 31166 43374 31218 43426
rect 31502 43374 31554 43426
rect 32062 43374 32114 43426
rect 32286 43374 32338 43426
rect 32622 43374 32674 43426
rect 33518 43374 33570 43426
rect 36654 43374 36706 43426
rect 40350 43374 40402 43426
rect 5182 43262 5234 43314
rect 6638 43262 6690 43314
rect 26014 43262 26066 43314
rect 26238 43262 26290 43314
rect 35870 43262 35922 43314
rect 36094 43262 36146 43314
rect 36206 43262 36258 43314
rect 38894 43262 38946 43314
rect 39342 43262 39394 43314
rect 39678 43262 39730 43314
rect 40350 43262 40402 43314
rect 43150 43262 43202 43314
rect 45390 43262 45442 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 4510 42926 4562 42978
rect 12686 42926 12738 42978
rect 14254 42926 14306 42978
rect 16382 42926 16434 42978
rect 17054 42926 17106 42978
rect 2606 42814 2658 42866
rect 3838 42814 3890 42866
rect 5630 42814 5682 42866
rect 8990 42814 9042 42866
rect 9886 42814 9938 42866
rect 16942 42814 16994 42866
rect 2382 42702 2434 42754
rect 2718 42702 2770 42754
rect 3614 42702 3666 42754
rect 4622 42702 4674 42754
rect 6414 42702 6466 42754
rect 6750 42702 6802 42754
rect 7534 42702 7586 42754
rect 10670 42702 10722 42754
rect 11342 42702 11394 42754
rect 12014 42702 12066 42754
rect 12126 42702 12178 42754
rect 14254 42702 14306 42754
rect 2158 42590 2210 42642
rect 6526 42590 6578 42642
rect 6638 42590 6690 42642
rect 7758 42590 7810 42642
rect 9550 42590 9602 42642
rect 10446 42590 10498 42642
rect 13694 42590 13746 42642
rect 13918 42590 13970 42642
rect 15822 42590 15874 42642
rect 18062 42926 18114 42978
rect 18286 42926 18338 42978
rect 18398 42926 18450 42978
rect 18958 42926 19010 42978
rect 26238 42926 26290 42978
rect 26686 42926 26738 42978
rect 27358 42926 27410 42978
rect 28030 42926 28082 42978
rect 39902 42926 39954 42978
rect 40350 42926 40402 42978
rect 43934 42926 43986 42978
rect 44158 42926 44210 42978
rect 19406 42814 19458 42866
rect 19742 42814 19794 42866
rect 20862 42814 20914 42866
rect 22990 42814 23042 42866
rect 26014 42814 26066 42866
rect 29486 42814 29538 42866
rect 29934 42814 29986 42866
rect 31726 42814 31778 42866
rect 34862 42814 34914 42866
rect 41022 42814 41074 42866
rect 43262 42814 43314 42866
rect 17950 42702 18002 42754
rect 19182 42702 19234 42754
rect 19854 42702 19906 42754
rect 25790 42702 25842 42754
rect 31502 42702 31554 42754
rect 31838 42702 31890 42754
rect 32062 42702 32114 42754
rect 34638 42702 34690 42754
rect 39678 42702 39730 42754
rect 40126 42702 40178 42754
rect 43710 42702 43762 42754
rect 44270 42702 44322 42754
rect 17838 42590 17890 42642
rect 22430 42590 22482 42642
rect 22542 42590 22594 42642
rect 22654 42590 22706 42642
rect 23662 42590 23714 42642
rect 23998 42590 24050 42642
rect 28254 42590 28306 42642
rect 28366 42590 28418 42642
rect 30494 42590 30546 42642
rect 30718 42590 30770 42642
rect 33070 42590 33122 42642
rect 34414 42590 34466 42642
rect 34974 42590 35026 42642
rect 35534 42590 35586 42642
rect 35758 42590 35810 42642
rect 35982 42590 36034 42642
rect 37774 42590 37826 42642
rect 38110 42590 38162 42642
rect 6302 42478 6354 42530
rect 8542 42478 8594 42530
rect 9774 42478 9826 42530
rect 14478 42478 14530 42530
rect 15374 42478 15426 42530
rect 16046 42478 16098 42530
rect 16270 42478 16322 42530
rect 17390 42478 17442 42530
rect 19630 42478 19682 42530
rect 20526 42478 20578 42530
rect 21646 42478 21698 42530
rect 22206 42478 22258 42530
rect 24446 42478 24498 42530
rect 25230 42478 25282 42530
rect 27358 42478 27410 42530
rect 27694 42478 27746 42530
rect 28590 42478 28642 42530
rect 30606 42478 30658 42530
rect 35422 42478 35474 42530
rect 38558 42478 38610 42530
rect 39006 42478 39058 42530
rect 40238 42478 40290 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 2830 42142 2882 42194
rect 3838 42142 3890 42194
rect 7310 42142 7362 42194
rect 8654 42142 8706 42194
rect 10782 42142 10834 42194
rect 10894 42142 10946 42194
rect 12126 42142 12178 42194
rect 12238 42142 12290 42194
rect 13134 42142 13186 42194
rect 15150 42142 15202 42194
rect 16606 42142 16658 42194
rect 23326 42142 23378 42194
rect 27582 42142 27634 42194
rect 30046 42142 30098 42194
rect 34190 42142 34242 42194
rect 34862 42142 34914 42194
rect 3166 42030 3218 42082
rect 4174 42030 4226 42082
rect 4846 42030 4898 42082
rect 5518 42030 5570 42082
rect 6862 42030 6914 42082
rect 7086 42030 7138 42082
rect 7422 42030 7474 42082
rect 8318 42030 8370 42082
rect 11006 42030 11058 42082
rect 14366 42030 14418 42082
rect 17726 42030 17778 42082
rect 25790 42030 25842 42082
rect 26014 42030 26066 42082
rect 26462 42030 26514 42082
rect 26686 42030 26738 42082
rect 26910 42030 26962 42082
rect 27022 42030 27074 42082
rect 29486 42030 29538 42082
rect 31838 42030 31890 42082
rect 31950 42030 32002 42082
rect 33742 42030 33794 42082
rect 33966 42030 34018 42082
rect 34302 42030 34354 42082
rect 35758 42030 35810 42082
rect 35870 42030 35922 42082
rect 36542 42030 36594 42082
rect 36878 42030 36930 42082
rect 37438 42030 37490 42082
rect 37774 42030 37826 42082
rect 40238 42030 40290 42082
rect 40686 42030 40738 42082
rect 4734 41918 4786 41970
rect 5966 41918 6018 41970
rect 6302 41918 6354 41970
rect 10334 41918 10386 41970
rect 14030 41918 14082 41970
rect 16046 41918 16098 41970
rect 16942 41918 16994 41970
rect 17950 41918 18002 41970
rect 18846 41918 18898 41970
rect 22094 41918 22146 41970
rect 22542 41918 22594 41970
rect 23102 41918 23154 41970
rect 23774 41918 23826 41970
rect 24670 41918 24722 41970
rect 25678 41918 25730 41970
rect 27806 41918 27858 41970
rect 28590 41918 28642 41970
rect 28814 41918 28866 41970
rect 30382 41918 30434 41970
rect 31614 41918 31666 41970
rect 32286 41918 32338 41970
rect 32846 41918 32898 41970
rect 35086 41918 35138 41970
rect 38670 41918 38722 41970
rect 38894 41918 38946 41970
rect 39118 41918 39170 41970
rect 40462 41918 40514 41970
rect 40798 41918 40850 41970
rect 41470 41918 41522 41970
rect 44158 41918 44210 41970
rect 44382 41918 44434 41970
rect 1934 41806 1986 41858
rect 2382 41806 2434 41858
rect 9886 41806 9938 41858
rect 11454 41806 11506 41858
rect 15598 41806 15650 41858
rect 18958 41806 19010 41858
rect 19966 41806 20018 41858
rect 20302 41806 20354 41858
rect 20750 41806 20802 41858
rect 21198 41806 21250 41858
rect 21758 41806 21810 41858
rect 23214 41806 23266 41858
rect 24558 41806 24610 41858
rect 31054 41806 31106 41858
rect 32398 41806 32450 41858
rect 9886 41694 9938 41746
rect 10222 41694 10274 41746
rect 12350 41694 12402 41746
rect 12910 41694 12962 41746
rect 13246 41694 13298 41746
rect 13918 41694 13970 41746
rect 14254 41694 14306 41746
rect 19070 41694 19122 41746
rect 20974 41694 21026 41746
rect 21758 41694 21810 41746
rect 35870 41694 35922 41746
rect 39342 41694 39394 41746
rect 39790 41694 39842 41746
rect 43486 41694 43538 41746
rect 43934 41694 43986 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 14030 41358 14082 41410
rect 17614 41358 17666 41410
rect 19854 41358 19906 41410
rect 21870 41358 21922 41410
rect 22206 41358 22258 41410
rect 25454 41358 25506 41410
rect 27582 41358 27634 41410
rect 39566 41358 39618 41410
rect 39790 41358 39842 41410
rect 2270 41246 2322 41298
rect 5966 41246 6018 41298
rect 7982 41246 8034 41298
rect 10670 41246 10722 41298
rect 13918 41246 13970 41298
rect 20638 41246 20690 41298
rect 24110 41246 24162 41298
rect 25230 41246 25282 41298
rect 26350 41246 26402 41298
rect 32846 41246 32898 41298
rect 35534 41246 35586 41298
rect 36318 41246 36370 41298
rect 38446 41246 38498 41298
rect 39006 41246 39058 41298
rect 55358 41246 55410 41298
rect 4622 41134 4674 41186
rect 7534 41134 7586 41186
rect 8430 41134 8482 41186
rect 9662 41134 9714 41186
rect 9886 41134 9938 41186
rect 10782 41134 10834 41186
rect 11790 41134 11842 41186
rect 12126 41134 12178 41186
rect 14030 41134 14082 41186
rect 14254 41134 14306 41186
rect 16494 41134 16546 41186
rect 17278 41134 17330 41186
rect 20078 41134 20130 41186
rect 20414 41134 20466 41186
rect 20750 41134 20802 41186
rect 22990 41134 23042 41186
rect 23774 41134 23826 41186
rect 28254 41134 28306 41186
rect 28478 41134 28530 41186
rect 29822 41134 29874 41186
rect 32174 41134 32226 41186
rect 32510 41134 32562 41186
rect 37774 41134 37826 41186
rect 39230 41134 39282 41186
rect 42926 41134 42978 41186
rect 43710 41134 43762 41186
rect 43822 41134 43874 41186
rect 45726 41134 45778 41186
rect 46062 41134 46114 41186
rect 56142 41134 56194 41186
rect 2494 41022 2546 41074
rect 3390 41022 3442 41074
rect 4062 41022 4114 41074
rect 4958 41022 5010 41074
rect 7310 41022 7362 41074
rect 11118 41022 11170 41074
rect 12014 41022 12066 41074
rect 16606 41022 16658 41074
rect 18846 41022 18898 41074
rect 19294 41022 19346 41074
rect 21646 41022 21698 41074
rect 24222 41022 24274 41074
rect 25790 41022 25842 41074
rect 27694 41022 27746 41074
rect 32286 41022 32338 41074
rect 37998 41022 38050 41074
rect 40462 41022 40514 41074
rect 40574 41022 40626 41074
rect 43038 41022 43090 41074
rect 44158 41022 44210 41074
rect 45502 41022 45554 41074
rect 2270 40910 2322 40962
rect 3054 40910 3106 40962
rect 12910 40910 12962 40962
rect 15486 40910 15538 40962
rect 15934 40910 15986 40962
rect 18510 40910 18562 40962
rect 20526 40910 20578 40962
rect 23102 40910 23154 40962
rect 27134 40910 27186 40962
rect 28814 40910 28866 40962
rect 29598 40910 29650 40962
rect 29710 40910 29762 40962
rect 30046 40910 30098 40962
rect 30606 40910 30658 40962
rect 31054 40910 31106 40962
rect 39902 40910 39954 40962
rect 40798 40910 40850 40962
rect 43262 40910 43314 40962
rect 43934 40910 43986 40962
rect 45726 40910 45778 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 1822 40574 1874 40626
rect 8766 40574 8818 40626
rect 8878 40574 8930 40626
rect 10110 40574 10162 40626
rect 10670 40574 10722 40626
rect 12238 40574 12290 40626
rect 13134 40574 13186 40626
rect 13694 40574 13746 40626
rect 16606 40574 16658 40626
rect 17614 40574 17666 40626
rect 17838 40574 17890 40626
rect 20414 40574 20466 40626
rect 21422 40574 21474 40626
rect 21982 40574 22034 40626
rect 24110 40574 24162 40626
rect 24558 40574 24610 40626
rect 26350 40574 26402 40626
rect 26798 40574 26850 40626
rect 27358 40574 27410 40626
rect 28030 40574 28082 40626
rect 28478 40574 28530 40626
rect 28926 40574 28978 40626
rect 34974 40574 35026 40626
rect 36542 40574 36594 40626
rect 38670 40574 38722 40626
rect 40014 40574 40066 40626
rect 40798 40574 40850 40626
rect 43934 40574 43986 40626
rect 44942 40574 44994 40626
rect 2942 40462 2994 40514
rect 7086 40462 7138 40514
rect 8430 40462 8482 40514
rect 12910 40462 12962 40514
rect 17950 40462 18002 40514
rect 20078 40462 20130 40514
rect 22430 40462 22482 40514
rect 23438 40462 23490 40514
rect 29374 40462 29426 40514
rect 31166 40462 31218 40514
rect 33966 40462 34018 40514
rect 34638 40462 34690 40514
rect 37774 40462 37826 40514
rect 43710 40462 43762 40514
rect 44494 40462 44546 40514
rect 2270 40350 2322 40402
rect 3950 40350 4002 40402
rect 4510 40350 4562 40402
rect 5854 40350 5906 40402
rect 8542 40350 8594 40402
rect 8990 40350 9042 40402
rect 9774 40350 9826 40402
rect 11230 40350 11282 40402
rect 11566 40350 11618 40402
rect 12798 40350 12850 40402
rect 15374 40350 15426 40402
rect 15822 40350 15874 40402
rect 16942 40350 16994 40402
rect 19070 40350 19122 40402
rect 20414 40350 20466 40402
rect 20638 40350 20690 40402
rect 22094 40350 22146 40402
rect 22206 40350 22258 40402
rect 23102 40350 23154 40402
rect 23550 40350 23602 40402
rect 23662 40350 23714 40402
rect 29598 40350 29650 40402
rect 29822 40350 29874 40402
rect 33854 40350 33906 40402
rect 36878 40350 36930 40402
rect 37438 40350 37490 40402
rect 41582 40350 41634 40402
rect 41806 40350 41858 40402
rect 42142 40350 42194 40402
rect 43598 40350 43650 40402
rect 44382 40350 44434 40402
rect 45390 40350 45442 40402
rect 46622 40350 46674 40402
rect 46846 40350 46898 40402
rect 3054 40238 3106 40290
rect 7198 40238 7250 40290
rect 14590 40238 14642 40290
rect 15150 40238 15202 40290
rect 18734 40238 18786 40290
rect 19518 40238 19570 40290
rect 26014 40238 26066 40290
rect 29486 40238 29538 40290
rect 45166 40238 45218 40290
rect 47518 40238 47570 40290
rect 7310 40126 7362 40178
rect 11118 40126 11170 40178
rect 11454 40126 11506 40178
rect 13582 40126 13634 40178
rect 13918 40126 13970 40178
rect 23886 40126 23938 40178
rect 24222 40126 24274 40178
rect 26126 40126 26178 40178
rect 27246 40126 27298 40178
rect 33966 40126 34018 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 7534 39790 7586 39842
rect 7758 39790 7810 39842
rect 14254 39790 14306 39842
rect 16942 39790 16994 39842
rect 17502 39790 17554 39842
rect 19854 39790 19906 39842
rect 20190 39790 20242 39842
rect 22094 39790 22146 39842
rect 23102 39790 23154 39842
rect 30942 39790 30994 39842
rect 37550 39790 37602 39842
rect 3726 39678 3778 39730
rect 5966 39678 6018 39730
rect 7534 39678 7586 39730
rect 8990 39678 9042 39730
rect 10446 39678 10498 39730
rect 12462 39678 12514 39730
rect 12910 39678 12962 39730
rect 15038 39678 15090 39730
rect 21646 39678 21698 39730
rect 24222 39678 24274 39730
rect 25006 39678 25058 39730
rect 25454 39678 25506 39730
rect 25902 39678 25954 39730
rect 33630 39678 33682 39730
rect 36878 39678 36930 39730
rect 37662 39678 37714 39730
rect 40686 39678 40738 39730
rect 43710 39678 43762 39730
rect 43934 39678 43986 39730
rect 2830 39566 2882 39618
rect 3502 39566 3554 39618
rect 3838 39566 3890 39618
rect 4174 39566 4226 39618
rect 7982 39566 8034 39618
rect 9550 39566 9602 39618
rect 9998 39566 10050 39618
rect 10222 39566 10274 39618
rect 11118 39566 11170 39618
rect 11342 39566 11394 39618
rect 11678 39566 11730 39618
rect 13918 39566 13970 39618
rect 14254 39566 14306 39618
rect 17054 39566 17106 39618
rect 17726 39566 17778 39618
rect 18398 39566 18450 39618
rect 21870 39566 21922 39618
rect 22542 39566 22594 39618
rect 22990 39566 23042 39618
rect 26462 39566 26514 39618
rect 27246 39566 27298 39618
rect 27694 39566 27746 39618
rect 31502 39566 31554 39618
rect 32622 39566 32674 39618
rect 33742 39566 33794 39618
rect 34190 39566 34242 39618
rect 38894 39566 38946 39618
rect 39342 39566 39394 39618
rect 40574 39566 40626 39618
rect 42030 39566 42082 39618
rect 44046 39566 44098 39618
rect 47518 39566 47570 39618
rect 57374 39566 57426 39618
rect 1934 39454 1986 39506
rect 6862 39454 6914 39506
rect 8318 39454 8370 39506
rect 9102 39454 9154 39506
rect 10558 39454 10610 39506
rect 13694 39454 13746 39506
rect 15934 39454 15986 39506
rect 18734 39454 18786 39506
rect 19630 39454 19682 39506
rect 26686 39454 26738 39506
rect 27806 39454 27858 39506
rect 30830 39454 30882 39506
rect 31838 39454 31890 39506
rect 42478 39454 42530 39506
rect 57150 39454 57202 39506
rect 4958 39342 5010 39394
rect 6526 39342 6578 39394
rect 8878 39342 8930 39394
rect 11230 39342 11282 39394
rect 14478 39342 14530 39394
rect 15598 39342 15650 39394
rect 16494 39342 16546 39394
rect 17838 39342 17890 39394
rect 20974 39342 21026 39394
rect 23102 39342 23154 39394
rect 23774 39342 23826 39394
rect 28366 39342 28418 39394
rect 28814 39342 28866 39394
rect 29934 39342 29986 39394
rect 30382 39342 30434 39394
rect 32398 39342 32450 39394
rect 35086 39342 35138 39394
rect 38110 39342 38162 39394
rect 39230 39342 39282 39394
rect 39454 39342 39506 39394
rect 47854 39342 47906 39394
rect 56702 39342 56754 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 2158 39006 2210 39058
rect 7758 39006 7810 39058
rect 8094 39006 8146 39058
rect 9998 39006 10050 39058
rect 12350 39006 12402 39058
rect 12574 39006 12626 39058
rect 13358 39006 13410 39058
rect 15710 39006 15762 39058
rect 30046 39006 30098 39058
rect 30494 39006 30546 39058
rect 38894 39006 38946 39058
rect 39454 39006 39506 39058
rect 41694 39006 41746 39058
rect 41918 39006 41970 39058
rect 42814 39006 42866 39058
rect 3838 38894 3890 38946
rect 6078 38894 6130 38946
rect 7982 38894 8034 38946
rect 10110 38894 10162 38946
rect 10782 38894 10834 38946
rect 11118 38894 11170 38946
rect 14254 38894 14306 38946
rect 14590 38894 14642 38946
rect 16382 38894 16434 38946
rect 16494 38894 16546 38946
rect 23214 38894 23266 38946
rect 27806 38894 27858 38946
rect 28702 38894 28754 38946
rect 32510 38894 32562 38946
rect 34638 38894 34690 38946
rect 36990 38894 37042 38946
rect 37214 38894 37266 38946
rect 38334 38894 38386 38946
rect 41582 38894 41634 38946
rect 42478 38894 42530 38946
rect 42590 38894 42642 38946
rect 1934 38782 1986 38834
rect 3166 38782 3218 38834
rect 5742 38782 5794 38834
rect 6302 38782 6354 38834
rect 6750 38782 6802 38834
rect 7422 38782 7474 38834
rect 8654 38782 8706 38834
rect 12686 38782 12738 38834
rect 13694 38782 13746 38834
rect 16158 38782 16210 38834
rect 16942 38782 16994 38834
rect 17726 38782 17778 38834
rect 18062 38782 18114 38834
rect 19630 38782 19682 38834
rect 20750 38782 20802 38834
rect 23774 38782 23826 38834
rect 24222 38782 24274 38834
rect 24558 38782 24610 38834
rect 25790 38782 25842 38834
rect 27358 38782 27410 38834
rect 27694 38782 27746 38834
rect 28366 38782 28418 38834
rect 28478 38782 28530 38834
rect 28814 38782 28866 38834
rect 31054 38782 31106 38834
rect 32622 38782 32674 38834
rect 35534 38782 35586 38834
rect 36206 38782 36258 38834
rect 36878 38782 36930 38834
rect 40014 38782 40066 38834
rect 2830 38670 2882 38722
rect 4286 38670 4338 38722
rect 5182 38670 5234 38722
rect 9102 38670 9154 38722
rect 9886 38670 9938 38722
rect 12014 38670 12066 38722
rect 15262 38670 15314 38722
rect 21422 38670 21474 38722
rect 22654 38670 22706 38722
rect 24670 38670 24722 38722
rect 26350 38670 26402 38722
rect 29598 38670 29650 38722
rect 31390 38670 31442 38722
rect 34190 38670 34242 38722
rect 37662 38670 37714 38722
rect 39566 38670 39618 38722
rect 40462 38670 40514 38722
rect 21646 38558 21698 38610
rect 31278 38558 31330 38610
rect 38558 38558 38610 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 1822 38222 1874 38274
rect 2270 38222 2322 38274
rect 2606 38222 2658 38274
rect 23662 38222 23714 38274
rect 24222 38222 24274 38274
rect 24558 38222 24610 38274
rect 26686 38222 26738 38274
rect 31054 38222 31106 38274
rect 31502 38222 31554 38274
rect 32286 38222 32338 38274
rect 34190 38222 34242 38274
rect 34526 38222 34578 38274
rect 35086 38222 35138 38274
rect 1934 38110 1986 38162
rect 3278 38110 3330 38162
rect 5070 38110 5122 38162
rect 9998 38110 10050 38162
rect 14478 38110 14530 38162
rect 18622 38110 18674 38162
rect 18734 38110 18786 38162
rect 20638 38110 20690 38162
rect 22094 38110 22146 38162
rect 23214 38110 23266 38162
rect 23438 38110 23490 38162
rect 24110 38110 24162 38162
rect 28814 38110 28866 38162
rect 31950 38110 32002 38162
rect 33518 38110 33570 38162
rect 34526 38110 34578 38162
rect 34974 38110 35026 38162
rect 36766 38110 36818 38162
rect 37998 38110 38050 38162
rect 41918 38110 41970 38162
rect 2830 37998 2882 38050
rect 5854 37998 5906 38050
rect 7086 37998 7138 38050
rect 7534 37998 7586 38050
rect 9102 37998 9154 38050
rect 11790 37998 11842 38050
rect 14030 37998 14082 38050
rect 14926 37998 14978 38050
rect 20302 37998 20354 38050
rect 24446 37998 24498 38050
rect 25566 37998 25618 38050
rect 26574 37998 26626 38050
rect 27358 37998 27410 38050
rect 27582 37998 27634 38050
rect 29598 37998 29650 38050
rect 30046 37998 30098 38050
rect 30606 37998 30658 38050
rect 30830 37998 30882 38050
rect 33070 37998 33122 38050
rect 33966 37998 34018 38050
rect 39454 37998 39506 38050
rect 42142 37998 42194 38050
rect 42366 37998 42418 38050
rect 2382 37886 2434 37938
rect 4286 37886 4338 37938
rect 6414 37886 6466 37938
rect 10110 37886 10162 37938
rect 12686 37886 12738 37938
rect 14366 37886 14418 37938
rect 16046 37886 16098 37938
rect 16494 37886 16546 37938
rect 16942 37886 16994 37938
rect 17502 37886 17554 37938
rect 19294 37886 19346 37938
rect 19630 37886 19682 37938
rect 20862 37886 20914 37938
rect 21646 37886 21698 37938
rect 22654 37886 22706 37938
rect 28254 37886 28306 37938
rect 32062 37886 32114 37938
rect 32958 37886 33010 37938
rect 38222 37886 38274 37938
rect 40126 37886 40178 37938
rect 41582 37886 41634 37938
rect 41806 37886 41858 37938
rect 3950 37774 4002 37826
rect 5854 37774 5906 37826
rect 11230 37774 11282 37826
rect 12350 37774 12402 37826
rect 15710 37774 15762 37826
rect 17838 37774 17890 37826
rect 18510 37774 18562 37826
rect 24894 37774 24946 37826
rect 25790 37774 25842 37826
rect 26462 37774 26514 37826
rect 32734 37774 32786 37826
rect 41134 37774 41186 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 2158 37438 2210 37490
rect 3838 37438 3890 37490
rect 4398 37438 4450 37490
rect 9886 37438 9938 37490
rect 14702 37438 14754 37490
rect 16942 37438 16994 37490
rect 21534 37438 21586 37490
rect 22206 37438 22258 37490
rect 22542 37438 22594 37490
rect 27246 37438 27298 37490
rect 27806 37438 27858 37490
rect 37550 37438 37602 37490
rect 38670 37438 38722 37490
rect 1822 37326 1874 37378
rect 7198 37326 7250 37378
rect 8990 37326 9042 37378
rect 10558 37326 10610 37378
rect 14478 37326 14530 37378
rect 21422 37326 21474 37378
rect 21646 37326 21698 37378
rect 23214 37326 23266 37378
rect 34414 37326 34466 37378
rect 34750 37326 34802 37378
rect 35422 37326 35474 37378
rect 2718 37214 2770 37266
rect 3278 37214 3330 37266
rect 4286 37214 4338 37266
rect 4510 37214 4562 37266
rect 4846 37214 4898 37266
rect 5742 37214 5794 37266
rect 6302 37214 6354 37266
rect 6974 37214 7026 37266
rect 7422 37214 7474 37266
rect 8766 37214 8818 37266
rect 10894 37214 10946 37266
rect 12238 37214 12290 37266
rect 14254 37214 14306 37266
rect 15150 37214 15202 37266
rect 15374 37214 15426 37266
rect 16606 37214 16658 37266
rect 18398 37214 18450 37266
rect 18622 37214 18674 37266
rect 20078 37214 20130 37266
rect 23550 37214 23602 37266
rect 24222 37214 24274 37266
rect 26238 37214 26290 37266
rect 26686 37214 26738 37266
rect 28142 37214 28194 37266
rect 29598 37214 29650 37266
rect 30606 37214 30658 37266
rect 31950 37214 32002 37266
rect 32398 37214 32450 37266
rect 35646 37214 35698 37266
rect 35870 37214 35922 37266
rect 38110 37214 38162 37266
rect 38334 37214 38386 37266
rect 42478 37214 42530 37266
rect 42814 37214 42866 37266
rect 17726 37102 17778 37154
rect 18846 37102 18898 37154
rect 19630 37102 19682 37154
rect 23774 37102 23826 37154
rect 24782 37102 24834 37154
rect 25678 37102 25730 37154
rect 29150 37102 29202 37154
rect 30046 37102 30098 37154
rect 32846 37102 32898 37154
rect 33966 37102 34018 37154
rect 35758 37102 35810 37154
rect 41806 37102 41858 37154
rect 42366 37102 42418 37154
rect 6862 36990 6914 37042
rect 7646 36990 7698 37042
rect 15710 36990 15762 37042
rect 19070 36990 19122 37042
rect 26910 36990 26962 37042
rect 30830 36990 30882 37042
rect 31166 36990 31218 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 2270 36654 2322 36706
rect 4062 36654 4114 36706
rect 9886 36654 9938 36706
rect 12574 36654 12626 36706
rect 27694 36654 27746 36706
rect 28478 36654 28530 36706
rect 31278 36654 31330 36706
rect 41470 36654 41522 36706
rect 1822 36542 1874 36594
rect 6078 36542 6130 36594
rect 6974 36542 7026 36594
rect 7982 36542 8034 36594
rect 9214 36542 9266 36594
rect 10894 36542 10946 36594
rect 26238 36542 26290 36594
rect 27358 36542 27410 36594
rect 28814 36542 28866 36594
rect 31390 36542 31442 36594
rect 31950 36542 32002 36594
rect 34862 36542 34914 36594
rect 38670 36542 38722 36594
rect 40798 36542 40850 36594
rect 42366 36542 42418 36594
rect 43150 36542 43202 36594
rect 4510 36430 4562 36482
rect 4734 36430 4786 36482
rect 4958 36430 5010 36482
rect 7422 36430 7474 36482
rect 8094 36430 8146 36482
rect 10558 36430 10610 36482
rect 11678 36430 11730 36482
rect 12350 36430 12402 36482
rect 12910 36430 12962 36482
rect 13806 36430 13858 36482
rect 15598 36430 15650 36482
rect 16270 36430 16322 36482
rect 17166 36430 17218 36482
rect 19854 36430 19906 36482
rect 21982 36430 22034 36482
rect 22542 36430 22594 36482
rect 22878 36430 22930 36482
rect 26910 36430 26962 36482
rect 29598 36430 29650 36482
rect 30494 36430 30546 36482
rect 33630 36430 33682 36482
rect 34638 36430 34690 36482
rect 35982 36430 36034 36482
rect 40126 36430 40178 36482
rect 41358 36430 41410 36482
rect 42478 36430 42530 36482
rect 2382 36318 2434 36370
rect 2942 36318 2994 36370
rect 3278 36318 3330 36370
rect 8318 36318 8370 36370
rect 9774 36318 9826 36370
rect 10670 36318 10722 36370
rect 14030 36318 14082 36370
rect 14254 36318 14306 36370
rect 14478 36318 14530 36370
rect 15486 36318 15538 36370
rect 16158 36318 16210 36370
rect 18510 36318 18562 36370
rect 19630 36318 19682 36370
rect 20526 36318 20578 36370
rect 21646 36318 21698 36370
rect 21758 36318 21810 36370
rect 23326 36318 23378 36370
rect 23662 36318 23714 36370
rect 24222 36318 24274 36370
rect 24558 36318 24610 36370
rect 28702 36318 28754 36370
rect 29710 36318 29762 36370
rect 33182 36318 33234 36370
rect 33742 36318 33794 36370
rect 36766 36318 36818 36370
rect 39118 36318 39170 36370
rect 6414 36206 6466 36258
rect 9886 36206 9938 36258
rect 17726 36206 17778 36258
rect 18174 36206 18226 36258
rect 19070 36206 19122 36258
rect 20638 36206 20690 36258
rect 20862 36206 20914 36258
rect 22654 36206 22706 36258
rect 25006 36206 25058 36258
rect 25454 36206 25506 36258
rect 30606 36206 30658 36258
rect 33966 36206 34018 36258
rect 41470 36206 41522 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 1822 35870 1874 35922
rect 2270 35870 2322 35922
rect 3950 35870 4002 35922
rect 4734 35870 4786 35922
rect 8206 35870 8258 35922
rect 14590 35870 14642 35922
rect 16606 35870 16658 35922
rect 21646 35870 21698 35922
rect 22430 35870 22482 35922
rect 23214 35870 23266 35922
rect 23774 35870 23826 35922
rect 26014 35870 26066 35922
rect 27246 35870 27298 35922
rect 27358 35870 27410 35922
rect 27918 35870 27970 35922
rect 32958 35870 33010 35922
rect 34190 35870 34242 35922
rect 35086 35870 35138 35922
rect 35758 35870 35810 35922
rect 36094 35870 36146 35922
rect 37214 35870 37266 35922
rect 38446 35870 38498 35922
rect 39006 35870 39058 35922
rect 39118 35870 39170 35922
rect 41694 35870 41746 35922
rect 41806 35870 41858 35922
rect 54350 35870 54402 35922
rect 3614 35758 3666 35810
rect 4174 35758 4226 35810
rect 5294 35758 5346 35810
rect 8878 35758 8930 35810
rect 11006 35758 11058 35810
rect 11902 35758 11954 35810
rect 12798 35758 12850 35810
rect 13246 35758 13298 35810
rect 17726 35758 17778 35810
rect 20638 35758 20690 35810
rect 21534 35758 21586 35810
rect 27470 35758 27522 35810
rect 32734 35758 32786 35810
rect 35870 35758 35922 35810
rect 39230 35758 39282 35810
rect 41582 35758 41634 35810
rect 3054 35646 3106 35698
rect 3838 35646 3890 35698
rect 5630 35646 5682 35698
rect 6302 35646 6354 35698
rect 6750 35646 6802 35698
rect 8654 35646 8706 35698
rect 8766 35646 8818 35698
rect 10334 35646 10386 35698
rect 11454 35646 11506 35698
rect 12462 35646 12514 35698
rect 13470 35646 13522 35698
rect 14030 35646 14082 35698
rect 14926 35646 14978 35698
rect 16942 35646 16994 35698
rect 18286 35646 18338 35698
rect 18958 35646 19010 35698
rect 19294 35646 19346 35698
rect 19406 35646 19458 35698
rect 20862 35646 20914 35698
rect 21870 35646 21922 35698
rect 22654 35646 22706 35698
rect 23998 35646 24050 35698
rect 29038 35646 29090 35698
rect 29486 35646 29538 35698
rect 32622 35646 32674 35698
rect 33630 35646 33682 35698
rect 33854 35646 33906 35698
rect 34862 35646 34914 35698
rect 34974 35646 35026 35698
rect 35422 35646 35474 35698
rect 36318 35646 36370 35698
rect 54910 35646 54962 35698
rect 7198 35534 7250 35586
rect 7646 35534 7698 35586
rect 9774 35534 9826 35586
rect 11342 35534 11394 35586
rect 15598 35534 15650 35586
rect 16046 35534 16098 35586
rect 24670 35534 24722 35586
rect 25566 35534 25618 35586
rect 28590 35534 28642 35586
rect 30046 35534 30098 35586
rect 30718 35534 30770 35586
rect 56030 35534 56082 35586
rect 2718 35422 2770 35474
rect 3054 35422 3106 35474
rect 7198 35422 7250 35474
rect 7870 35422 7922 35474
rect 19966 35422 20018 35474
rect 24782 35422 24834 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 9102 35086 9154 35138
rect 11566 35086 11618 35138
rect 28590 35086 28642 35138
rect 37550 35086 37602 35138
rect 5630 34974 5682 35026
rect 6638 34974 6690 35026
rect 7310 34974 7362 35026
rect 9326 34974 9378 35026
rect 11454 34974 11506 35026
rect 12574 34974 12626 35026
rect 15710 34974 15762 35026
rect 25230 34974 25282 35026
rect 26350 34974 26402 35026
rect 26910 34974 26962 35026
rect 27918 34974 27970 35026
rect 32062 34974 32114 35026
rect 34526 34974 34578 35026
rect 35646 34974 35698 35026
rect 37774 34974 37826 35026
rect 2158 34862 2210 34914
rect 3838 34862 3890 34914
rect 4734 34862 4786 34914
rect 6190 34862 6242 34914
rect 10334 34862 10386 34914
rect 11118 34862 11170 34914
rect 12910 34862 12962 34914
rect 14926 34862 14978 34914
rect 16942 34862 16994 34914
rect 17838 34862 17890 34914
rect 18286 34862 18338 34914
rect 19182 34862 19234 34914
rect 20862 34862 20914 34914
rect 24670 34862 24722 34914
rect 25790 34862 25842 34914
rect 26574 34862 26626 34914
rect 28478 34862 28530 34914
rect 29934 34862 29986 34914
rect 31390 34862 31442 34914
rect 31838 34862 31890 34914
rect 32510 34862 32562 34914
rect 39902 34862 39954 34914
rect 40462 34862 40514 34914
rect 7870 34750 7922 34802
rect 8206 34750 8258 34802
rect 8766 34750 8818 34802
rect 10558 34750 10610 34802
rect 13694 34750 13746 34802
rect 14030 34750 14082 34802
rect 15150 34750 15202 34802
rect 15822 34750 15874 34802
rect 16606 34750 16658 34802
rect 16718 34750 16770 34802
rect 17502 34750 17554 34802
rect 18398 34750 18450 34802
rect 20526 34750 20578 34802
rect 23886 34750 23938 34802
rect 24782 34750 24834 34802
rect 29598 34750 29650 34802
rect 2606 34638 2658 34690
rect 2942 34638 2994 34690
rect 3502 34638 3554 34690
rect 4958 34638 5010 34690
rect 18510 34638 18562 34690
rect 21534 34638 21586 34690
rect 30606 34638 30658 34690
rect 33742 34638 33794 34690
rect 36766 34638 36818 34690
rect 37774 34638 37826 34690
rect 39006 34638 39058 34690
rect 39454 34638 39506 34690
rect 43038 34638 43090 34690
rect 43598 34638 43650 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 4398 34302 4450 34354
rect 4958 34302 5010 34354
rect 5406 34302 5458 34354
rect 5742 34302 5794 34354
rect 6302 34302 6354 34354
rect 8430 34302 8482 34354
rect 9886 34302 9938 34354
rect 10334 34302 10386 34354
rect 10782 34302 10834 34354
rect 11230 34302 11282 34354
rect 11678 34302 11730 34354
rect 12126 34302 12178 34354
rect 12574 34302 12626 34354
rect 14030 34302 14082 34354
rect 14926 34302 14978 34354
rect 15710 34302 15762 34354
rect 16158 34302 16210 34354
rect 16942 34302 16994 34354
rect 19294 34302 19346 34354
rect 21086 34302 21138 34354
rect 21646 34302 21698 34354
rect 22766 34302 22818 34354
rect 24222 34302 24274 34354
rect 25566 34302 25618 34354
rect 28254 34302 28306 34354
rect 29262 34302 29314 34354
rect 29710 34302 29762 34354
rect 31726 34302 31778 34354
rect 32734 34302 32786 34354
rect 3950 34190 4002 34242
rect 7646 34190 7698 34242
rect 17950 34190 18002 34242
rect 18622 34190 18674 34242
rect 18734 34190 18786 34242
rect 18846 34190 18898 34242
rect 23102 34190 23154 34242
rect 23886 34190 23938 34242
rect 24446 34190 24498 34242
rect 32622 34190 32674 34242
rect 34078 34190 34130 34242
rect 37102 34190 37154 34242
rect 2830 34078 2882 34130
rect 3726 34078 3778 34130
rect 6862 34078 6914 34130
rect 7982 34078 8034 34130
rect 13470 34078 13522 34130
rect 13806 34078 13858 34130
rect 14590 34078 14642 34130
rect 16494 34078 16546 34130
rect 19742 34078 19794 34130
rect 20750 34078 20802 34130
rect 21870 34078 21922 34130
rect 22430 34078 22482 34130
rect 22766 34078 22818 34130
rect 24670 34078 24722 34130
rect 27806 34078 27858 34130
rect 29934 34078 29986 34130
rect 30382 34078 30434 34130
rect 32958 34078 33010 34130
rect 1934 33966 1986 34018
rect 8878 33966 8930 34018
rect 13022 33966 13074 34018
rect 20190 33966 20242 34018
rect 26014 33966 26066 34018
rect 28702 33966 28754 34018
rect 29822 33966 29874 34018
rect 31166 33966 31218 34018
rect 31614 33966 31666 34018
rect 36318 33966 36370 34018
rect 38222 33966 38274 34018
rect 6638 33854 6690 33906
rect 14142 33854 14194 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 3726 33518 3778 33570
rect 6638 33518 6690 33570
rect 9550 33518 9602 33570
rect 9886 33518 9938 33570
rect 11230 33518 11282 33570
rect 11790 33518 11842 33570
rect 17278 33518 17330 33570
rect 23886 33518 23938 33570
rect 24670 33518 24722 33570
rect 28926 33518 28978 33570
rect 31726 33518 31778 33570
rect 36878 33518 36930 33570
rect 1934 33406 1986 33458
rect 2382 33406 2434 33458
rect 4622 33406 4674 33458
rect 5742 33406 5794 33458
rect 8094 33406 8146 33458
rect 10558 33406 10610 33458
rect 11006 33406 11058 33458
rect 11454 33406 11506 33458
rect 11902 33406 11954 33458
rect 14366 33406 14418 33458
rect 18734 33406 18786 33458
rect 20414 33406 20466 33458
rect 22094 33406 22146 33458
rect 44494 33406 44546 33458
rect 2942 33294 2994 33346
rect 8878 33294 8930 33346
rect 12910 33294 12962 33346
rect 14926 33294 14978 33346
rect 15934 33294 15986 33346
rect 16718 33294 16770 33346
rect 16942 33294 16994 33346
rect 23438 33294 23490 33346
rect 23774 33294 23826 33346
rect 25454 33294 25506 33346
rect 25902 33294 25954 33346
rect 29710 33294 29762 33346
rect 30046 33294 30098 33346
rect 30382 33294 30434 33346
rect 31054 33294 31106 33346
rect 32734 33294 32786 33346
rect 33406 33294 33458 33346
rect 33854 33294 33906 33346
rect 37662 33294 37714 33346
rect 37998 33294 38050 33346
rect 41470 33294 41522 33346
rect 3166 33182 3218 33234
rect 3838 33182 3890 33234
rect 5854 33182 5906 33234
rect 6750 33182 6802 33234
rect 7310 33182 7362 33234
rect 7422 33182 7474 33234
rect 8990 33182 9042 33234
rect 13694 33182 13746 33234
rect 13806 33182 13858 33234
rect 16158 33182 16210 33234
rect 17838 33182 17890 33234
rect 18174 33182 18226 33234
rect 21646 33182 21698 33234
rect 22654 33182 22706 33234
rect 22766 33182 22818 33234
rect 31838 33182 31890 33234
rect 42366 33182 42418 33234
rect 7646 33070 7698 33122
rect 12238 33070 12290 33122
rect 14030 33070 14082 33122
rect 15262 33070 15314 33122
rect 19294 33070 19346 33122
rect 20862 33070 20914 33122
rect 22990 33070 23042 33122
rect 23550 33070 23602 33122
rect 24110 33070 24162 33122
rect 24558 33070 24610 33122
rect 28254 33070 28306 33122
rect 29822 33070 29874 33122
rect 30830 33070 30882 33122
rect 30942 33070 30994 33122
rect 31726 33070 31778 33122
rect 32398 33070 32450 33122
rect 36318 33070 36370 33122
rect 40350 33070 40402 33122
rect 41134 33070 41186 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 1934 32734 1986 32786
rect 6078 32734 6130 32786
rect 6414 32734 6466 32786
rect 7198 32734 7250 32786
rect 11006 32734 11058 32786
rect 11230 32734 11282 32786
rect 11678 32734 11730 32786
rect 13134 32734 13186 32786
rect 14142 32734 14194 32786
rect 15150 32734 15202 32786
rect 17614 32734 17666 32786
rect 18174 32734 18226 32786
rect 22094 32734 22146 32786
rect 24110 32734 24162 32786
rect 26910 32734 26962 32786
rect 29374 32734 29426 32786
rect 32062 32734 32114 32786
rect 37214 32734 37266 32786
rect 37550 32734 37602 32786
rect 46622 32734 46674 32786
rect 3950 32622 4002 32674
rect 4958 32622 5010 32674
rect 14814 32622 14866 32674
rect 25678 32622 25730 32674
rect 26014 32622 26066 32674
rect 27806 32622 27858 32674
rect 30382 32622 30434 32674
rect 36430 32622 36482 32674
rect 37998 32622 38050 32674
rect 40350 32622 40402 32674
rect 51662 32622 51714 32674
rect 52670 32622 52722 32674
rect 2718 32510 2770 32562
rect 3278 32510 3330 32562
rect 4286 32510 4338 32562
rect 5406 32510 5458 32562
rect 7422 32510 7474 32562
rect 8430 32510 8482 32562
rect 8766 32510 8818 32562
rect 8990 32510 9042 32562
rect 9998 32510 10050 32562
rect 10894 32510 10946 32562
rect 11902 32510 11954 32562
rect 12798 32510 12850 32562
rect 13582 32510 13634 32562
rect 14030 32510 14082 32562
rect 14254 32510 14306 32562
rect 16270 32510 16322 32562
rect 16942 32510 16994 32562
rect 18958 32510 19010 32562
rect 19518 32510 19570 32562
rect 22878 32510 22930 32562
rect 27134 32510 27186 32562
rect 28478 32510 28530 32562
rect 33518 32510 33570 32562
rect 34190 32510 34242 32562
rect 47518 32510 47570 32562
rect 48078 32510 48130 32562
rect 51998 32510 52050 32562
rect 3390 32398 3442 32450
rect 8542 32398 8594 32450
rect 12574 32398 12626 32450
rect 16606 32398 16658 32450
rect 19630 32398 19682 32450
rect 23102 32398 23154 32450
rect 23550 32398 23602 32450
rect 28926 32398 28978 32450
rect 38670 32398 38722 32450
rect 39118 32398 39170 32450
rect 41470 32398 41522 32450
rect 46174 32398 46226 32450
rect 48190 32398 48242 32450
rect 51102 32398 51154 32450
rect 53230 32398 53282 32450
rect 53678 32398 53730 32450
rect 55022 32398 55074 32450
rect 55918 32398 55970 32450
rect 56366 32398 56418 32450
rect 56814 32398 56866 32450
rect 57374 32398 57426 32450
rect 5182 32286 5234 32338
rect 5630 32286 5682 32338
rect 9886 32286 9938 32338
rect 10222 32286 10274 32338
rect 10334 32286 10386 32338
rect 52558 32286 52610 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 11118 31950 11170 32002
rect 19518 31950 19570 32002
rect 23326 31950 23378 32002
rect 7758 31838 7810 31890
rect 14590 31838 14642 31890
rect 14926 31838 14978 31890
rect 15710 31838 15762 31890
rect 16158 31838 16210 31890
rect 17054 31838 17106 31890
rect 20302 31838 20354 31890
rect 21982 31838 22034 31890
rect 22430 31838 22482 31890
rect 27358 31838 27410 31890
rect 29486 31838 29538 31890
rect 31390 31838 31442 31890
rect 39454 31838 39506 31890
rect 45726 31838 45778 31890
rect 53902 31838 53954 31890
rect 56926 31838 56978 31890
rect 57262 31838 57314 31890
rect 2830 31726 2882 31778
rect 4734 31726 4786 31778
rect 5966 31726 6018 31778
rect 6862 31726 6914 31778
rect 10110 31726 10162 31778
rect 10782 31726 10834 31778
rect 11902 31726 11954 31778
rect 12462 31726 12514 31778
rect 19854 31726 19906 31778
rect 23662 31726 23714 31778
rect 33854 31726 33906 31778
rect 34190 31726 34242 31778
rect 36766 31726 36818 31778
rect 40126 31726 40178 31778
rect 40462 31726 40514 31778
rect 46062 31726 46114 31778
rect 47630 31726 47682 31778
rect 48190 31726 48242 31778
rect 51550 31726 51602 31778
rect 52446 31726 52498 31778
rect 54686 31726 54738 31778
rect 55358 31726 55410 31778
rect 1822 31614 1874 31666
rect 2158 31614 2210 31666
rect 3054 31614 3106 31666
rect 3614 31614 3666 31666
rect 3950 31614 4002 31666
rect 4958 31614 5010 31666
rect 8430 31614 8482 31666
rect 8766 31614 8818 31666
rect 9550 31614 9602 31666
rect 9998 31614 10050 31666
rect 10558 31614 10610 31666
rect 11678 31614 11730 31666
rect 14142 31614 14194 31666
rect 22542 31614 22594 31666
rect 22766 31614 22818 31666
rect 28590 31614 28642 31666
rect 33966 31614 34018 31666
rect 36430 31614 36482 31666
rect 38446 31614 38498 31666
rect 46510 31614 46562 31666
rect 5742 31502 5794 31554
rect 6638 31502 6690 31554
rect 9774 31502 9826 31554
rect 13022 31502 13074 31554
rect 13582 31502 13634 31554
rect 19630 31502 19682 31554
rect 23438 31502 23490 31554
rect 24110 31502 24162 31554
rect 26574 31502 26626 31554
rect 43038 31502 43090 31554
rect 43598 31502 43650 31554
rect 47294 31502 47346 31554
rect 47518 31502 47570 31554
rect 48526 31502 48578 31554
rect 49086 31502 49138 31554
rect 50206 31502 50258 31554
rect 50766 31502 50818 31554
rect 51214 31502 51266 31554
rect 52110 31502 52162 31554
rect 53342 31502 53394 31554
rect 54462 31502 54514 31554
rect 55694 31502 55746 31554
rect 56254 31502 56306 31554
rect 57710 31502 57762 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 2046 31166 2098 31218
rect 3166 31166 3218 31218
rect 3614 31166 3666 31218
rect 4734 31166 4786 31218
rect 6414 31166 6466 31218
rect 7310 31166 7362 31218
rect 8094 31166 8146 31218
rect 8542 31166 8594 31218
rect 9998 31166 10050 31218
rect 11454 31166 11506 31218
rect 14142 31166 14194 31218
rect 14590 31166 14642 31218
rect 15486 31166 15538 31218
rect 17614 31166 17666 31218
rect 22654 31166 22706 31218
rect 22766 31166 22818 31218
rect 23774 31166 23826 31218
rect 27134 31166 27186 31218
rect 31278 31166 31330 31218
rect 40350 31166 40402 31218
rect 45838 31166 45890 31218
rect 47854 31166 47906 31218
rect 48638 31166 48690 31218
rect 50654 31166 50706 31218
rect 13358 31054 13410 31106
rect 15262 31054 15314 31106
rect 30494 31054 30546 31106
rect 32062 31054 32114 31106
rect 36206 31054 36258 31106
rect 42926 31054 42978 31106
rect 44270 31054 44322 31106
rect 48190 31054 48242 31106
rect 49534 31054 49586 31106
rect 51326 31054 51378 31106
rect 51662 31054 51714 31106
rect 54910 31054 54962 31106
rect 5070 30942 5122 30994
rect 6750 30942 6802 30994
rect 7646 30942 7698 30994
rect 9102 30942 9154 30994
rect 10334 30942 10386 30994
rect 15038 30942 15090 30994
rect 18398 30942 18450 30994
rect 18846 30942 18898 30994
rect 21086 30942 21138 30994
rect 27582 30942 27634 30994
rect 28142 30942 28194 30994
rect 37438 30942 37490 30994
rect 37774 30942 37826 30994
rect 44046 30942 44098 30994
rect 45390 30942 45442 30994
rect 45726 30942 45778 30994
rect 45950 30942 46002 30994
rect 46510 30942 46562 30994
rect 49870 30942 49922 30994
rect 50430 30942 50482 30994
rect 53118 30942 53170 30994
rect 55246 30942 55298 30994
rect 2382 30830 2434 30882
rect 4174 30830 4226 30882
rect 5518 30830 5570 30882
rect 10894 30830 10946 30882
rect 11118 30830 11170 30882
rect 12014 30830 12066 30882
rect 15150 30830 15202 30882
rect 16046 30830 16098 30882
rect 23438 30830 23490 30882
rect 24334 30830 24386 30882
rect 31614 30830 31666 30882
rect 32622 30830 32674 30882
rect 35422 30830 35474 30882
rect 35870 30830 35922 30882
rect 41582 30830 41634 30882
rect 44718 30830 44770 30882
rect 46846 30830 46898 30882
rect 47294 30830 47346 30882
rect 52670 30830 52722 30882
rect 53790 30830 53842 30882
rect 54350 30830 54402 30882
rect 55694 30830 55746 30882
rect 56142 30830 56194 30882
rect 56702 30830 56754 30882
rect 57486 30830 57538 30882
rect 57822 30830 57874 30882
rect 3614 30718 3666 30770
rect 4174 30718 4226 30770
rect 21982 30718 22034 30770
rect 22878 30718 22930 30770
rect 23214 30718 23266 30770
rect 23438 30718 23490 30770
rect 35422 30718 35474 30770
rect 36094 30718 36146 30770
rect 40910 30718 40962 30770
rect 50766 30718 50818 30770
rect 52334 30718 52386 30770
rect 53902 30718 53954 30770
rect 54686 30718 54738 30770
rect 55806 30718 55858 30770
rect 56142 30718 56194 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 3726 30382 3778 30434
rect 3950 30382 4002 30434
rect 14702 30382 14754 30434
rect 19182 30382 19234 30434
rect 22878 30382 22930 30434
rect 23214 30382 23266 30434
rect 33182 30382 33234 30434
rect 34078 30382 34130 30434
rect 38110 30382 38162 30434
rect 3726 30270 3778 30322
rect 19742 30270 19794 30322
rect 21982 30270 22034 30322
rect 33742 30270 33794 30322
rect 36430 30270 36482 30322
rect 36654 30270 36706 30322
rect 43262 30270 43314 30322
rect 50654 30270 50706 30322
rect 1934 30158 1986 30210
rect 5742 30158 5794 30210
rect 7310 30158 7362 30210
rect 7982 30158 8034 30210
rect 11902 30158 11954 30210
rect 14926 30158 14978 30210
rect 15598 30158 15650 30210
rect 15710 30158 15762 30210
rect 16270 30158 16322 30210
rect 16942 30158 16994 30210
rect 17950 30158 18002 30210
rect 18958 30158 19010 30210
rect 19630 30158 19682 30210
rect 20190 30158 20242 30210
rect 20526 30158 20578 30210
rect 23326 30158 23378 30210
rect 23886 30158 23938 30210
rect 27022 30158 27074 30210
rect 30270 30158 30322 30210
rect 31950 30158 32002 30210
rect 41134 30158 41186 30210
rect 43934 30158 43986 30210
rect 44494 30158 44546 30210
rect 46062 30158 46114 30210
rect 50878 30158 50930 30210
rect 52558 30158 52610 30210
rect 53790 30158 53842 30210
rect 57038 30158 57090 30210
rect 2382 30046 2434 30098
rect 2718 30046 2770 30098
rect 6414 30046 6466 30098
rect 8206 30046 8258 30098
rect 8766 30046 8818 30098
rect 9102 30046 9154 30098
rect 10222 30046 10274 30098
rect 10558 30046 10610 30098
rect 11454 30046 11506 30098
rect 12910 30046 12962 30098
rect 17166 30046 17218 30098
rect 17726 30046 17778 30098
rect 19406 30046 19458 30098
rect 20414 30046 20466 30098
rect 29598 30046 29650 30098
rect 29710 30046 29762 30098
rect 32286 30046 32338 30098
rect 32846 30046 32898 30098
rect 35086 30046 35138 30098
rect 35422 30046 35474 30098
rect 35870 30046 35922 30098
rect 36094 30046 36146 30098
rect 40238 30046 40290 30098
rect 41694 30046 41746 30098
rect 42478 30046 42530 30098
rect 44158 30046 44210 30098
rect 46510 30046 46562 30098
rect 46734 30046 46786 30098
rect 48526 30046 48578 30098
rect 49310 30046 49362 30098
rect 49646 30046 49698 30098
rect 50206 30046 50258 30098
rect 50430 30046 50482 30098
rect 55582 30046 55634 30098
rect 56478 30046 56530 30098
rect 3278 29934 3330 29986
rect 4286 29934 4338 29986
rect 4622 29934 4674 29986
rect 9662 29934 9714 29986
rect 11118 29934 11170 29986
rect 12350 29934 12402 29986
rect 13694 29934 13746 29986
rect 14366 29934 14418 29986
rect 21534 29934 21586 29986
rect 22430 29934 22482 29986
rect 22878 29934 22930 29986
rect 26238 29934 26290 29986
rect 27358 29934 27410 29986
rect 29934 29934 29986 29986
rect 30830 29934 30882 29986
rect 31278 29934 31330 29986
rect 32174 29934 32226 29986
rect 33070 29934 33122 29986
rect 33966 29934 34018 29986
rect 34526 29934 34578 29986
rect 35198 29934 35250 29986
rect 36766 29934 36818 29986
rect 37438 29934 37490 29986
rect 42030 29934 42082 29986
rect 44270 29934 44322 29986
rect 45390 29934 45442 29986
rect 46286 29934 46338 29986
rect 47294 29934 47346 29986
rect 47630 29934 47682 29986
rect 48190 29934 48242 29986
rect 51326 29934 51378 29986
rect 51662 29934 51714 29986
rect 52222 29934 52274 29986
rect 53454 29934 53506 29986
rect 54574 29934 54626 29986
rect 54910 29934 54962 29986
rect 55470 29934 55522 29986
rect 56142 29934 56194 29986
rect 57374 29934 57426 29986
rect 57822 29934 57874 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 2830 29598 2882 29650
rect 3278 29598 3330 29650
rect 4734 29598 4786 29650
rect 6078 29598 6130 29650
rect 6638 29598 6690 29650
rect 7198 29598 7250 29650
rect 7646 29598 7698 29650
rect 8318 29598 8370 29650
rect 8654 29598 8706 29650
rect 16942 29598 16994 29650
rect 18286 29598 18338 29650
rect 21534 29598 21586 29650
rect 22318 29598 22370 29650
rect 22654 29598 22706 29650
rect 28478 29598 28530 29650
rect 29262 29598 29314 29650
rect 30046 29598 30098 29650
rect 30718 29598 30770 29650
rect 35310 29598 35362 29650
rect 37662 29598 37714 29650
rect 41918 29598 41970 29650
rect 42366 29598 42418 29650
rect 43262 29598 43314 29650
rect 43710 29598 43762 29650
rect 44382 29598 44434 29650
rect 44606 29598 44658 29650
rect 47406 29598 47458 29650
rect 49646 29598 49698 29650
rect 54238 29598 54290 29650
rect 56702 29598 56754 29650
rect 4286 29486 4338 29538
rect 5182 29486 5234 29538
rect 9662 29486 9714 29538
rect 15374 29486 15426 29538
rect 23550 29486 23602 29538
rect 32510 29486 32562 29538
rect 35534 29486 35586 29538
rect 36542 29486 36594 29538
rect 38334 29486 38386 29538
rect 38670 29486 38722 29538
rect 39118 29486 39170 29538
rect 41582 29486 41634 29538
rect 42926 29486 42978 29538
rect 44830 29486 44882 29538
rect 45950 29486 46002 29538
rect 50318 29486 50370 29538
rect 51214 29486 51266 29538
rect 54350 29486 54402 29538
rect 57486 29486 57538 29538
rect 57822 29486 57874 29538
rect 10446 29374 10498 29426
rect 11454 29374 11506 29426
rect 14254 29374 14306 29426
rect 14702 29374 14754 29426
rect 14814 29374 14866 29426
rect 15598 29374 15650 29426
rect 18622 29374 18674 29426
rect 19294 29374 19346 29426
rect 23326 29374 23378 29426
rect 25566 29374 25618 29426
rect 26126 29374 26178 29426
rect 31838 29374 31890 29426
rect 33518 29374 33570 29426
rect 34862 29374 34914 29426
rect 35086 29374 35138 29426
rect 36430 29374 36482 29426
rect 36766 29374 36818 29426
rect 37102 29374 37154 29426
rect 37550 29374 37602 29426
rect 37774 29374 37826 29426
rect 46062 29374 46114 29426
rect 46622 29374 46674 29426
rect 47742 29374 47794 29426
rect 49758 29374 49810 29426
rect 50654 29374 50706 29426
rect 51438 29374 51490 29426
rect 51774 29374 51826 29426
rect 53566 29374 53618 29426
rect 54910 29374 54962 29426
rect 1934 29262 1986 29314
rect 2270 29262 2322 29314
rect 3726 29262 3778 29314
rect 5742 29262 5794 29314
rect 10894 29262 10946 29314
rect 11678 29262 11730 29314
rect 13358 29262 13410 29314
rect 16270 29262 16322 29314
rect 17614 29262 17666 29314
rect 23998 29262 24050 29314
rect 24894 29262 24946 29314
rect 30606 29262 30658 29314
rect 32062 29262 32114 29314
rect 34078 29262 34130 29314
rect 45950 29262 46002 29314
rect 48190 29262 48242 29314
rect 48862 29262 48914 29314
rect 51326 29262 51378 29314
rect 52110 29262 52162 29314
rect 52558 29262 52610 29314
rect 53006 29262 53058 29314
rect 56030 29262 56082 29314
rect 2270 29150 2322 29202
rect 3054 29150 3106 29202
rect 3390 29150 3442 29202
rect 4958 29150 5010 29202
rect 5406 29150 5458 29202
rect 5742 29150 5794 29202
rect 30494 29150 30546 29202
rect 35422 29150 35474 29202
rect 44718 29150 44770 29202
rect 49646 29150 49698 29202
rect 52558 29150 52610 29202
rect 53902 29150 53954 29202
rect 54238 29150 54290 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 3502 28814 3554 28866
rect 4062 28814 4114 28866
rect 35646 28814 35698 28866
rect 35982 28814 36034 28866
rect 36542 28814 36594 28866
rect 42478 28814 42530 28866
rect 48750 28814 48802 28866
rect 2606 28702 2658 28754
rect 3054 28702 3106 28754
rect 3614 28702 3666 28754
rect 4062 28702 4114 28754
rect 19966 28702 20018 28754
rect 22430 28702 22482 28754
rect 25902 28702 25954 28754
rect 26462 28702 26514 28754
rect 28814 28702 28866 28754
rect 29822 28702 29874 28754
rect 30606 28702 30658 28754
rect 32062 28702 32114 28754
rect 35758 28702 35810 28754
rect 36094 28702 36146 28754
rect 36542 28702 36594 28754
rect 40350 28702 40402 28754
rect 46174 28702 46226 28754
rect 46622 28702 46674 28754
rect 48414 28702 48466 28754
rect 49870 28702 49922 28754
rect 50430 28702 50482 28754
rect 52558 28702 52610 28754
rect 4510 28590 4562 28642
rect 4958 28590 5010 28642
rect 14030 28590 14082 28642
rect 14478 28590 14530 28642
rect 16606 28590 16658 28642
rect 30942 28590 30994 28642
rect 31726 28590 31778 28642
rect 32734 28590 32786 28642
rect 34638 28590 34690 28642
rect 35198 28590 35250 28642
rect 37774 28590 37826 28642
rect 38222 28590 38274 28642
rect 40798 28590 40850 28642
rect 41470 28590 41522 28642
rect 42590 28590 42642 28642
rect 42814 28590 42866 28642
rect 49310 28590 49362 28642
rect 50878 28590 50930 28642
rect 52110 28590 52162 28642
rect 53678 28590 53730 28642
rect 54574 28590 54626 28642
rect 55358 28590 55410 28642
rect 56590 28590 56642 28642
rect 57598 28590 57650 28642
rect 58046 28590 58098 28642
rect 25118 28478 25170 28530
rect 25454 28478 25506 28530
rect 27022 28478 27074 28530
rect 27358 28478 27410 28530
rect 30270 28478 30322 28530
rect 32286 28478 32338 28530
rect 33406 28478 33458 28530
rect 35086 28478 35138 28530
rect 41358 28478 41410 28530
rect 43486 28478 43538 28530
rect 44718 28478 44770 28530
rect 45614 28478 45666 28530
rect 45726 28478 45778 28530
rect 48526 28478 48578 28530
rect 51662 28478 51714 28530
rect 53454 28478 53506 28530
rect 54014 28478 54066 28530
rect 56366 28478 56418 28530
rect 57262 28478 57314 28530
rect 2158 28366 2210 28418
rect 17614 28366 17666 28418
rect 18062 28366 18114 28418
rect 32062 28366 32114 28418
rect 33742 28366 33794 28418
rect 34974 28366 35026 28418
rect 37438 28366 37490 28418
rect 37662 28366 37714 28418
rect 41134 28366 41186 28418
rect 42478 28366 42530 28418
rect 43822 28366 43874 28418
rect 44382 28366 44434 28418
rect 45390 28366 45442 28418
rect 47182 28366 47234 28418
rect 47630 28366 47682 28418
rect 51326 28366 51378 28418
rect 53566 28366 53618 28418
rect 55694 28366 55746 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 3502 28030 3554 28082
rect 4062 28030 4114 28082
rect 10334 28030 10386 28082
rect 15486 28030 15538 28082
rect 16942 28030 16994 28082
rect 23998 28030 24050 28082
rect 25678 28030 25730 28082
rect 26686 28030 26738 28082
rect 29710 28030 29762 28082
rect 32510 28030 32562 28082
rect 33630 28030 33682 28082
rect 37550 28030 37602 28082
rect 44046 28030 44098 28082
rect 47854 28030 47906 28082
rect 49646 28030 49698 28082
rect 50206 28030 50258 28082
rect 51774 28030 51826 28082
rect 53902 28030 53954 28082
rect 54686 28030 54738 28082
rect 14590 27918 14642 27970
rect 19182 27918 19234 27970
rect 28142 27918 28194 27970
rect 28478 27918 28530 27970
rect 29374 27918 29426 27970
rect 31278 27918 31330 27970
rect 35758 27918 35810 27970
rect 38446 27918 38498 27970
rect 39678 27918 39730 27970
rect 40686 27918 40738 27970
rect 40798 27918 40850 27970
rect 41582 27918 41634 27970
rect 42478 27918 42530 27970
rect 46958 27918 47010 27970
rect 47966 27918 48018 27970
rect 48190 27918 48242 27970
rect 49758 27918 49810 27970
rect 53006 27918 53058 27970
rect 55470 27918 55522 27970
rect 56366 27918 56418 27970
rect 57374 27918 57426 27970
rect 3054 27806 3106 27858
rect 11342 27806 11394 27858
rect 13470 27806 13522 27858
rect 14030 27806 14082 27858
rect 14926 27806 14978 27858
rect 17726 27806 17778 27858
rect 17950 27806 18002 27858
rect 18286 27806 18338 27858
rect 18846 27806 18898 27858
rect 21310 27806 21362 27858
rect 21646 27806 21698 27858
rect 26238 27806 26290 27858
rect 33966 27806 34018 27858
rect 35086 27806 35138 27858
rect 35982 27806 36034 27858
rect 38110 27806 38162 27858
rect 40014 27806 40066 27858
rect 40462 27806 40514 27858
rect 41918 27806 41970 27858
rect 42702 27806 42754 27858
rect 43262 27806 43314 27858
rect 43822 27806 43874 27858
rect 44494 27806 44546 27858
rect 45614 27806 45666 27858
rect 46398 27806 46450 27858
rect 46846 27806 46898 27858
rect 47630 27806 47682 27858
rect 49422 27806 49474 27858
rect 51662 27806 51714 27858
rect 51886 27806 51938 27858
rect 53230 27806 53282 27858
rect 55694 27806 55746 27858
rect 56702 27806 56754 27858
rect 1934 27694 1986 27746
rect 15822 27694 15874 27746
rect 16270 27694 16322 27746
rect 30270 27694 30322 27746
rect 36542 27694 36594 27746
rect 36990 27694 37042 27746
rect 39006 27694 39058 27746
rect 42590 27694 42642 27746
rect 43934 27694 43986 27746
rect 45726 27694 45778 27746
rect 48638 27694 48690 27746
rect 52334 27694 52386 27746
rect 54238 27694 54290 27746
rect 57822 27694 57874 27746
rect 24782 27582 24834 27634
rect 26014 27582 26066 27634
rect 34638 27582 34690 27634
rect 34750 27582 34802 27634
rect 34974 27582 35026 27634
rect 43038 27582 43090 27634
rect 45502 27582 45554 27634
rect 46958 27582 47010 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 43710 27246 43762 27298
rect 44046 27246 44098 27298
rect 56254 27246 56306 27298
rect 56590 27246 56642 27298
rect 2158 27134 2210 27186
rect 15150 27134 15202 27186
rect 18510 27134 18562 27186
rect 26126 27134 26178 27186
rect 28142 27134 28194 27186
rect 28590 27134 28642 27186
rect 30046 27134 30098 27186
rect 30382 27134 30434 27186
rect 30942 27134 30994 27186
rect 31390 27134 31442 27186
rect 32734 27134 32786 27186
rect 39678 27134 39730 27186
rect 43150 27134 43202 27186
rect 43598 27134 43650 27186
rect 44158 27134 44210 27186
rect 48190 27134 48242 27186
rect 56814 27134 56866 27186
rect 11006 27022 11058 27074
rect 25678 27022 25730 27074
rect 26686 27022 26738 27074
rect 27470 27022 27522 27074
rect 28030 27022 28082 27074
rect 34078 27022 34130 27074
rect 34862 27022 34914 27074
rect 35758 27022 35810 27074
rect 37662 27022 37714 27074
rect 37998 27022 38050 27074
rect 38222 27022 38274 27074
rect 38894 27022 38946 27074
rect 41582 27022 41634 27074
rect 41918 27022 41970 27074
rect 46062 27022 46114 27074
rect 47070 27022 47122 27074
rect 49086 27022 49138 27074
rect 49310 27022 49362 27074
rect 50206 27022 50258 27074
rect 51662 27022 51714 27074
rect 52670 27022 52722 27074
rect 53566 27022 53618 27074
rect 54350 27022 54402 27074
rect 57710 27022 57762 27074
rect 13022 26910 13074 26962
rect 13806 26910 13858 26962
rect 17166 26910 17218 26962
rect 21982 26910 22034 26962
rect 24558 26910 24610 26962
rect 27246 26910 27298 26962
rect 33966 26910 34018 26962
rect 34638 26910 34690 26962
rect 36878 26910 36930 26962
rect 37774 26910 37826 26962
rect 38670 26910 38722 26962
rect 39230 26910 39282 26962
rect 41358 26910 41410 26962
rect 42366 26910 42418 26962
rect 42702 26910 42754 26962
rect 44494 26910 44546 26962
rect 45614 26910 45666 26962
rect 47742 26910 47794 26962
rect 49198 26910 49250 26962
rect 50430 26910 50482 26962
rect 55582 26910 55634 26962
rect 11342 26798 11394 26850
rect 21646 26798 21698 26850
rect 24894 26798 24946 26850
rect 25342 26798 25394 26850
rect 25566 26798 25618 26850
rect 32174 26798 32226 26850
rect 34302 26798 34354 26850
rect 36318 26798 36370 26850
rect 39006 26798 39058 26850
rect 40126 26798 40178 26850
rect 40798 26798 40850 26850
rect 41582 26798 41634 26850
rect 42590 26798 42642 26850
rect 45838 26798 45890 26850
rect 45950 26798 46002 26850
rect 46846 26798 46898 26850
rect 50206 26798 50258 26850
rect 51326 26798 51378 26850
rect 52334 26798 52386 26850
rect 53790 26798 53842 26850
rect 54686 26798 54738 26850
rect 55246 26798 55298 26850
rect 57374 26798 57426 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 16270 26462 16322 26514
rect 24446 26462 24498 26514
rect 25006 26462 25058 26514
rect 25678 26462 25730 26514
rect 26350 26462 26402 26514
rect 27694 26462 27746 26514
rect 31502 26462 31554 26514
rect 33518 26462 33570 26514
rect 34750 26462 34802 26514
rect 35422 26462 35474 26514
rect 37102 26462 37154 26514
rect 37662 26462 37714 26514
rect 38446 26462 38498 26514
rect 38894 26462 38946 26514
rect 41582 26462 41634 26514
rect 43374 26462 43426 26514
rect 46622 26462 46674 26514
rect 47518 26462 47570 26514
rect 48526 26462 48578 26514
rect 18062 26350 18114 26402
rect 32062 26350 32114 26402
rect 35982 26350 36034 26402
rect 37998 26350 38050 26402
rect 39790 26350 39842 26402
rect 43934 26350 43986 26402
rect 48750 26350 48802 26402
rect 54910 26350 54962 26402
rect 56030 26350 56082 26402
rect 57374 26350 57426 26402
rect 13582 26238 13634 26290
rect 14030 26238 14082 26290
rect 18398 26238 18450 26290
rect 18958 26238 19010 26290
rect 19630 26238 19682 26290
rect 19854 26238 19906 26290
rect 20414 26238 20466 26290
rect 21310 26238 21362 26290
rect 21870 26238 21922 26290
rect 29934 26238 29986 26290
rect 30606 26238 30658 26290
rect 31614 26238 31666 26290
rect 32510 26238 32562 26290
rect 34526 26238 34578 26290
rect 35534 26238 35586 26290
rect 36542 26238 36594 26290
rect 36878 26238 36930 26290
rect 39342 26238 39394 26290
rect 44270 26238 44322 26290
rect 44830 26238 44882 26290
rect 45838 26238 45890 26290
rect 46174 26238 46226 26290
rect 47070 26238 47122 26290
rect 48302 26238 48354 26290
rect 50766 26238 50818 26290
rect 52670 26238 52722 26290
rect 53454 26238 53506 26290
rect 53678 26238 53730 26290
rect 56254 26238 56306 26290
rect 20862 26126 20914 26178
rect 40350 26126 40402 26178
rect 40686 26126 40738 26178
rect 42142 26126 42194 26178
rect 42590 26126 42642 26178
rect 49422 26126 49474 26178
rect 49870 26126 49922 26178
rect 50990 26126 51042 26178
rect 51550 26126 51602 26178
rect 53118 26126 53170 26178
rect 54462 26126 54514 26178
rect 55358 26126 55410 26178
rect 57822 26126 57874 26178
rect 17054 26014 17106 26066
rect 26126 26014 26178 26066
rect 26910 26014 26962 26066
rect 35422 26014 35474 26066
rect 37214 26014 37266 26066
rect 44270 26014 44322 26066
rect 48862 26014 48914 26066
rect 50430 26014 50482 26066
rect 51774 26014 51826 26066
rect 52110 26014 52162 26066
rect 57934 26014 57986 26066
rect 58270 26014 58322 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 20974 25678 21026 25730
rect 28142 25678 28194 25730
rect 35646 25678 35698 25730
rect 35870 25678 35922 25730
rect 37550 25678 37602 25730
rect 38110 25678 38162 25730
rect 38334 25678 38386 25730
rect 48862 25678 48914 25730
rect 49646 25678 49698 25730
rect 50878 25678 50930 25730
rect 51438 25678 51490 25730
rect 57598 25678 57650 25730
rect 16046 25566 16098 25618
rect 26014 25566 26066 25618
rect 27022 25566 27074 25618
rect 31502 25566 31554 25618
rect 41806 25566 41858 25618
rect 43150 25566 43202 25618
rect 47406 25566 47458 25618
rect 49534 25566 49586 25618
rect 51326 25566 51378 25618
rect 51774 25566 51826 25618
rect 52334 25566 52386 25618
rect 52670 25566 52722 25618
rect 56366 25566 56418 25618
rect 14590 25454 14642 25506
rect 15598 25454 15650 25506
rect 17502 25454 17554 25506
rect 17950 25454 18002 25506
rect 27582 25454 27634 25506
rect 27806 25454 27858 25506
rect 28030 25454 28082 25506
rect 31166 25454 31218 25506
rect 33966 25454 34018 25506
rect 35422 25454 35474 25506
rect 37662 25454 37714 25506
rect 38894 25454 38946 25506
rect 39118 25454 39170 25506
rect 39342 25454 39394 25506
rect 40574 25454 40626 25506
rect 43822 25454 43874 25506
rect 44158 25454 44210 25506
rect 47742 25454 47794 25506
rect 53790 25454 53842 25506
rect 55134 25454 55186 25506
rect 56478 25454 56530 25506
rect 57934 25454 57986 25506
rect 14366 25342 14418 25394
rect 15262 25342 15314 25394
rect 24670 25342 24722 25394
rect 31838 25342 31890 25394
rect 32398 25342 32450 25394
rect 32622 25342 32674 25394
rect 32734 25342 32786 25394
rect 32846 25342 32898 25394
rect 33742 25342 33794 25394
rect 34302 25342 34354 25394
rect 36430 25342 36482 25394
rect 36766 25342 36818 25394
rect 37886 25342 37938 25394
rect 39566 25342 39618 25394
rect 40238 25342 40290 25394
rect 41134 25342 41186 25394
rect 43038 25342 43090 25394
rect 43262 25342 43314 25394
rect 44494 25342 44546 25394
rect 46174 25342 46226 25394
rect 46846 25342 46898 25394
rect 47630 25342 47682 25394
rect 47966 25342 48018 25394
rect 50430 25342 50482 25394
rect 50878 25342 50930 25394
rect 54238 25342 54290 25394
rect 56030 25342 56082 25394
rect 20414 25230 20466 25282
rect 21534 25230 21586 25282
rect 24110 25230 24162 25282
rect 26462 25230 26514 25282
rect 28590 25230 28642 25282
rect 30046 25230 30098 25282
rect 32510 25230 32562 25282
rect 33966 25230 34018 25282
rect 34974 25230 35026 25282
rect 35086 25230 35138 25282
rect 35198 25230 35250 25282
rect 41246 25230 41298 25282
rect 41470 25230 41522 25282
rect 42254 25230 42306 25282
rect 44046 25230 44098 25282
rect 45838 25230 45890 25282
rect 46734 25230 46786 25282
rect 48190 25230 48242 25282
rect 48638 25230 48690 25282
rect 49086 25230 49138 25282
rect 50094 25230 50146 25282
rect 53454 25230 53506 25282
rect 54798 25230 54850 25282
rect 57710 25230 57762 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 14366 24894 14418 24946
rect 21422 24894 21474 24946
rect 21870 24894 21922 24946
rect 25902 24894 25954 24946
rect 27582 24894 27634 24946
rect 29710 24894 29762 24946
rect 30270 24894 30322 24946
rect 31390 24894 31442 24946
rect 32734 24894 32786 24946
rect 34302 24894 34354 24946
rect 37774 24894 37826 24946
rect 38222 24894 38274 24946
rect 40574 24894 40626 24946
rect 43822 24894 43874 24946
rect 46846 24894 46898 24946
rect 48078 24894 48130 24946
rect 51774 24894 51826 24946
rect 52334 24894 52386 24946
rect 52782 24894 52834 24946
rect 57486 24894 57538 24946
rect 14702 24782 14754 24834
rect 15262 24782 15314 24834
rect 18846 24782 18898 24834
rect 22878 24782 22930 24834
rect 24670 24782 24722 24834
rect 26910 24782 26962 24834
rect 27022 24782 27074 24834
rect 29822 24782 29874 24834
rect 36766 24782 36818 24834
rect 37326 24782 37378 24834
rect 38670 24782 38722 24834
rect 40126 24782 40178 24834
rect 46062 24782 46114 24834
rect 46958 24782 47010 24834
rect 47182 24782 47234 24834
rect 49982 24782 50034 24834
rect 51102 24782 51154 24834
rect 53902 24782 53954 24834
rect 54798 24782 54850 24834
rect 55134 24782 55186 24834
rect 56030 24782 56082 24834
rect 25678 24670 25730 24722
rect 26350 24670 26402 24722
rect 26686 24670 26738 24722
rect 27918 24670 27970 24722
rect 31950 24670 32002 24722
rect 33630 24670 33682 24722
rect 33966 24670 34018 24722
rect 34078 24670 34130 24722
rect 35198 24670 35250 24722
rect 35646 24670 35698 24722
rect 35870 24670 35922 24722
rect 39454 24670 39506 24722
rect 39678 24670 39730 24722
rect 39902 24670 39954 24722
rect 42254 24670 42306 24722
rect 42926 24670 42978 24722
rect 43934 24670 43986 24722
rect 44158 24670 44210 24722
rect 44382 24670 44434 24722
rect 45502 24670 45554 24722
rect 45726 24670 45778 24722
rect 46734 24670 46786 24722
rect 49646 24670 49698 24722
rect 49758 24670 49810 24722
rect 50206 24670 50258 24722
rect 50878 24670 50930 24722
rect 51886 24670 51938 24722
rect 54126 24670 54178 24722
rect 56366 24670 56418 24722
rect 56590 24670 56642 24722
rect 58046 24670 58098 24722
rect 20638 24558 20690 24610
rect 25790 24558 25842 24610
rect 30830 24558 30882 24610
rect 34190 24558 34242 24610
rect 36654 24558 36706 24610
rect 39790 24558 39842 24610
rect 41470 24558 41522 24610
rect 42702 24558 42754 24610
rect 44046 24558 44098 24610
rect 45950 24558 46002 24610
rect 47630 24558 47682 24610
rect 48526 24558 48578 24610
rect 53230 24558 53282 24610
rect 56142 24558 56194 24610
rect 29710 24446 29762 24498
rect 31838 24446 31890 24498
rect 32398 24446 32450 24498
rect 32622 24446 32674 24498
rect 35422 24446 35474 24498
rect 35982 24446 36034 24498
rect 36542 24446 36594 24498
rect 37550 24446 37602 24498
rect 37998 24446 38050 24498
rect 42478 24446 42530 24498
rect 43038 24446 43090 24498
rect 45614 24446 45666 24498
rect 47518 24446 47570 24498
rect 49646 24446 49698 24498
rect 51774 24446 51826 24498
rect 52110 24446 52162 24498
rect 53006 24446 53058 24498
rect 53678 24446 53730 24498
rect 55806 24446 55858 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 38894 24110 38946 24162
rect 39902 24110 39954 24162
rect 57150 24110 57202 24162
rect 57598 24110 57650 24162
rect 22542 23998 22594 24050
rect 23102 23998 23154 24050
rect 24334 23998 24386 24050
rect 27918 23998 27970 24050
rect 30606 23998 30658 24050
rect 32174 23998 32226 24050
rect 32958 23998 33010 24050
rect 34190 23998 34242 24050
rect 34974 23998 35026 24050
rect 47630 23998 47682 24050
rect 50766 23998 50818 24050
rect 56702 23998 56754 24050
rect 17502 23886 17554 23938
rect 17838 23886 17890 23938
rect 21758 23886 21810 23938
rect 23214 23886 23266 23938
rect 29934 23886 29986 23938
rect 31726 23886 31778 23938
rect 32734 23886 32786 23938
rect 34078 23886 34130 23938
rect 35198 23886 35250 23938
rect 38446 23886 38498 23938
rect 38670 23886 38722 23938
rect 39118 23886 39170 23938
rect 39454 23886 39506 23938
rect 40238 23886 40290 23938
rect 40462 23886 40514 23938
rect 40910 23886 40962 23938
rect 41246 23886 41298 23938
rect 41918 23886 41970 23938
rect 42366 23886 42418 23938
rect 42702 23886 42754 23938
rect 43710 23886 43762 23938
rect 46622 23886 46674 23938
rect 46734 23886 46786 23938
rect 46958 23886 47010 23938
rect 48638 23886 48690 23938
rect 49870 23886 49922 23938
rect 50990 23886 51042 23938
rect 52110 23886 52162 23938
rect 52670 23886 52722 23938
rect 53454 23886 53506 23938
rect 53678 23886 53730 23938
rect 55022 23886 55074 23938
rect 56926 23886 56978 23938
rect 22990 23774 23042 23826
rect 23550 23774 23602 23826
rect 26126 23774 26178 23826
rect 27470 23774 27522 23826
rect 33182 23774 33234 23826
rect 35422 23774 35474 23826
rect 35982 23774 36034 23826
rect 36318 23774 36370 23826
rect 37550 23774 37602 23826
rect 37886 23774 37938 23826
rect 43822 23774 43874 23826
rect 43934 23774 43986 23826
rect 44046 23774 44098 23826
rect 46286 23774 46338 23826
rect 47182 23774 47234 23826
rect 48974 23774 49026 23826
rect 51886 23774 51938 23826
rect 54014 23774 54066 23826
rect 56030 23774 56082 23826
rect 20414 23662 20466 23714
rect 20974 23662 21026 23714
rect 21982 23662 22034 23714
rect 27134 23662 27186 23714
rect 28926 23662 28978 23714
rect 30046 23662 30098 23714
rect 30270 23662 30322 23714
rect 34862 23662 34914 23714
rect 34974 23662 35026 23714
rect 36766 23662 36818 23714
rect 38894 23662 38946 23714
rect 41134 23662 41186 23714
rect 42030 23662 42082 23714
rect 42142 23662 42194 23714
rect 43598 23662 43650 23714
rect 45390 23662 45442 23714
rect 46622 23662 46674 23714
rect 48190 23662 48242 23714
rect 48862 23662 48914 23714
rect 49534 23662 49586 23714
rect 50430 23662 50482 23714
rect 52446 23662 52498 23714
rect 53902 23662 53954 23714
rect 57934 23662 57986 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 17950 23326 18002 23378
rect 20302 23326 20354 23378
rect 23774 23326 23826 23378
rect 24670 23326 24722 23378
rect 30382 23326 30434 23378
rect 31054 23326 31106 23378
rect 33966 23326 34018 23378
rect 36542 23326 36594 23378
rect 37102 23326 37154 23378
rect 37438 23326 37490 23378
rect 38782 23326 38834 23378
rect 39566 23326 39618 23378
rect 41470 23326 41522 23378
rect 44718 23326 44770 23378
rect 45950 23326 46002 23378
rect 46846 23326 46898 23378
rect 47294 23326 47346 23378
rect 47742 23326 47794 23378
rect 48750 23326 48802 23378
rect 51886 23326 51938 23378
rect 52110 23326 52162 23378
rect 55022 23326 55074 23378
rect 55470 23326 55522 23378
rect 56142 23326 56194 23378
rect 57486 23326 57538 23378
rect 21310 23214 21362 23266
rect 24894 23214 24946 23266
rect 27358 23214 27410 23266
rect 29150 23214 29202 23266
rect 35870 23214 35922 23266
rect 42814 23214 42866 23266
rect 53790 23214 53842 23266
rect 19182 23102 19234 23154
rect 19406 23102 19458 23154
rect 20750 23102 20802 23154
rect 25678 23102 25730 23154
rect 26126 23102 26178 23154
rect 27246 23102 27298 23154
rect 27582 23102 27634 23154
rect 28478 23102 28530 23154
rect 29262 23102 29314 23154
rect 29934 23102 29986 23154
rect 30158 23102 30210 23154
rect 31390 23102 31442 23154
rect 34638 23102 34690 23154
rect 34974 23102 35026 23154
rect 35086 23102 35138 23154
rect 40126 23102 40178 23154
rect 40350 23102 40402 23154
rect 40574 23102 40626 23154
rect 40798 23102 40850 23154
rect 42478 23102 42530 23154
rect 49534 23102 49586 23154
rect 49758 23102 49810 23154
rect 50094 23102 50146 23154
rect 50990 23102 51042 23154
rect 51662 23102 51714 23154
rect 53342 23102 53394 23154
rect 54014 23102 54066 23154
rect 55246 23102 55298 23154
rect 56478 23102 56530 23154
rect 18510 22990 18562 23042
rect 24558 22990 24610 23042
rect 26462 22990 26514 23042
rect 30046 22990 30098 23042
rect 31838 22990 31890 23042
rect 32398 22990 32450 23042
rect 32846 22990 32898 23042
rect 33518 22990 33570 23042
rect 34750 22990 34802 23042
rect 35758 22990 35810 23042
rect 37886 22990 37938 23042
rect 38334 22990 38386 23042
rect 40462 22990 40514 23042
rect 41918 22990 41970 23042
rect 43262 22990 43314 23042
rect 43710 22990 43762 23042
rect 44158 22990 44210 23042
rect 45054 22990 45106 23042
rect 45502 22990 45554 23042
rect 46398 22990 46450 23042
rect 48190 22990 48242 23042
rect 49646 22990 49698 23042
rect 50542 22990 50594 23042
rect 51774 22990 51826 23042
rect 53454 22990 53506 23042
rect 55134 22990 55186 23042
rect 56702 22990 56754 23042
rect 57934 22990 57986 23042
rect 28142 22878 28194 22930
rect 36094 22878 36146 22930
rect 36318 22878 36370 22930
rect 36654 22878 36706 22930
rect 37886 22878 37938 22930
rect 38446 22878 38498 22930
rect 47630 22878 47682 22930
rect 48526 22878 48578 22930
rect 53342 22878 53394 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 26014 22542 26066 22594
rect 32398 22542 32450 22594
rect 33406 22542 33458 22594
rect 34974 22542 35026 22594
rect 36094 22542 36146 22594
rect 42142 22542 42194 22594
rect 43262 22542 43314 22594
rect 52558 22542 52610 22594
rect 19742 22430 19794 22482
rect 23774 22430 23826 22482
rect 24782 22430 24834 22482
rect 25118 22430 25170 22482
rect 26238 22430 26290 22482
rect 26798 22430 26850 22482
rect 27470 22430 27522 22482
rect 27582 22430 27634 22482
rect 32174 22430 32226 22482
rect 35198 22430 35250 22482
rect 35758 22430 35810 22482
rect 36094 22430 36146 22482
rect 36542 22430 36594 22482
rect 37998 22430 38050 22482
rect 40014 22430 40066 22482
rect 41806 22430 41858 22482
rect 42142 22430 42194 22482
rect 43598 22430 43650 22482
rect 50430 22430 50482 22482
rect 57038 22430 57090 22482
rect 2830 22318 2882 22370
rect 18958 22318 19010 22370
rect 27246 22318 27298 22370
rect 27694 22318 27746 22370
rect 27918 22318 27970 22370
rect 28926 22318 28978 22370
rect 29710 22318 29762 22370
rect 33742 22318 33794 22370
rect 37662 22318 37714 22370
rect 39902 22318 39954 22370
rect 40350 22318 40402 22370
rect 42590 22318 42642 22370
rect 44382 22318 44434 22370
rect 46286 22318 46338 22370
rect 47294 22318 47346 22370
rect 47406 22318 47458 22370
rect 47630 22318 47682 22370
rect 48414 22318 48466 22370
rect 48638 22318 48690 22370
rect 53902 22318 53954 22370
rect 54014 22318 54066 22370
rect 54238 22318 54290 22370
rect 56814 22318 56866 22370
rect 57934 22318 57986 22370
rect 1934 22206 1986 22258
rect 18734 22206 18786 22258
rect 22094 22206 22146 22258
rect 22430 22206 22482 22258
rect 23214 22206 23266 22258
rect 23326 22206 23378 22258
rect 28030 22206 28082 22258
rect 31390 22206 31442 22258
rect 31726 22206 31778 22258
rect 34078 22206 34130 22258
rect 34302 22206 34354 22258
rect 39230 22206 39282 22258
rect 40238 22206 40290 22258
rect 40910 22206 40962 22258
rect 41246 22206 41298 22258
rect 45390 22206 45442 22258
rect 48190 22206 48242 22258
rect 48862 22206 48914 22258
rect 49086 22206 49138 22258
rect 52558 22206 52610 22258
rect 52670 22206 52722 22258
rect 54798 22206 54850 22258
rect 57598 22206 57650 22258
rect 22990 22094 23042 22146
rect 25678 22094 25730 22146
rect 29934 22094 29986 22146
rect 30718 22094 30770 22146
rect 32734 22094 32786 22146
rect 33182 22094 33234 22146
rect 33854 22094 33906 22146
rect 34862 22094 34914 22146
rect 37326 22094 37378 22146
rect 37550 22094 37602 22146
rect 37998 22094 38050 22146
rect 38222 22094 38274 22146
rect 38670 22094 38722 22146
rect 38782 22094 38834 22146
rect 39006 22094 39058 22146
rect 41134 22094 41186 22146
rect 43038 22094 43090 22146
rect 44046 22094 44098 22146
rect 45950 22094 46002 22146
rect 46174 22094 46226 22146
rect 46846 22094 46898 22146
rect 48638 22094 48690 22146
rect 49534 22094 49586 22146
rect 49982 22094 50034 22146
rect 50878 22094 50930 22146
rect 51326 22094 51378 22146
rect 51774 22094 51826 22146
rect 53454 22094 53506 22146
rect 55134 22094 55186 22146
rect 55582 22094 55634 22146
rect 56478 22094 56530 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 23550 21758 23602 21810
rect 26126 21758 26178 21810
rect 30718 21758 30770 21810
rect 34078 21758 34130 21810
rect 34638 21758 34690 21810
rect 35982 21758 36034 21810
rect 37326 21758 37378 21810
rect 39454 21758 39506 21810
rect 40238 21758 40290 21810
rect 41694 21758 41746 21810
rect 42142 21758 42194 21810
rect 42702 21758 42754 21810
rect 48190 21758 48242 21810
rect 49646 21758 49698 21810
rect 52894 21758 52946 21810
rect 53678 21758 53730 21810
rect 23326 21646 23378 21698
rect 24782 21646 24834 21698
rect 29150 21646 29202 21698
rect 29486 21646 29538 21698
rect 30606 21646 30658 21698
rect 30942 21646 30994 21698
rect 31950 21646 32002 21698
rect 37102 21646 37154 21698
rect 39342 21646 39394 21698
rect 39566 21646 39618 21698
rect 43486 21646 43538 21698
rect 22430 21534 22482 21586
rect 22654 21534 22706 21586
rect 23998 21534 24050 21586
rect 31390 21534 31442 21586
rect 31726 21534 31778 21586
rect 32174 21534 32226 21586
rect 33742 21534 33794 21586
rect 35422 21534 35474 21586
rect 36990 21534 37042 21586
rect 37998 21534 38050 21586
rect 40462 21534 40514 21586
rect 40910 21534 40962 21586
rect 41918 21534 41970 21586
rect 43598 21590 43650 21642
rect 45166 21646 45218 21698
rect 45390 21646 45442 21698
rect 45950 21646 46002 21698
rect 50654 21646 50706 21698
rect 54798 21646 54850 21698
rect 55022 21646 55074 21698
rect 55918 21646 55970 21698
rect 57822 21646 57874 21698
rect 44046 21534 44098 21586
rect 45054 21534 45106 21586
rect 46286 21534 46338 21586
rect 46958 21534 47010 21586
rect 47966 21534 48018 21586
rect 48750 21534 48802 21586
rect 49534 21534 49586 21586
rect 49758 21534 49810 21586
rect 50094 21534 50146 21586
rect 50990 21534 51042 21586
rect 51886 21534 51938 21586
rect 54126 21534 54178 21586
rect 55470 21534 55522 21586
rect 56030 21534 56082 21586
rect 57934 21534 57986 21586
rect 58270 21534 58322 21586
rect 21758 21422 21810 21474
rect 23438 21422 23490 21474
rect 24334 21422 24386 21474
rect 28254 21422 28306 21474
rect 28702 21422 28754 21474
rect 30046 21422 30098 21474
rect 31950 21422 32002 21474
rect 32622 21422 32674 21474
rect 34078 21422 34130 21474
rect 36430 21422 36482 21474
rect 37774 21422 37826 21474
rect 38782 21422 38834 21474
rect 40350 21422 40402 21474
rect 41806 21422 41858 21474
rect 44494 21422 44546 21474
rect 46510 21422 46562 21474
rect 46734 21422 46786 21474
rect 51438 21422 51490 21474
rect 52334 21422 52386 21474
rect 53230 21422 53282 21474
rect 54910 21422 54962 21474
rect 55694 21422 55746 21474
rect 56590 21422 56642 21474
rect 57486 21422 57538 21474
rect 24334 21310 24386 21362
rect 24670 21310 24722 21362
rect 25118 21310 25170 21362
rect 33966 21310 34018 21362
rect 35534 21310 35586 21362
rect 35758 21310 35810 21362
rect 36766 21310 36818 21362
rect 38334 21310 38386 21362
rect 43486 21310 43538 21362
rect 48302 21310 48354 21362
rect 52334 21310 52386 21362
rect 52894 21310 52946 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 33294 20974 33346 21026
rect 33518 20974 33570 21026
rect 34862 20974 34914 21026
rect 39342 20974 39394 21026
rect 40238 20974 40290 21026
rect 49534 20974 49586 21026
rect 50542 20974 50594 21026
rect 51438 20974 51490 21026
rect 51998 20974 52050 21026
rect 52334 20974 52386 21026
rect 52782 20974 52834 21026
rect 21758 20862 21810 20914
rect 22206 20862 22258 20914
rect 31054 20862 31106 20914
rect 31278 20862 31330 20914
rect 32622 20862 32674 20914
rect 33182 20862 33234 20914
rect 33518 20862 33570 20914
rect 36766 20862 36818 20914
rect 38446 20862 38498 20914
rect 39454 20862 39506 20914
rect 40238 20862 40290 20914
rect 44718 20862 44770 20914
rect 45390 20862 45442 20914
rect 51438 20862 51490 20914
rect 52222 20862 52274 20914
rect 54686 20862 54738 20914
rect 22542 20750 22594 20802
rect 23774 20750 23826 20802
rect 25902 20750 25954 20802
rect 26686 20750 26738 20802
rect 28478 20750 28530 20802
rect 29934 20750 29986 20802
rect 30718 20750 30770 20802
rect 32174 20750 32226 20802
rect 34414 20750 34466 20802
rect 34750 20750 34802 20802
rect 34974 20750 35026 20802
rect 38110 20750 38162 20802
rect 38222 20750 38274 20802
rect 38670 20750 38722 20802
rect 38894 20750 38946 20802
rect 40910 20750 40962 20802
rect 41246 20750 41298 20802
rect 41470 20750 41522 20802
rect 42366 20750 42418 20802
rect 42590 20750 42642 20802
rect 43822 20750 43874 20802
rect 46286 20750 46338 20802
rect 46734 20750 46786 20802
rect 47070 20750 47122 20802
rect 47966 20750 48018 20802
rect 49422 20750 49474 20802
rect 50878 20750 50930 20802
rect 53454 20750 53506 20802
rect 53790 20750 53842 20802
rect 54014 20750 54066 20802
rect 54126 20750 54178 20802
rect 54238 20750 54290 20802
rect 55694 20750 55746 20802
rect 57262 20750 57314 20802
rect 2382 20638 2434 20690
rect 2718 20638 2770 20690
rect 24110 20638 24162 20690
rect 24670 20638 24722 20690
rect 25006 20638 25058 20690
rect 25566 20638 25618 20690
rect 27134 20638 27186 20690
rect 28030 20638 28082 20690
rect 28702 20638 28754 20690
rect 35982 20638 36034 20690
rect 36094 20638 36146 20690
rect 36206 20638 36258 20690
rect 43710 20638 43762 20690
rect 44046 20638 44098 20690
rect 46510 20638 46562 20690
rect 48638 20638 48690 20690
rect 48862 20638 48914 20690
rect 50094 20638 50146 20690
rect 50318 20638 50370 20690
rect 57710 20638 57762 20690
rect 3278 20526 3330 20578
rect 23438 20526 23490 20578
rect 23998 20526 24050 20578
rect 27246 20526 27298 20578
rect 27358 20526 27410 20578
rect 27470 20526 27522 20578
rect 27918 20526 27970 20578
rect 28254 20526 28306 20578
rect 30158 20526 30210 20578
rect 31838 20526 31890 20578
rect 34526 20526 34578 20578
rect 35534 20526 35586 20578
rect 37998 20526 38050 20578
rect 39790 20526 39842 20578
rect 41246 20526 41298 20578
rect 42478 20526 42530 20578
rect 42814 20526 42866 20578
rect 44158 20526 44210 20578
rect 44270 20526 44322 20578
rect 46734 20526 46786 20578
rect 47630 20526 47682 20578
rect 48750 20526 48802 20578
rect 49086 20526 49138 20578
rect 50878 20526 50930 20578
rect 51774 20526 51826 20578
rect 52670 20526 52722 20578
rect 55582 20526 55634 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 23102 20190 23154 20242
rect 24782 20190 24834 20242
rect 26462 20190 26514 20242
rect 29038 20190 29090 20242
rect 30606 20190 30658 20242
rect 31838 20190 31890 20242
rect 33966 20190 34018 20242
rect 37326 20190 37378 20242
rect 38222 20190 38274 20242
rect 42926 20190 42978 20242
rect 43934 20190 43986 20242
rect 44158 20190 44210 20242
rect 45502 20190 45554 20242
rect 52334 20190 52386 20242
rect 53342 20190 53394 20242
rect 56366 20190 56418 20242
rect 57486 20190 57538 20242
rect 24334 20078 24386 20130
rect 25566 20078 25618 20130
rect 28142 20078 28194 20130
rect 28366 20078 28418 20130
rect 29934 20078 29986 20130
rect 31054 20078 31106 20130
rect 34862 20078 34914 20130
rect 35422 20078 35474 20130
rect 35870 20078 35922 20130
rect 36878 20078 36930 20130
rect 36990 20078 37042 20130
rect 39006 20078 39058 20130
rect 39454 20078 39506 20130
rect 40350 20078 40402 20130
rect 40798 20078 40850 20130
rect 42030 20078 42082 20130
rect 45390 20078 45442 20130
rect 50766 20078 50818 20130
rect 50878 20078 50930 20130
rect 52110 20078 52162 20130
rect 26686 19966 26738 20018
rect 27134 19966 27186 20018
rect 28478 19966 28530 20018
rect 29374 19966 29426 20018
rect 30718 19966 30770 20018
rect 30830 19966 30882 20018
rect 34302 19966 34354 20018
rect 35086 19966 35138 20018
rect 37102 19966 37154 20018
rect 38222 19966 38274 20018
rect 38558 19966 38610 20018
rect 38782 19966 38834 20018
rect 42366 19966 42418 20018
rect 43150 19966 43202 20018
rect 44382 19966 44434 20018
rect 45502 19966 45554 20018
rect 48190 19966 48242 20018
rect 48638 19966 48690 20018
rect 50542 19966 50594 20018
rect 51214 19966 51266 20018
rect 51886 19966 51938 20018
rect 53006 19966 53058 20018
rect 53790 19966 53842 20018
rect 54798 19966 54850 20018
rect 55246 19966 55298 20018
rect 57710 19966 57762 20018
rect 22430 19854 22482 19906
rect 23550 19854 23602 19906
rect 26574 19854 26626 19906
rect 27694 19854 27746 19906
rect 32510 19854 32562 19906
rect 34974 19854 35026 19906
rect 36318 19854 36370 19906
rect 39902 19854 39954 19906
rect 41470 19854 41522 19906
rect 43822 19854 43874 19906
rect 49422 19854 49474 19906
rect 49870 19854 49922 19906
rect 51326 19854 51378 19906
rect 51998 19854 52050 19906
rect 55358 19854 55410 19906
rect 24222 19742 24274 19794
rect 31726 19742 31778 19794
rect 32062 19742 32114 19794
rect 55582 19742 55634 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 25902 19406 25954 19458
rect 30830 19406 30882 19458
rect 31166 19406 31218 19458
rect 31614 19406 31666 19458
rect 44270 19406 44322 19458
rect 46958 19406 47010 19458
rect 47630 19406 47682 19458
rect 51102 19406 51154 19458
rect 26126 19294 26178 19346
rect 26574 19294 26626 19346
rect 32398 19294 32450 19346
rect 32846 19294 32898 19346
rect 36206 19294 36258 19346
rect 36542 19294 36594 19346
rect 39566 19294 39618 19346
rect 42030 19294 42082 19346
rect 46286 19294 46338 19346
rect 46734 19294 46786 19346
rect 47182 19294 47234 19346
rect 47630 19294 47682 19346
rect 48078 19294 48130 19346
rect 48526 19294 48578 19346
rect 48974 19294 49026 19346
rect 49422 19294 49474 19346
rect 49870 19294 49922 19346
rect 53342 19294 53394 19346
rect 24110 19182 24162 19234
rect 24446 19182 24498 19234
rect 33630 19182 33682 19234
rect 34526 19182 34578 19234
rect 34862 19182 34914 19234
rect 35310 19182 35362 19234
rect 38334 19182 38386 19234
rect 43150 19182 43202 19234
rect 44382 19182 44434 19234
rect 50542 19182 50594 19234
rect 50990 19182 51042 19234
rect 51326 19182 51378 19234
rect 55470 19182 55522 19234
rect 56254 19182 56306 19234
rect 57150 19182 57202 19234
rect 21646 19070 21698 19122
rect 21870 19070 21922 19122
rect 22206 19070 22258 19122
rect 25006 19070 25058 19122
rect 30830 19070 30882 19122
rect 31390 19070 31442 19122
rect 33518 19070 33570 19122
rect 34750 19070 34802 19122
rect 35646 19070 35698 19122
rect 39118 19070 39170 19122
rect 40014 19070 40066 19122
rect 45950 19070 46002 19122
rect 51550 19070 51602 19122
rect 54350 19070 54402 19122
rect 55022 19070 55074 19122
rect 55246 19070 55298 19122
rect 58046 19070 58098 19122
rect 22094 18958 22146 19010
rect 22654 18958 22706 19010
rect 23550 18958 23602 19010
rect 25566 18958 25618 19010
rect 27246 18958 27298 19010
rect 28702 18958 28754 19010
rect 29598 18958 29650 19010
rect 31950 18958 32002 19010
rect 33294 18958 33346 19010
rect 34190 18958 34242 19010
rect 35534 18958 35586 19010
rect 37550 18958 37602 19010
rect 37998 18958 38050 19010
rect 38222 18958 38274 19010
rect 38782 18958 38834 19010
rect 39006 18958 39058 19010
rect 40798 18958 40850 19010
rect 41134 18958 41186 19010
rect 41582 18958 41634 19010
rect 42814 18958 42866 19010
rect 43598 18958 43650 19010
rect 44270 18958 44322 19010
rect 45390 18958 45442 19010
rect 51662 18958 51714 19010
rect 51998 18958 52050 19010
rect 52446 18958 52498 19010
rect 54014 18958 54066 19010
rect 55358 18958 55410 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 24222 18622 24274 18674
rect 24894 18622 24946 18674
rect 27582 18622 27634 18674
rect 28030 18622 28082 18674
rect 31390 18622 31442 18674
rect 33518 18622 33570 18674
rect 37886 18622 37938 18674
rect 39006 18622 39058 18674
rect 39342 18622 39394 18674
rect 40126 18622 40178 18674
rect 42814 18622 42866 18674
rect 43934 18622 43986 18674
rect 44158 18622 44210 18674
rect 47294 18622 47346 18674
rect 48190 18622 48242 18674
rect 48414 18622 48466 18674
rect 16942 18510 16994 18562
rect 23214 18510 23266 18562
rect 23550 18510 23602 18562
rect 24446 18510 24498 18562
rect 25790 18510 25842 18562
rect 25902 18510 25954 18562
rect 26462 18510 26514 18562
rect 27694 18510 27746 18562
rect 31614 18510 31666 18562
rect 35310 18510 35362 18562
rect 35982 18510 36034 18562
rect 36094 18510 36146 18562
rect 38782 18510 38834 18562
rect 40238 18510 40290 18562
rect 42366 18510 42418 18562
rect 44046 18510 44098 18562
rect 44382 18510 44434 18562
rect 46622 18510 46674 18562
rect 47630 18510 47682 18562
rect 48302 18510 48354 18562
rect 51662 18510 51714 18562
rect 53454 18510 53506 18562
rect 54350 18510 54402 18562
rect 56254 18510 56306 18562
rect 57486 18510 57538 18562
rect 57822 18510 57874 18562
rect 16494 18398 16546 18450
rect 18174 18398 18226 18450
rect 18958 18398 19010 18450
rect 19630 18398 19682 18450
rect 20190 18398 20242 18450
rect 21198 18398 21250 18450
rect 21646 18398 21698 18450
rect 22094 18398 22146 18450
rect 26798 18398 26850 18450
rect 27022 18398 27074 18450
rect 27806 18398 27858 18450
rect 29262 18398 29314 18450
rect 29822 18398 29874 18450
rect 30718 18398 30770 18450
rect 32062 18398 32114 18450
rect 34974 18398 35026 18450
rect 35758 18398 35810 18450
rect 36542 18398 36594 18450
rect 36990 18398 37042 18450
rect 39230 18398 39282 18450
rect 40798 18398 40850 18450
rect 41918 18398 41970 18450
rect 42030 18398 42082 18450
rect 43822 18398 43874 18450
rect 44942 18398 44994 18450
rect 46734 18398 46786 18450
rect 48862 18398 48914 18450
rect 49646 18398 49698 18450
rect 49982 18398 50034 18450
rect 50766 18398 50818 18450
rect 51326 18398 51378 18450
rect 52782 18398 52834 18450
rect 53678 18398 53730 18450
rect 53902 18398 53954 18450
rect 54462 18398 54514 18450
rect 55134 18398 55186 18450
rect 55694 18398 55746 18450
rect 56478 18398 56530 18450
rect 16718 18286 16770 18338
rect 22766 18286 22818 18338
rect 24110 18286 24162 18338
rect 26910 18286 26962 18338
rect 28814 18286 28866 18338
rect 30382 18286 30434 18338
rect 31502 18286 31554 18338
rect 32398 18286 32450 18338
rect 32846 18286 32898 18338
rect 33966 18286 34018 18338
rect 34750 18286 34802 18338
rect 37438 18286 37490 18338
rect 39118 18286 39170 18338
rect 42254 18286 42306 18338
rect 45726 18286 45778 18338
rect 56030 18286 56082 18338
rect 25790 18174 25842 18226
rect 29822 18174 29874 18226
rect 30718 18174 30770 18226
rect 32174 18174 32226 18226
rect 32846 18174 32898 18226
rect 40014 18174 40066 18226
rect 45838 18174 45890 18226
rect 46622 18174 46674 18226
rect 49758 18174 49810 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 16606 17838 16658 17890
rect 17502 17838 17554 17890
rect 20862 17838 20914 17890
rect 30606 17838 30658 17890
rect 30830 17838 30882 17890
rect 39006 17838 39058 17890
rect 39902 17838 39954 17890
rect 44382 17838 44434 17890
rect 50990 17838 51042 17890
rect 51326 17838 51378 17890
rect 15150 17726 15202 17778
rect 16270 17726 16322 17778
rect 19854 17726 19906 17778
rect 20526 17726 20578 17778
rect 26126 17726 26178 17778
rect 28030 17726 28082 17778
rect 48302 17726 48354 17778
rect 55918 17726 55970 17778
rect 57934 17726 57986 17778
rect 2830 17614 2882 17666
rect 14366 17614 14418 17666
rect 15262 17614 15314 17666
rect 16830 17614 16882 17666
rect 20302 17614 20354 17666
rect 22654 17614 22706 17666
rect 23214 17614 23266 17666
rect 23886 17614 23938 17666
rect 24110 17614 24162 17666
rect 24558 17614 24610 17666
rect 24894 17614 24946 17666
rect 27246 17614 27298 17666
rect 29822 17614 29874 17666
rect 32398 17614 32450 17666
rect 32622 17614 32674 17666
rect 33518 17614 33570 17666
rect 33854 17614 33906 17666
rect 34414 17614 34466 17666
rect 35086 17614 35138 17666
rect 35310 17614 35362 17666
rect 36206 17614 36258 17666
rect 36542 17614 36594 17666
rect 36878 17614 36930 17666
rect 38894 17614 38946 17666
rect 39230 17614 39282 17666
rect 40238 17614 40290 17666
rect 41246 17614 41298 17666
rect 42142 17614 42194 17666
rect 42702 17614 42754 17666
rect 44158 17614 44210 17666
rect 44718 17614 44770 17666
rect 46062 17614 46114 17666
rect 47406 17614 47458 17666
rect 49646 17614 49698 17666
rect 51214 17614 51266 17666
rect 52558 17614 52610 17666
rect 53454 17614 53506 17666
rect 54910 17614 54962 17666
rect 56814 17614 56866 17666
rect 57262 17614 57314 17666
rect 1934 17502 1986 17554
rect 16046 17502 16098 17554
rect 16270 17502 16322 17554
rect 17838 17502 17890 17554
rect 18398 17502 18450 17554
rect 18622 17502 18674 17554
rect 21646 17502 21698 17554
rect 25342 17502 25394 17554
rect 25566 17502 25618 17554
rect 28254 17502 28306 17554
rect 28478 17502 28530 17554
rect 28590 17502 28642 17554
rect 29486 17502 29538 17554
rect 29710 17502 29762 17554
rect 31166 17502 31218 17554
rect 31390 17502 31442 17554
rect 31950 17502 32002 17554
rect 33742 17502 33794 17554
rect 35198 17502 35250 17554
rect 37662 17502 37714 17554
rect 38558 17502 38610 17554
rect 41918 17502 41970 17554
rect 42590 17502 42642 17554
rect 43934 17502 43986 17554
rect 45726 17502 45778 17554
rect 49758 17502 49810 17554
rect 50878 17502 50930 17554
rect 56702 17502 56754 17554
rect 17614 17390 17666 17442
rect 18510 17390 18562 17442
rect 23998 17390 24050 17442
rect 25230 17390 25282 17442
rect 26686 17390 26738 17442
rect 26798 17390 26850 17442
rect 26910 17390 26962 17442
rect 28814 17390 28866 17442
rect 30494 17390 30546 17442
rect 32174 17390 32226 17442
rect 32286 17390 32338 17442
rect 33406 17390 33458 17442
rect 33630 17390 33682 17442
rect 35758 17390 35810 17442
rect 36318 17390 36370 17442
rect 37550 17390 37602 17442
rect 38670 17390 38722 17442
rect 40014 17390 40066 17442
rect 40686 17390 40738 17442
rect 44718 17390 44770 17442
rect 50318 17390 50370 17442
rect 52334 17390 52386 17442
rect 53790 17390 53842 17442
rect 54238 17390 54290 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 2382 17054 2434 17106
rect 3278 17054 3330 17106
rect 16718 17054 16770 17106
rect 22990 17054 23042 17106
rect 25790 17054 25842 17106
rect 25902 17054 25954 17106
rect 26462 17054 26514 17106
rect 27246 17054 27298 17106
rect 28478 17054 28530 17106
rect 28702 17054 28754 17106
rect 28926 17054 28978 17106
rect 29598 17054 29650 17106
rect 29934 17054 29986 17106
rect 30494 17054 30546 17106
rect 31278 17054 31330 17106
rect 31950 17054 32002 17106
rect 32958 17054 33010 17106
rect 34750 17054 34802 17106
rect 35198 17054 35250 17106
rect 36766 17054 36818 17106
rect 39342 17054 39394 17106
rect 40462 17054 40514 17106
rect 42254 17054 42306 17106
rect 43934 17054 43986 17106
rect 45166 17054 45218 17106
rect 45838 17054 45890 17106
rect 46846 17054 46898 17106
rect 48190 17054 48242 17106
rect 51774 17054 51826 17106
rect 51998 17054 52050 17106
rect 53006 17054 53058 17106
rect 57486 17054 57538 17106
rect 2718 16942 2770 16994
rect 15374 16942 15426 16994
rect 16942 16942 16994 16994
rect 24222 16942 24274 16994
rect 27470 16942 27522 16994
rect 27582 16942 27634 16994
rect 33966 16942 34018 16994
rect 34526 16942 34578 16994
rect 37438 16942 37490 16994
rect 37998 16942 38050 16994
rect 38110 16942 38162 16994
rect 38222 16942 38274 16994
rect 40686 16942 40738 16994
rect 40798 16942 40850 16994
rect 42926 16942 42978 16994
rect 44718 16942 44770 16994
rect 46174 16942 46226 16994
rect 50206 16942 50258 16994
rect 53454 16942 53506 16994
rect 54126 16942 54178 16994
rect 54238 16942 54290 16994
rect 55358 16942 55410 16994
rect 56702 16942 56754 16994
rect 15934 16830 15986 16882
rect 16382 16830 16434 16882
rect 19966 16830 20018 16882
rect 21310 16830 21362 16882
rect 21646 16830 21698 16882
rect 22990 16830 23042 16882
rect 24670 16830 24722 16882
rect 30830 16830 30882 16882
rect 31838 16830 31890 16882
rect 32062 16830 32114 16882
rect 32510 16830 32562 16882
rect 33630 16830 33682 16882
rect 34974 16830 35026 16882
rect 35198 16830 35250 16882
rect 36318 16830 36370 16882
rect 36542 16830 36594 16882
rect 39454 16830 39506 16882
rect 39902 16830 39954 16882
rect 41470 16830 41522 16882
rect 42030 16830 42082 16882
rect 43150 16830 43202 16882
rect 43934 16830 43986 16882
rect 44494 16830 44546 16882
rect 47406 16830 47458 16882
rect 49870 16830 49922 16882
rect 50878 16830 50930 16882
rect 52446 16830 52498 16882
rect 53230 16830 53282 16882
rect 53902 16830 53954 16882
rect 54686 16830 54738 16882
rect 55134 16830 55186 16882
rect 28814 16718 28866 16770
rect 36094 16718 36146 16770
rect 36654 16718 36706 16770
rect 48750 16718 48802 16770
rect 49758 16718 49810 16770
rect 50766 16718 50818 16770
rect 51886 16718 51938 16770
rect 53342 16718 53394 16770
rect 25678 16606 25730 16658
rect 33630 16606 33682 16658
rect 35870 16606 35922 16658
rect 38670 16606 38722 16658
rect 44158 16606 44210 16658
rect 54462 16606 54514 16658
rect 57822 16830 57874 16882
rect 55582 16606 55634 16658
rect 56030 16606 56082 16658
rect 56254 16606 56306 16658
rect 56478 16606 56530 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 14814 16270 14866 16322
rect 28702 16270 28754 16322
rect 28926 16270 28978 16322
rect 33518 16270 33570 16322
rect 34750 16270 34802 16322
rect 36430 16270 36482 16322
rect 36766 16270 36818 16322
rect 43262 16270 43314 16322
rect 44382 16270 44434 16322
rect 47182 16270 47234 16322
rect 48526 16270 48578 16322
rect 50542 16270 50594 16322
rect 16494 16158 16546 16210
rect 19182 16158 19234 16210
rect 19966 16158 20018 16210
rect 21534 16158 21586 16210
rect 23214 16158 23266 16210
rect 25566 16158 25618 16210
rect 26350 16158 26402 16210
rect 28926 16158 28978 16210
rect 29598 16158 29650 16210
rect 29934 16158 29986 16210
rect 33406 16158 33458 16210
rect 34190 16158 34242 16210
rect 34750 16158 34802 16210
rect 35646 16158 35698 16210
rect 41806 16158 41858 16210
rect 44158 16158 44210 16210
rect 45390 16158 45442 16210
rect 47854 16158 47906 16210
rect 51998 16158 52050 16210
rect 52446 16158 52498 16210
rect 53902 16158 53954 16210
rect 55694 16158 55746 16210
rect 55918 16158 55970 16210
rect 16046 16046 16098 16098
rect 16382 16046 16434 16098
rect 17166 16046 17218 16098
rect 24110 16046 24162 16098
rect 24894 16046 24946 16098
rect 31390 16046 31442 16098
rect 32510 16046 32562 16098
rect 38670 16046 38722 16098
rect 39678 16046 39730 16098
rect 40686 16046 40738 16098
rect 42926 16046 42978 16098
rect 43486 16046 43538 16098
rect 46398 16046 46450 16098
rect 47294 16046 47346 16098
rect 48414 16046 48466 16098
rect 49086 16046 49138 16098
rect 49870 16046 49922 16098
rect 50318 16046 50370 16098
rect 56814 16046 56866 16098
rect 14702 15934 14754 15986
rect 18958 15934 19010 15986
rect 24670 15934 24722 15986
rect 28030 15934 28082 15986
rect 28366 15934 28418 15986
rect 32846 15934 32898 15986
rect 33742 15934 33794 15986
rect 36654 15934 36706 15986
rect 37774 15934 37826 15986
rect 38110 15934 38162 15986
rect 40126 15934 40178 15986
rect 40798 15934 40850 15986
rect 41918 15934 41970 15986
rect 42142 15934 42194 15986
rect 42702 15934 42754 15986
rect 44158 15934 44210 15986
rect 46174 15934 46226 15986
rect 47182 15934 47234 15986
rect 48526 15934 48578 15986
rect 49758 15934 49810 15986
rect 50094 15934 50146 15986
rect 51102 15934 51154 15986
rect 55694 15934 55746 15986
rect 57374 15934 57426 15986
rect 57710 15934 57762 15986
rect 14814 15822 14866 15874
rect 17054 15822 17106 15874
rect 19518 15822 19570 15874
rect 20414 15822 20466 15874
rect 21982 15822 22034 15874
rect 23774 15822 23826 15874
rect 26686 15822 26738 15874
rect 27134 15822 27186 15874
rect 31838 15822 31890 15874
rect 31950 15822 32002 15874
rect 32062 15822 32114 15874
rect 32734 15822 32786 15874
rect 35198 15822 35250 15874
rect 39790 15822 39842 15874
rect 42814 15822 42866 15874
rect 51550 15822 51602 15874
rect 53342 15822 53394 15874
rect 54462 15822 54514 15874
rect 54798 15822 54850 15874
rect 56478 15822 56530 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 16046 15486 16098 15538
rect 16830 15486 16882 15538
rect 18398 15486 18450 15538
rect 27918 15486 27970 15538
rect 28254 15486 28306 15538
rect 29598 15486 29650 15538
rect 30046 15486 30098 15538
rect 37774 15486 37826 15538
rect 38222 15486 38274 15538
rect 40350 15486 40402 15538
rect 42366 15486 42418 15538
rect 43710 15486 43762 15538
rect 44270 15486 44322 15538
rect 45502 15486 45554 15538
rect 46958 15486 47010 15538
rect 49422 15486 49474 15538
rect 52894 15486 52946 15538
rect 55022 15486 55074 15538
rect 57822 15486 57874 15538
rect 14478 15374 14530 15426
rect 15934 15374 15986 15426
rect 20526 15374 20578 15426
rect 21422 15374 21474 15426
rect 26574 15374 26626 15426
rect 34862 15374 34914 15426
rect 37326 15374 37378 15426
rect 42814 15374 42866 15426
rect 44606 15374 44658 15426
rect 45726 15374 45778 15426
rect 48414 15374 48466 15426
rect 50990 15374 51042 15426
rect 51438 15374 51490 15426
rect 52670 15374 52722 15426
rect 54126 15374 54178 15426
rect 56702 15374 56754 15426
rect 14702 15262 14754 15314
rect 19182 15262 19234 15314
rect 22654 15262 22706 15314
rect 24558 15262 24610 15314
rect 25566 15262 25618 15314
rect 26238 15262 26290 15314
rect 29150 15262 29202 15314
rect 33630 15262 33682 15314
rect 33966 15262 34018 15314
rect 35086 15262 35138 15314
rect 35982 15262 36034 15314
rect 36430 15262 36482 15314
rect 39342 15262 39394 15314
rect 39566 15262 39618 15314
rect 40798 15262 40850 15314
rect 41470 15262 41522 15314
rect 46174 15262 46226 15314
rect 47182 15262 47234 15314
rect 47518 15262 47570 15314
rect 50206 15262 50258 15314
rect 50542 15262 50594 15314
rect 51774 15262 51826 15314
rect 52558 15262 52610 15314
rect 53230 15262 53282 15314
rect 53678 15262 53730 15314
rect 53902 15262 53954 15314
rect 54798 15262 54850 15314
rect 55806 15262 55858 15314
rect 56366 15262 56418 15314
rect 57486 15262 57538 15314
rect 20414 15150 20466 15202
rect 22542 15150 22594 15202
rect 24446 15150 24498 15202
rect 26462 15150 26514 15202
rect 27358 15150 27410 15202
rect 32286 15150 32338 15202
rect 32734 15150 32786 15202
rect 34974 15150 35026 15202
rect 35758 15150 35810 15202
rect 38894 15150 38946 15202
rect 41918 15150 41970 15202
rect 43262 15150 43314 15202
rect 47070 15150 47122 15202
rect 47966 15150 48018 15202
rect 55694 15150 55746 15202
rect 23774 15038 23826 15090
rect 28814 15038 28866 15090
rect 29150 15038 29202 15090
rect 38782 15038 38834 15090
rect 40238 15038 40290 15090
rect 41022 15038 41074 15090
rect 43150 15038 43202 15090
rect 44158 15038 44210 15090
rect 45390 15038 45442 15090
rect 54238 15038 54290 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 14926 14702 14978 14754
rect 16158 14702 16210 14754
rect 36206 14702 36258 14754
rect 52670 14702 52722 14754
rect 14254 14590 14306 14642
rect 17614 14590 17666 14642
rect 18846 14590 18898 14642
rect 20302 14590 20354 14642
rect 21870 14590 21922 14642
rect 22542 14590 22594 14642
rect 25678 14590 25730 14642
rect 28702 14590 28754 14642
rect 31390 14590 31442 14642
rect 33742 14590 33794 14642
rect 35310 14590 35362 14642
rect 36766 14590 36818 14642
rect 37438 14590 37490 14642
rect 37886 14590 37938 14642
rect 48414 14590 48466 14642
rect 48862 14590 48914 14642
rect 50206 14590 50258 14642
rect 53902 14590 53954 14642
rect 58046 14590 58098 14642
rect 14702 14478 14754 14530
rect 18958 14478 19010 14530
rect 19406 14478 19458 14530
rect 20638 14478 20690 14530
rect 21534 14478 21586 14530
rect 22654 14478 22706 14530
rect 24222 14478 24274 14530
rect 24782 14478 24834 14530
rect 25790 14478 25842 14530
rect 26798 14478 26850 14530
rect 27358 14478 27410 14530
rect 28478 14478 28530 14530
rect 29486 14478 29538 14530
rect 31950 14478 32002 14530
rect 35646 14478 35698 14530
rect 36318 14478 36370 14530
rect 39230 14478 39282 14530
rect 40238 14478 40290 14530
rect 40798 14478 40850 14530
rect 41694 14478 41746 14530
rect 41806 14478 41858 14530
rect 42590 14478 42642 14530
rect 42814 14478 42866 14530
rect 43150 14478 43202 14530
rect 45838 14478 45890 14530
rect 47742 14478 47794 14530
rect 50542 14478 50594 14530
rect 53454 14478 53506 14530
rect 54238 14478 54290 14530
rect 55022 14478 55074 14530
rect 57374 14478 57426 14530
rect 13806 14366 13858 14418
rect 15934 14366 15986 14418
rect 17054 14366 17106 14418
rect 20862 14366 20914 14418
rect 24110 14366 24162 14418
rect 27806 14366 27858 14418
rect 29822 14366 29874 14418
rect 31054 14366 31106 14418
rect 35422 14366 35474 14418
rect 39006 14366 39058 14418
rect 40686 14366 40738 14418
rect 44270 14366 44322 14418
rect 45502 14366 45554 14418
rect 47070 14366 47122 14418
rect 49310 14366 49362 14418
rect 51438 14366 51490 14418
rect 54126 14366 54178 14418
rect 55134 14366 55186 14418
rect 55582 14366 55634 14418
rect 56142 14366 56194 14418
rect 15262 14254 15314 14306
rect 16046 14254 16098 14306
rect 16606 14254 16658 14306
rect 17950 14254 18002 14306
rect 18734 14254 18786 14306
rect 23438 14254 23490 14306
rect 24334 14254 24386 14306
rect 25342 14254 25394 14306
rect 25566 14254 25618 14306
rect 26686 14254 26738 14306
rect 26910 14254 26962 14306
rect 29710 14254 29762 14306
rect 30270 14254 30322 14306
rect 33294 14254 33346 14306
rect 35870 14254 35922 14306
rect 38446 14254 38498 14306
rect 39454 14254 39506 14306
rect 39566 14254 39618 14306
rect 40462 14254 40514 14306
rect 41358 14254 41410 14306
rect 41470 14254 41522 14306
rect 41582 14254 41634 14306
rect 42814 14254 42866 14306
rect 44046 14254 44098 14306
rect 44382 14254 44434 14306
rect 44494 14254 44546 14306
rect 46734 14254 46786 14306
rect 47966 14254 48018 14306
rect 50318 14254 50370 14306
rect 51102 14254 51154 14306
rect 52446 14254 52498 14306
rect 52558 14254 52610 14306
rect 55358 14254 55410 14306
rect 56478 14254 56530 14306
rect 57038 14254 57090 14306
rect 57934 14254 57986 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 13918 13918 13970 13970
rect 15710 13918 15762 13970
rect 16494 13918 16546 13970
rect 18734 13918 18786 13970
rect 19742 13918 19794 13970
rect 20190 13918 20242 13970
rect 22990 13918 23042 13970
rect 24558 13918 24610 13970
rect 26014 13918 26066 13970
rect 26126 13918 26178 13970
rect 26238 13918 26290 13970
rect 31390 13918 31442 13970
rect 35198 13918 35250 13970
rect 37214 13918 37266 13970
rect 40574 13918 40626 13970
rect 42590 13918 42642 13970
rect 43934 13918 43986 13970
rect 44046 13918 44098 13970
rect 44830 13918 44882 13970
rect 45726 13918 45778 13970
rect 46846 13918 46898 13970
rect 48190 13918 48242 13970
rect 50542 13918 50594 13970
rect 51438 13918 51490 13970
rect 52446 13918 52498 13970
rect 55134 13918 55186 13970
rect 55806 13918 55858 13970
rect 56142 13918 56194 13970
rect 57374 13918 57426 13970
rect 15822 13806 15874 13858
rect 16718 13806 16770 13858
rect 22542 13806 22594 13858
rect 24894 13806 24946 13858
rect 28366 13806 28418 13858
rect 31278 13806 31330 13858
rect 36206 13806 36258 13858
rect 38110 13806 38162 13858
rect 39342 13806 39394 13858
rect 39566 13806 39618 13858
rect 39678 13806 39730 13858
rect 40350 13806 40402 13858
rect 41918 13806 41970 13858
rect 46734 13806 46786 13858
rect 49982 13806 50034 13858
rect 50878 13806 50930 13858
rect 53118 13806 53170 13858
rect 53454 13806 53506 13858
rect 54126 13806 54178 13858
rect 54462 13806 54514 13858
rect 55358 13806 55410 13858
rect 14478 13694 14530 13746
rect 14702 13694 14754 13746
rect 14926 13694 14978 13746
rect 15486 13694 15538 13746
rect 16046 13694 16098 13746
rect 16830 13694 16882 13746
rect 19070 13694 19122 13746
rect 21982 13694 22034 13746
rect 22318 13694 22370 13746
rect 25566 13694 25618 13746
rect 27806 13694 27858 13746
rect 28478 13694 28530 13746
rect 29262 13694 29314 13746
rect 30270 13694 30322 13746
rect 35758 13694 35810 13746
rect 36542 13694 36594 13746
rect 38334 13694 38386 13746
rect 38670 13694 38722 13746
rect 39902 13694 39954 13746
rect 40686 13694 40738 13746
rect 41806 13694 41858 13746
rect 42142 13694 42194 13746
rect 43374 13694 43426 13746
rect 43710 13694 43762 13746
rect 46510 13694 46562 13746
rect 47182 13694 47234 13746
rect 48414 13694 48466 13746
rect 49422 13694 49474 13746
rect 49758 13694 49810 13746
rect 51774 13694 51826 13746
rect 52222 13694 52274 13746
rect 52558 13694 52610 13746
rect 55022 13694 55074 13746
rect 19294 13582 19346 13634
rect 20862 13582 20914 13634
rect 23438 13582 23490 13634
rect 28926 13582 28978 13634
rect 29150 13582 29202 13634
rect 32398 13582 32450 13634
rect 39118 13582 39170 13634
rect 42926 13582 42978 13634
rect 44382 13582 44434 13634
rect 45278 13582 45330 13634
rect 48302 13582 48354 13634
rect 49982 13582 50034 13634
rect 56590 13582 56642 13634
rect 57822 13582 57874 13634
rect 14366 13470 14418 13522
rect 19518 13470 19570 13522
rect 20190 13470 20242 13522
rect 31502 13470 31554 13522
rect 37998 13470 38050 13522
rect 47070 13470 47122 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 15262 13134 15314 13186
rect 15934 13134 15986 13186
rect 16382 13134 16434 13186
rect 28254 13134 28306 13186
rect 29934 13134 29986 13186
rect 36094 13134 36146 13186
rect 15038 13022 15090 13074
rect 16494 13022 16546 13074
rect 20862 13022 20914 13074
rect 21534 13022 21586 13074
rect 28590 13022 28642 13074
rect 29598 13022 29650 13074
rect 30494 13022 30546 13074
rect 31614 13022 31666 13074
rect 34862 13022 34914 13074
rect 37550 13022 37602 13074
rect 38334 13022 38386 13074
rect 39230 13022 39282 13074
rect 39454 13022 39506 13074
rect 41246 13022 41298 13074
rect 41582 13022 41634 13074
rect 43486 13022 43538 13074
rect 45502 13022 45554 13074
rect 45950 13022 46002 13074
rect 52670 13022 52722 13074
rect 53790 13022 53842 13074
rect 54910 13022 54962 13074
rect 57262 13022 57314 13074
rect 15486 12910 15538 12962
rect 24670 12910 24722 12962
rect 25118 12910 25170 12962
rect 26014 12910 26066 12962
rect 31950 12910 32002 12962
rect 32958 12910 33010 12962
rect 33182 12910 33234 12962
rect 33966 12910 34018 12962
rect 35086 12910 35138 12962
rect 42702 12910 42754 12962
rect 42926 12910 42978 12962
rect 44158 12910 44210 12962
rect 44382 12910 44434 12962
rect 46510 12910 46562 12962
rect 46734 12910 46786 12962
rect 48638 12910 48690 12962
rect 50318 12910 50370 12962
rect 51886 12910 51938 12962
rect 54238 12910 54290 12962
rect 18958 12798 19010 12850
rect 19854 12798 19906 12850
rect 19966 12798 20018 12850
rect 25454 12798 25506 12850
rect 28814 12798 28866 12850
rect 31502 12798 31554 12850
rect 31838 12798 31890 12850
rect 32622 12798 32674 12850
rect 33854 12798 33906 12850
rect 34750 12798 34802 12850
rect 35310 12798 35362 12850
rect 35870 12798 35922 12850
rect 42366 12798 42418 12850
rect 48862 12798 48914 12850
rect 51438 12798 51490 12850
rect 53454 12798 53506 12850
rect 53790 12798 53842 12850
rect 56142 12798 56194 12850
rect 18510 12686 18562 12738
rect 19070 12686 19122 12738
rect 19294 12686 19346 12738
rect 19630 12686 19682 12738
rect 20526 12686 20578 12738
rect 26350 12686 26402 12738
rect 26462 12686 26514 12738
rect 26574 12686 26626 12738
rect 29710 12686 29762 12738
rect 30942 12686 30994 12738
rect 33630 12686 33682 12738
rect 36430 12686 36482 12738
rect 37886 12686 37938 12738
rect 39790 12686 39842 12738
rect 40350 12686 40402 12738
rect 40686 12686 40738 12738
rect 42814 12686 42866 12738
rect 44718 12686 44770 12738
rect 46622 12686 46674 12738
rect 46958 12686 47010 12738
rect 47518 12686 47570 12738
rect 49646 12686 49698 12738
rect 53678 12686 53730 12738
rect 56814 12686 56866 12738
rect 57710 12686 57762 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 2718 12350 2770 12402
rect 15150 12350 15202 12402
rect 15374 12350 15426 12402
rect 24894 12350 24946 12402
rect 29262 12350 29314 12402
rect 30382 12350 30434 12402
rect 31166 12350 31218 12402
rect 34750 12350 34802 12402
rect 35198 12350 35250 12402
rect 36654 12350 36706 12402
rect 39342 12350 39394 12402
rect 39678 12350 39730 12402
rect 40238 12350 40290 12402
rect 42030 12350 42082 12402
rect 42814 12350 42866 12402
rect 43710 12350 43762 12402
rect 44270 12350 44322 12402
rect 47182 12350 47234 12402
rect 48750 12350 48802 12402
rect 49534 12350 49586 12402
rect 51662 12350 51714 12402
rect 52222 12350 52274 12402
rect 53454 12350 53506 12402
rect 54126 12350 54178 12402
rect 54686 12350 54738 12402
rect 55134 12350 55186 12402
rect 56030 12350 56082 12402
rect 56590 12350 56642 12402
rect 57374 12350 57426 12402
rect 27246 12238 27298 12290
rect 28254 12238 28306 12290
rect 28590 12238 28642 12290
rect 32622 12238 32674 12290
rect 37102 12238 37154 12290
rect 40574 12238 40626 12290
rect 45502 12238 45554 12290
rect 46174 12238 46226 12290
rect 50990 12238 51042 12290
rect 54238 12238 54290 12290
rect 2494 12126 2546 12178
rect 15262 12126 15314 12178
rect 15710 12126 15762 12178
rect 18622 12126 18674 12178
rect 19518 12126 19570 12178
rect 20862 12126 20914 12178
rect 21198 12126 21250 12178
rect 21982 12126 22034 12178
rect 22654 12126 22706 12178
rect 25902 12126 25954 12178
rect 26350 12126 26402 12178
rect 27582 12126 27634 12178
rect 28702 12126 28754 12178
rect 31054 12126 31106 12178
rect 31278 12126 31330 12178
rect 31502 12126 31554 12178
rect 31838 12126 31890 12178
rect 32510 12126 32562 12178
rect 35534 12126 35586 12178
rect 35870 12126 35922 12178
rect 37214 12126 37266 12178
rect 37326 12126 37378 12178
rect 38782 12126 38834 12178
rect 42590 12126 42642 12178
rect 43262 12126 43314 12178
rect 44830 12126 44882 12178
rect 45726 12126 45778 12178
rect 46510 12126 46562 12178
rect 47406 12126 47458 12178
rect 47854 12126 47906 12178
rect 49870 12126 49922 12178
rect 50094 12126 50146 12178
rect 50766 12126 50818 12178
rect 51550 12126 51602 12178
rect 53230 12126 53282 12178
rect 53566 12126 53618 12178
rect 3166 12014 3218 12066
rect 19406 12014 19458 12066
rect 20302 12014 20354 12066
rect 22878 12014 22930 12066
rect 27358 12014 27410 12066
rect 28366 12014 28418 12066
rect 29934 12014 29986 12066
rect 30494 12014 30546 12066
rect 33518 12014 33570 12066
rect 33966 12014 34018 12066
rect 41470 12014 41522 12066
rect 42702 12014 42754 12066
rect 47294 12014 47346 12066
rect 48190 12014 48242 12066
rect 52670 12014 52722 12066
rect 55694 12014 55746 12066
rect 57822 12014 57874 12066
rect 26126 11902 26178 11954
rect 26798 11902 26850 11954
rect 32398 11902 32450 11954
rect 35310 11902 35362 11954
rect 36094 11902 36146 11954
rect 51662 11902 51714 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 22878 11566 22930 11618
rect 25678 11566 25730 11618
rect 28814 11566 28866 11618
rect 29038 11566 29090 11618
rect 31390 11566 31442 11618
rect 32510 11566 32562 11618
rect 39230 11566 39282 11618
rect 39790 11566 39842 11618
rect 42814 11566 42866 11618
rect 43150 11566 43202 11618
rect 44158 11566 44210 11618
rect 44382 11566 44434 11618
rect 44830 11566 44882 11618
rect 46958 11566 47010 11618
rect 47406 11566 47458 11618
rect 48190 11566 48242 11618
rect 54574 11566 54626 11618
rect 55470 11566 55522 11618
rect 55918 11566 55970 11618
rect 56366 11566 56418 11618
rect 56814 11566 56866 11618
rect 14254 11454 14306 11506
rect 18286 11454 18338 11506
rect 20526 11454 20578 11506
rect 21870 11454 21922 11506
rect 23214 11454 23266 11506
rect 28814 11454 28866 11506
rect 32062 11454 32114 11506
rect 34190 11454 34242 11506
rect 36206 11454 36258 11506
rect 36766 11454 36818 11506
rect 38782 11454 38834 11506
rect 39118 11454 39170 11506
rect 39790 11454 39842 11506
rect 40126 11454 40178 11506
rect 40574 11454 40626 11506
rect 41582 11454 41634 11506
rect 43262 11454 43314 11506
rect 48302 11454 48354 11506
rect 49198 11454 49250 11506
rect 51102 11454 51154 11506
rect 51662 11454 51714 11506
rect 55134 11454 55186 11506
rect 55582 11454 55634 11506
rect 55918 11454 55970 11506
rect 56814 11454 56866 11506
rect 57374 11454 57426 11506
rect 2830 11342 2882 11394
rect 14926 11342 14978 11394
rect 15150 11342 15202 11394
rect 15710 11342 15762 11394
rect 19742 11342 19794 11394
rect 19854 11342 19906 11394
rect 23102 11342 23154 11394
rect 23998 11342 24050 11394
rect 25006 11342 25058 11394
rect 25230 11342 25282 11394
rect 26350 11342 26402 11394
rect 27918 11342 27970 11394
rect 28254 11342 28306 11394
rect 29598 11342 29650 11394
rect 30606 11342 30658 11394
rect 31054 11342 31106 11394
rect 31950 11342 32002 11394
rect 32622 11342 32674 11394
rect 33630 11342 33682 11394
rect 42926 11342 42978 11394
rect 43934 11342 43986 11394
rect 45614 11342 45666 11394
rect 45950 11342 46002 11394
rect 46174 11342 46226 11394
rect 46398 11342 46450 11394
rect 46734 11342 46786 11394
rect 49982 11342 50034 11394
rect 50430 11342 50482 11394
rect 50654 11342 50706 11394
rect 53566 11342 53618 11394
rect 53678 11342 53730 11394
rect 53790 11342 53842 11394
rect 54014 11342 54066 11394
rect 1934 11230 1986 11282
rect 15934 11230 15986 11282
rect 16046 11230 16098 11282
rect 19630 11230 19682 11282
rect 27582 11230 27634 11282
rect 29934 11230 29986 11282
rect 32174 11230 32226 11282
rect 35870 11230 35922 11282
rect 35982 11230 36034 11282
rect 37550 11230 37602 11282
rect 37886 11230 37938 11282
rect 46846 11230 46898 11282
rect 48750 11230 48802 11282
rect 50318 11230 50370 11282
rect 52446 11230 52498 11282
rect 18174 11118 18226 11170
rect 19182 11118 19234 11170
rect 24110 11118 24162 11170
rect 24334 11118 24386 11170
rect 26686 11118 26738 11170
rect 28030 11118 28082 11170
rect 29822 11118 29874 11170
rect 31278 11118 31330 11170
rect 33182 11118 33234 11170
rect 36094 11118 36146 11170
rect 36318 11118 36370 11170
rect 41134 11118 41186 11170
rect 42030 11118 42082 11170
rect 45726 11118 45778 11170
rect 45838 11118 45890 11170
rect 47406 11118 47458 11170
rect 47854 11118 47906 11170
rect 49646 11118 49698 11170
rect 52558 11118 52610 11170
rect 53902 11118 53954 11170
rect 54574 11118 54626 11170
rect 56366 11118 56418 11170
rect 57710 11118 57762 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 2382 10782 2434 10834
rect 3278 10782 3330 10834
rect 14814 10782 14866 10834
rect 16606 10782 16658 10834
rect 17950 10782 18002 10834
rect 24894 10782 24946 10834
rect 28366 10782 28418 10834
rect 37102 10782 37154 10834
rect 37438 10782 37490 10834
rect 39342 10782 39394 10834
rect 41582 10782 41634 10834
rect 42478 10782 42530 10834
rect 42926 10782 42978 10834
rect 43262 10782 43314 10834
rect 43822 10782 43874 10834
rect 44494 10782 44546 10834
rect 45054 10782 45106 10834
rect 46062 10782 46114 10834
rect 47182 10782 47234 10834
rect 47742 10782 47794 10834
rect 48078 10782 48130 10834
rect 48638 10782 48690 10834
rect 49534 10782 49586 10834
rect 50318 10782 50370 10834
rect 51214 10782 51266 10834
rect 51774 10782 51826 10834
rect 53566 10782 53618 10834
rect 54126 10782 54178 10834
rect 54574 10782 54626 10834
rect 55134 10782 55186 10834
rect 55694 10782 55746 10834
rect 56478 10782 56530 10834
rect 57374 10782 57426 10834
rect 57822 10782 57874 10834
rect 2718 10670 2770 10722
rect 15934 10670 15986 10722
rect 16830 10670 16882 10722
rect 18062 10670 18114 10722
rect 19182 10670 19234 10722
rect 19518 10670 19570 10722
rect 23998 10670 24050 10722
rect 30494 10670 30546 10722
rect 32062 10670 32114 10722
rect 35758 10670 35810 10722
rect 36094 10670 36146 10722
rect 37662 10670 37714 10722
rect 38670 10670 38722 10722
rect 44942 10670 44994 10722
rect 50206 10670 50258 10722
rect 50542 10670 50594 10722
rect 51102 10670 51154 10722
rect 52782 10670 52834 10722
rect 52894 10670 52946 10722
rect 53342 10670 53394 10722
rect 53678 10670 53730 10722
rect 15598 10558 15650 10610
rect 16158 10558 16210 10610
rect 16942 10558 16994 10610
rect 17726 10558 17778 10610
rect 18286 10558 18338 10610
rect 19630 10558 19682 10610
rect 22542 10558 22594 10610
rect 24334 10558 24386 10610
rect 25902 10558 25954 10610
rect 26126 10558 26178 10610
rect 27582 10558 27634 10610
rect 29150 10558 29202 10610
rect 29374 10558 29426 10610
rect 31166 10558 31218 10610
rect 31390 10558 31442 10610
rect 32398 10558 32450 10610
rect 34302 10558 34354 10610
rect 34638 10558 34690 10610
rect 34750 10558 34802 10610
rect 37774 10558 37826 10610
rect 38446 10558 38498 10610
rect 39454 10558 39506 10610
rect 40014 10558 40066 10610
rect 40238 10558 40290 10610
rect 50094 10558 50146 10610
rect 15038 10446 15090 10498
rect 16046 10446 16098 10498
rect 19294 10446 19346 10498
rect 22878 10446 22930 10498
rect 25678 10446 25730 10498
rect 27806 10446 27858 10498
rect 28926 10446 28978 10498
rect 32846 10446 32898 10498
rect 33742 10446 33794 10498
rect 34414 10446 34466 10498
rect 36542 10446 36594 10498
rect 41918 10446 41970 10498
rect 45726 10446 45778 10498
rect 46734 10446 46786 10498
rect 56030 10446 56082 10498
rect 14702 10334 14754 10386
rect 22990 10334 23042 10386
rect 27246 10334 27298 10386
rect 36318 10334 36370 10386
rect 36878 10334 36930 10386
rect 39342 10334 39394 10386
rect 40574 10334 40626 10386
rect 45054 10334 45106 10386
rect 51214 10334 51266 10386
rect 52782 10334 52834 10386
rect 57374 10334 57426 10386
rect 57934 10334 57986 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 17502 9998 17554 10050
rect 17838 9998 17890 10050
rect 26350 9998 26402 10050
rect 32174 9998 32226 10050
rect 32398 9998 32450 10050
rect 32846 9998 32898 10050
rect 33182 9998 33234 10050
rect 33406 9998 33458 10050
rect 33966 9998 34018 10050
rect 44718 9998 44770 10050
rect 48078 9998 48130 10050
rect 48526 9998 48578 10050
rect 51550 9998 51602 10050
rect 14590 9886 14642 9938
rect 15598 9886 15650 9938
rect 16494 9886 16546 9938
rect 21534 9886 21586 9938
rect 23102 9886 23154 9938
rect 28814 9886 28866 9938
rect 34750 9886 34802 9938
rect 34862 9886 34914 9938
rect 35534 9886 35586 9938
rect 35758 9886 35810 9938
rect 37886 9886 37938 9938
rect 38334 9886 38386 9938
rect 41918 9886 41970 9938
rect 45390 9886 45442 9938
rect 46174 9886 46226 9938
rect 46510 9886 46562 9938
rect 48526 9886 48578 9938
rect 49086 9886 49138 9938
rect 49646 9886 49698 9938
rect 50318 9886 50370 9938
rect 52558 9886 52610 9938
rect 53790 9886 53842 9938
rect 54686 9886 54738 9938
rect 55246 9886 55298 9938
rect 55582 9886 55634 9938
rect 57038 9886 57090 9938
rect 57374 9886 57426 9938
rect 14702 9774 14754 9826
rect 16270 9774 16322 9826
rect 24110 9774 24162 9826
rect 25230 9774 25282 9826
rect 26014 9774 26066 9826
rect 29486 9774 29538 9826
rect 29822 9774 29874 9826
rect 30046 9774 30098 9826
rect 33854 9774 33906 9826
rect 36766 9774 36818 9826
rect 38558 9774 38610 9826
rect 40014 9774 40066 9826
rect 40686 9774 40738 9826
rect 41470 9774 41522 9826
rect 42142 9774 42194 9826
rect 42814 9774 42866 9826
rect 47518 9774 47570 9826
rect 50206 9774 50258 9826
rect 53342 9774 53394 9826
rect 58046 9774 58098 9826
rect 2382 9662 2434 9714
rect 2718 9662 2770 9714
rect 3278 9662 3330 9714
rect 13806 9662 13858 9714
rect 17614 9662 17666 9714
rect 22990 9662 23042 9714
rect 23214 9662 23266 9714
rect 25790 9662 25842 9714
rect 36094 9662 36146 9714
rect 36318 9662 36370 9714
rect 39902 9662 39954 9714
rect 40238 9662 40290 9714
rect 42478 9662 42530 9714
rect 42702 9662 42754 9714
rect 43822 9662 43874 9714
rect 51326 9662 51378 9714
rect 52110 9662 52162 9714
rect 54350 9662 54402 9714
rect 23774 9550 23826 9602
rect 24894 9550 24946 9602
rect 26238 9550 26290 9602
rect 26686 9550 26738 9602
rect 27134 9550 27186 9602
rect 29822 9550 29874 9602
rect 30606 9550 30658 9602
rect 32510 9550 32562 9602
rect 33070 9550 33122 9602
rect 35422 9550 35474 9602
rect 39342 9550 39394 9602
rect 43486 9550 43538 9602
rect 44494 9550 44546 9602
rect 44606 9550 44658 9602
rect 47294 9550 47346 9602
rect 48190 9550 48242 9602
rect 51438 9550 51490 9602
rect 56030 9550 56082 9602
rect 56478 9550 56530 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 21982 9214 22034 9266
rect 25006 9214 25058 9266
rect 25678 9214 25730 9266
rect 27470 9214 27522 9266
rect 29038 9214 29090 9266
rect 31614 9214 31666 9266
rect 32846 9214 32898 9266
rect 35982 9214 36034 9266
rect 36206 9214 36258 9266
rect 37214 9214 37266 9266
rect 38446 9214 38498 9266
rect 39230 9214 39282 9266
rect 40350 9214 40402 9266
rect 40910 9214 40962 9266
rect 41694 9214 41746 9266
rect 46062 9214 46114 9266
rect 46510 9214 46562 9266
rect 47294 9214 47346 9266
rect 48638 9214 48690 9266
rect 51886 9214 51938 9266
rect 55582 9214 55634 9266
rect 56030 9214 56082 9266
rect 56478 9214 56530 9266
rect 57374 9214 57426 9266
rect 58046 9214 58098 9266
rect 12686 9102 12738 9154
rect 13022 9102 13074 9154
rect 26686 9102 26738 9154
rect 26910 9102 26962 9154
rect 29822 9102 29874 9154
rect 31390 9102 31442 9154
rect 34974 9102 35026 9154
rect 35198 9102 35250 9154
rect 35534 9102 35586 9154
rect 39342 9102 39394 9154
rect 39678 9102 39730 9154
rect 42478 9102 42530 9154
rect 42926 9102 42978 9154
rect 43374 9102 43426 9154
rect 47742 9102 47794 9154
rect 19630 8990 19682 9042
rect 21086 8990 21138 9042
rect 25902 8990 25954 9042
rect 26126 8990 26178 9042
rect 30158 8990 30210 9042
rect 33742 8990 33794 9042
rect 33966 8990 34018 9042
rect 34190 8990 34242 9042
rect 34414 8990 34466 9042
rect 36318 8990 36370 9042
rect 38222 8990 38274 9042
rect 38334 8990 38386 9042
rect 38782 8990 38834 9042
rect 39454 8990 39506 9042
rect 42030 8990 42082 9042
rect 43598 8990 43650 9042
rect 44718 8990 44770 9042
rect 45054 8990 45106 9042
rect 47854 8990 47906 9042
rect 47966 8990 48018 9042
rect 50318 8990 50370 9042
rect 50766 8990 50818 9042
rect 51438 8990 51490 9042
rect 52894 8990 52946 9042
rect 54462 8990 54514 9042
rect 55022 8990 55074 9042
rect 20638 8878 20690 8930
rect 22542 8878 22594 8930
rect 22990 8878 23042 8930
rect 25790 8878 25842 8930
rect 26910 8878 26962 8930
rect 32174 8878 32226 8930
rect 35422 8878 35474 8930
rect 36766 8878 36818 8930
rect 45614 8878 45666 8930
rect 49870 8878 49922 8930
rect 52670 8878 52722 8930
rect 53566 8878 53618 8930
rect 55134 8878 55186 8930
rect 19518 8766 19570 8818
rect 33630 8766 33682 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 16494 8430 16546 8482
rect 21982 8430 22034 8482
rect 25678 8430 25730 8482
rect 25902 8430 25954 8482
rect 36542 8430 36594 8482
rect 42926 8430 42978 8482
rect 43598 8430 43650 8482
rect 17166 8318 17218 8370
rect 19630 8318 19682 8370
rect 20414 8318 20466 8370
rect 22766 8318 22818 8370
rect 23550 8318 23602 8370
rect 24446 8318 24498 8370
rect 25342 8318 25394 8370
rect 27022 8318 27074 8370
rect 30494 8318 30546 8370
rect 31166 8318 31218 8370
rect 33294 8318 33346 8370
rect 34638 8318 34690 8370
rect 36430 8318 36482 8370
rect 39230 8318 39282 8370
rect 42142 8318 42194 8370
rect 43150 8318 43202 8370
rect 48078 8318 48130 8370
rect 48526 8318 48578 8370
rect 48974 8318 49026 8370
rect 49534 8318 49586 8370
rect 49870 8318 49922 8370
rect 53790 8318 53842 8370
rect 56366 8318 56418 8370
rect 57486 8318 57538 8370
rect 58046 8318 58098 8370
rect 17278 8206 17330 8258
rect 18510 8206 18562 8258
rect 18622 8206 18674 8258
rect 20638 8206 20690 8258
rect 25006 8206 25058 8258
rect 25118 8206 25170 8258
rect 25566 8206 25618 8258
rect 25902 8206 25954 8258
rect 26574 8206 26626 8258
rect 26910 8206 26962 8258
rect 28030 8206 28082 8258
rect 30046 8206 30098 8258
rect 34190 8206 34242 8258
rect 34974 8206 35026 8258
rect 37550 8206 37602 8258
rect 39006 8206 39058 8258
rect 40910 8206 40962 8258
rect 41134 8206 41186 8258
rect 41358 8206 41410 8258
rect 42702 8206 42754 8258
rect 44046 8206 44098 8258
rect 45502 8206 45554 8258
rect 45838 8206 45890 8258
rect 47742 8206 47794 8258
rect 51998 8206 52050 8258
rect 52446 8206 52498 8258
rect 53678 8206 53730 8258
rect 54574 8206 54626 8258
rect 55134 8206 55186 8258
rect 18062 8094 18114 8146
rect 18286 8094 18338 8146
rect 22206 8094 22258 8146
rect 23774 8094 23826 8146
rect 27694 8094 27746 8146
rect 27806 8094 27858 8146
rect 29598 8094 29650 8146
rect 33070 8094 33122 8146
rect 34638 8094 34690 8146
rect 35086 8094 35138 8146
rect 38782 8094 38834 8146
rect 39342 8094 39394 8146
rect 41582 8094 41634 8146
rect 46734 8094 46786 8146
rect 50990 8094 51042 8146
rect 51662 8094 51714 8146
rect 52558 8094 52610 8146
rect 18846 7982 18898 8034
rect 20078 7982 20130 8034
rect 21646 7982 21698 8034
rect 23214 7982 23266 8034
rect 27134 7982 27186 8034
rect 28478 7982 28530 8034
rect 33182 7982 33234 8034
rect 35982 7982 36034 8034
rect 37886 7982 37938 8034
rect 39902 7982 39954 8034
rect 44382 7982 44434 8034
rect 45614 7982 45666 8034
rect 46958 7982 47010 8034
rect 47070 7982 47122 8034
rect 47182 7982 47234 8034
rect 47966 7982 48018 8034
rect 50318 7982 50370 8034
rect 51774 7982 51826 8034
rect 52782 7982 52834 8034
rect 55246 7982 55298 8034
rect 55470 7982 55522 8034
rect 55806 7982 55858 8034
rect 56926 7982 56978 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 20414 7646 20466 7698
rect 31614 7646 31666 7698
rect 36990 7646 37042 7698
rect 37886 7646 37938 7698
rect 38334 7646 38386 7698
rect 42478 7646 42530 7698
rect 42702 7646 42754 7698
rect 42814 7646 42866 7698
rect 43822 7646 43874 7698
rect 44382 7646 44434 7698
rect 45054 7646 45106 7698
rect 47518 7646 47570 7698
rect 48190 7646 48242 7698
rect 50654 7646 50706 7698
rect 51662 7646 51714 7698
rect 54350 7646 54402 7698
rect 56814 7646 56866 7698
rect 57598 7646 57650 7698
rect 58046 7646 58098 7698
rect 17726 7534 17778 7586
rect 18062 7534 18114 7586
rect 18286 7534 18338 7586
rect 20078 7534 20130 7586
rect 20302 7534 20354 7586
rect 24894 7534 24946 7586
rect 28478 7534 28530 7586
rect 29374 7534 29426 7586
rect 36206 7534 36258 7586
rect 36542 7534 36594 7586
rect 43486 7534 43538 7586
rect 45502 7534 45554 7586
rect 45726 7534 45778 7586
rect 48414 7534 48466 7586
rect 49646 7534 49698 7586
rect 49758 7534 49810 7586
rect 52782 7534 52834 7586
rect 20750 7422 20802 7474
rect 22094 7422 22146 7474
rect 23438 7422 23490 7474
rect 23886 7422 23938 7474
rect 24558 7422 24610 7474
rect 25678 7422 25730 7474
rect 26574 7422 26626 7474
rect 27022 7422 27074 7474
rect 28142 7422 28194 7474
rect 29038 7422 29090 7474
rect 31726 7422 31778 7474
rect 31950 7422 32002 7474
rect 32174 7422 32226 7474
rect 35198 7422 35250 7474
rect 35646 7422 35698 7474
rect 42926 7422 42978 7474
rect 46174 7422 46226 7474
rect 46622 7422 46674 7474
rect 46846 7422 46898 7474
rect 47854 7422 47906 7474
rect 53230 7422 53282 7474
rect 53566 7422 53618 7474
rect 56142 7422 56194 7474
rect 17838 7310 17890 7362
rect 21422 7310 21474 7362
rect 22318 7310 22370 7362
rect 22990 7310 23042 7362
rect 25790 7310 25842 7362
rect 27470 7310 27522 7362
rect 28254 7310 28306 7362
rect 29822 7310 29874 7362
rect 30942 7310 30994 7362
rect 31838 7310 31890 7362
rect 37438 7310 37490 7362
rect 45950 7310 46002 7362
rect 47070 7310 47122 7362
rect 50206 7310 50258 7362
rect 51102 7310 51154 7362
rect 51998 7310 52050 7362
rect 52782 7310 52834 7362
rect 55358 7310 55410 7362
rect 24558 7198 24610 7250
rect 29038 7198 29090 7250
rect 35086 7198 35138 7250
rect 35422 7198 35474 7250
rect 48526 7198 48578 7250
rect 49646 7198 49698 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19182 6862 19234 6914
rect 41918 6862 41970 6914
rect 51326 6862 51378 6914
rect 20974 6750 21026 6802
rect 21646 6750 21698 6802
rect 28702 6750 28754 6802
rect 33294 6750 33346 6802
rect 42702 6750 42754 6802
rect 49198 6750 49250 6802
rect 57822 6750 57874 6802
rect 19294 6638 19346 6690
rect 19630 6638 19682 6690
rect 22878 6638 22930 6690
rect 23214 6638 23266 6690
rect 23438 6638 23490 6690
rect 23998 6638 24050 6690
rect 24222 6638 24274 6690
rect 24670 6638 24722 6690
rect 27470 6638 27522 6690
rect 28030 6638 28082 6690
rect 30830 6638 30882 6690
rect 31390 6638 31442 6690
rect 31614 6638 31666 6690
rect 32174 6638 32226 6690
rect 32846 6638 32898 6690
rect 33070 6638 33122 6690
rect 34638 6638 34690 6690
rect 35310 6638 35362 6690
rect 35758 6638 35810 6690
rect 36542 6638 36594 6690
rect 38222 6638 38274 6690
rect 38782 6638 38834 6690
rect 43598 6638 43650 6690
rect 45390 6638 45442 6690
rect 46174 6638 46226 6690
rect 46622 6638 46674 6690
rect 47966 6638 48018 6690
rect 48190 6638 48242 6690
rect 49310 6638 49362 6690
rect 50654 6638 50706 6690
rect 52558 6638 52610 6690
rect 53454 6638 53506 6690
rect 53790 6638 53842 6690
rect 54238 6638 54290 6690
rect 54798 6638 54850 6690
rect 55918 6638 55970 6690
rect 56814 6638 56866 6690
rect 2718 6526 2770 6578
rect 27134 6526 27186 6578
rect 28142 6526 28194 6578
rect 30718 6526 30770 6578
rect 31726 6526 31778 6578
rect 36206 6526 36258 6578
rect 46062 6526 46114 6578
rect 48526 6526 48578 6578
rect 55358 6526 55410 6578
rect 56254 6526 56306 6578
rect 2382 6414 2434 6466
rect 3166 6414 3218 6466
rect 22990 6414 23042 6466
rect 24110 6414 24162 6466
rect 29486 6414 29538 6466
rect 30494 6414 30546 6466
rect 32398 6414 32450 6466
rect 32958 6414 33010 6466
rect 33854 6414 33906 6466
rect 35086 6414 35138 6466
rect 35198 6414 35250 6466
rect 37438 6414 37490 6466
rect 41134 6414 41186 6466
rect 43038 6414 43090 6466
rect 44046 6414 44098 6466
rect 44382 6414 44434 6466
rect 48078 6414 48130 6466
rect 51998 6414 52050 6466
rect 57150 6414 57202 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 20638 6078 20690 6130
rect 24558 6078 24610 6130
rect 27582 6078 27634 6130
rect 32510 6078 32562 6130
rect 42702 6078 42754 6130
rect 44494 6078 44546 6130
rect 45278 6078 45330 6130
rect 45390 6078 45442 6130
rect 45950 6078 46002 6130
rect 46510 6078 46562 6130
rect 47182 6078 47234 6130
rect 48078 6078 48130 6130
rect 48414 6078 48466 6130
rect 49758 6078 49810 6130
rect 51326 6078 51378 6130
rect 52446 6078 52498 6130
rect 53342 6078 53394 6130
rect 53790 6078 53842 6130
rect 54462 6078 54514 6130
rect 55918 6078 55970 6130
rect 56366 6078 56418 6130
rect 57934 6078 57986 6130
rect 20414 5966 20466 6018
rect 24334 5966 24386 6018
rect 27246 5966 27298 6018
rect 31166 5966 31218 6018
rect 32622 5966 32674 6018
rect 33630 5966 33682 6018
rect 40126 5966 40178 6018
rect 40910 5966 40962 6018
rect 42814 5966 42866 6018
rect 43486 5966 43538 6018
rect 43822 5966 43874 6018
rect 44382 5966 44434 6018
rect 45502 5966 45554 6018
rect 49870 5966 49922 6018
rect 53006 5966 53058 6018
rect 54910 5966 54962 6018
rect 2830 5854 2882 5906
rect 22094 5854 22146 5906
rect 28366 5854 28418 5906
rect 33966 5854 34018 5906
rect 35758 5854 35810 5906
rect 36206 5854 36258 5906
rect 37214 5854 37266 5906
rect 37886 5854 37938 5906
rect 49534 5854 49586 5906
rect 57374 5854 57426 5906
rect 1934 5742 1986 5794
rect 28142 5742 28194 5794
rect 30718 5742 30770 5794
rect 34190 5742 34242 5794
rect 34638 5742 34690 5794
rect 35310 5742 35362 5794
rect 35982 5742 36034 5794
rect 36654 5742 36706 5794
rect 50318 5742 50370 5794
rect 50878 5742 50930 5794
rect 51774 5742 51826 5794
rect 55246 5742 55298 5794
rect 56814 5742 56866 5794
rect 20750 5630 20802 5682
rect 22094 5630 22146 5682
rect 22430 5630 22482 5682
rect 24670 5630 24722 5682
rect 28702 5630 28754 5682
rect 42590 5630 42642 5682
rect 50878 5630 50930 5682
rect 51774 5630 51826 5682
rect 53902 5630 53954 5682
rect 55246 5630 55298 5682
rect 56030 5630 56082 5682
rect 56814 5630 56866 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 22094 5294 22146 5346
rect 31502 5294 31554 5346
rect 47854 5294 47906 5346
rect 49198 5294 49250 5346
rect 21646 5182 21698 5234
rect 28030 5182 28082 5234
rect 31166 5182 31218 5234
rect 33742 5182 33794 5234
rect 36542 5182 36594 5234
rect 43822 5182 43874 5234
rect 45390 5182 45442 5234
rect 46398 5182 46450 5234
rect 46734 5182 46786 5234
rect 47854 5182 47906 5234
rect 48302 5182 48354 5234
rect 48750 5182 48802 5234
rect 49198 5182 49250 5234
rect 50430 5182 50482 5234
rect 50990 5182 51042 5234
rect 51662 5182 51714 5234
rect 52110 5182 52162 5234
rect 52446 5182 52498 5234
rect 53902 5182 53954 5234
rect 54350 5182 54402 5234
rect 54798 5182 54850 5234
rect 55246 5182 55298 5234
rect 55582 5182 55634 5234
rect 20526 5070 20578 5122
rect 20638 5070 20690 5122
rect 21870 5070 21922 5122
rect 24110 5070 24162 5122
rect 24222 5070 24274 5122
rect 24894 5070 24946 5122
rect 28366 5070 28418 5122
rect 32510 5070 32562 5122
rect 32958 5070 33010 5122
rect 37774 5070 37826 5122
rect 38222 5070 38274 5122
rect 38894 5070 38946 5122
rect 41918 5070 41970 5122
rect 49646 5070 49698 5122
rect 20750 4958 20802 5010
rect 23774 4958 23826 5010
rect 23998 4958 24050 5010
rect 25118 4958 25170 5010
rect 25454 4958 25506 5010
rect 28814 4958 28866 5010
rect 31278 4958 31330 5010
rect 32398 4958 32450 5010
rect 34638 4958 34690 5010
rect 37662 4958 37714 5010
rect 47518 4958 47570 5010
rect 22542 4846 22594 4898
rect 23886 4846 23938 4898
rect 25342 4846 25394 4898
rect 32958 4846 33010 4898
rect 37438 4846 37490 4898
rect 41134 4846 41186 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 3278 4510 3330 4562
rect 33518 4510 33570 4562
rect 37438 4510 37490 4562
rect 37998 4510 38050 4562
rect 38446 4510 38498 4562
rect 38782 4510 38834 4562
rect 46846 4510 46898 4562
rect 47294 4510 47346 4562
rect 47742 4510 47794 4562
rect 54350 4510 54402 4562
rect 2382 4398 2434 4450
rect 2718 4398 2770 4450
rect 26350 4398 26402 4450
rect 30606 4398 30658 4450
rect 39342 4398 39394 4450
rect 39454 4398 39506 4450
rect 48526 4398 48578 4450
rect 57486 4398 57538 4450
rect 21982 4286 22034 4338
rect 22430 4286 22482 4338
rect 23102 4286 23154 4338
rect 26686 4286 26738 4338
rect 28478 4286 28530 4338
rect 29374 4286 29426 4338
rect 30270 4286 30322 4338
rect 31838 4286 31890 4338
rect 32398 4286 32450 4338
rect 34526 4286 34578 4338
rect 34974 4286 35026 4338
rect 40014 4286 40066 4338
rect 48302 4286 48354 4338
rect 54910 4286 54962 4338
rect 56702 4286 56754 4338
rect 57710 4286 57762 4338
rect 23886 4174 23938 4226
rect 28590 4174 28642 4226
rect 28926 4174 28978 4226
rect 32622 4174 32674 4226
rect 55806 4174 55858 4226
rect 39454 4062 39506 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 6974 3614 7026 3666
rect 19294 3614 19346 3666
rect 27582 3614 27634 3666
rect 29374 3614 29426 3666
rect 30270 3614 30322 3666
rect 33182 3614 33234 3666
rect 34526 3614 34578 3666
rect 35646 3614 35698 3666
rect 37102 3614 37154 3666
rect 37550 3614 37602 3666
rect 37998 3614 38050 3666
rect 38446 3614 38498 3666
rect 47966 3614 48018 3666
rect 51326 3614 51378 3666
rect 55246 3614 55298 3666
rect 2830 3502 2882 3554
rect 12238 3502 12290 3554
rect 18734 3502 18786 3554
rect 23662 3502 23714 3554
rect 26798 3502 26850 3554
rect 28478 3502 28530 3554
rect 29822 3502 29874 3554
rect 33854 3502 33906 3554
rect 40014 3502 40066 3554
rect 40910 3502 40962 3554
rect 44270 3502 44322 3554
rect 45166 3502 45218 3554
rect 50654 3502 50706 3554
rect 55918 3502 55970 3554
rect 1934 3390 1986 3442
rect 5070 3390 5122 3442
rect 5854 3390 5906 3442
rect 11118 3390 11170 3442
rect 17614 3390 17666 3442
rect 22542 3390 22594 3442
rect 39118 3390 39170 3442
rect 44942 3278 44994 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 1344 59200 1456 59800
rect 6720 59200 6832 59800
rect 12096 59200 12208 59800
rect 18144 59200 18256 59800
rect 23520 59200 23632 59800
rect 28896 59200 29008 59800
rect 34944 59200 35056 59800
rect 40320 59200 40432 59800
rect 46368 59200 46480 59800
rect 51744 59200 51856 59800
rect 57120 59200 57232 59800
rect 1372 58100 1428 59200
rect 2604 58436 2660 58446
rect 1372 58034 1428 58044
rect 2268 58100 2324 58110
rect 2268 56194 2324 58044
rect 2268 56142 2270 56194
rect 2322 56142 2324 56194
rect 2268 56130 2324 56142
rect 1260 55972 1316 55982
rect 1148 52276 1204 52286
rect 1148 47236 1204 52220
rect 1148 47170 1204 47180
rect 1260 28196 1316 55916
rect 1932 55860 1988 55870
rect 1932 55410 1988 55804
rect 1932 55358 1934 55410
rect 1986 55358 1988 55410
rect 1932 55346 1988 55358
rect 2044 54402 2100 54414
rect 2044 54350 2046 54402
rect 2098 54350 2100 54402
rect 1820 53620 1876 53630
rect 1820 53526 1876 53564
rect 2044 53396 2100 54350
rect 2492 54404 2548 54414
rect 2492 54310 2548 54348
rect 2268 53508 2324 53518
rect 2268 53414 2324 53452
rect 2044 53330 2100 53340
rect 1484 53284 1540 53294
rect 1372 52836 1428 52846
rect 1372 42980 1428 52780
rect 1484 48468 1540 53228
rect 2492 53172 2548 53182
rect 2156 52836 2212 52846
rect 2156 52742 2212 52780
rect 2044 52722 2100 52734
rect 2044 52670 2046 52722
rect 2098 52670 2100 52722
rect 1820 52612 1876 52622
rect 1820 51602 1876 52556
rect 1932 51940 1988 51950
rect 1932 51846 1988 51884
rect 1820 51550 1822 51602
rect 1874 51550 1876 51602
rect 1820 51538 1876 51550
rect 1932 50484 1988 50494
rect 1932 50390 1988 50428
rect 1932 50036 1988 50046
rect 2044 50036 2100 52670
rect 1932 50034 2100 50036
rect 1932 49982 1934 50034
rect 1986 49982 2100 50034
rect 1932 49980 2100 49982
rect 2156 51940 2212 51950
rect 2380 51940 2436 51950
rect 2212 51938 2436 51940
rect 2212 51886 2382 51938
rect 2434 51886 2436 51938
rect 2212 51884 2436 51886
rect 1932 49970 1988 49980
rect 1820 48916 1876 48926
rect 1820 48822 1876 48860
rect 2044 48916 2100 48926
rect 1484 48402 1540 48412
rect 1596 48356 1652 48366
rect 1372 42914 1428 42924
rect 1484 47236 1540 47246
rect 1484 35924 1540 47180
rect 1596 44548 1652 48300
rect 1932 48132 1988 48142
rect 1820 48130 1988 48132
rect 1820 48078 1934 48130
rect 1986 48078 1988 48130
rect 1820 48076 1988 48078
rect 1596 44482 1652 44492
rect 1708 47124 1764 47134
rect 1708 39956 1764 47068
rect 1820 43428 1876 48076
rect 1932 48066 1988 48076
rect 2044 47460 2100 48860
rect 2156 48802 2212 51884
rect 2380 51874 2436 51884
rect 2268 51266 2324 51278
rect 2268 51214 2270 51266
rect 2322 51214 2324 51266
rect 2268 50820 2324 51214
rect 2268 50754 2324 50764
rect 2380 50708 2436 50718
rect 2380 50034 2436 50652
rect 2380 49982 2382 50034
rect 2434 49982 2436 50034
rect 2380 49970 2436 49982
rect 2156 48750 2158 48802
rect 2210 48750 2212 48802
rect 2156 48132 2212 48750
rect 2156 48066 2212 48076
rect 2380 48132 2436 48142
rect 2492 48132 2548 53116
rect 2604 53060 2660 58380
rect 4620 57428 4676 57438
rect 4620 56306 4676 57372
rect 6636 57316 6692 57326
rect 4620 56254 4622 56306
rect 4674 56254 4676 56306
rect 4620 56242 4676 56254
rect 5852 57204 5908 57214
rect 3052 55972 3108 55982
rect 3052 55878 3108 55916
rect 4172 55970 4228 55982
rect 4172 55918 4174 55970
rect 4226 55918 4228 55970
rect 2828 55300 2884 55310
rect 2828 55206 2884 55244
rect 4172 55300 4228 55918
rect 5068 55972 5124 55982
rect 5068 55878 5124 55916
rect 5404 55972 5460 55982
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 5180 55636 5236 55646
rect 4172 55234 4228 55244
rect 5068 55188 5124 55198
rect 5068 55094 5124 55132
rect 3724 55074 3780 55086
rect 3724 55022 3726 55074
rect 3778 55022 3780 55074
rect 3724 54516 3780 55022
rect 4172 55076 4228 55086
rect 4172 55074 4340 55076
rect 4172 55022 4174 55074
rect 4226 55022 4340 55074
rect 4172 55020 4340 55022
rect 4172 55010 4228 55020
rect 3724 54450 3780 54460
rect 3948 54740 4004 54750
rect 2940 54404 2996 54414
rect 3388 54404 3444 54414
rect 3836 54404 3892 54414
rect 2940 54402 3108 54404
rect 2940 54350 2942 54402
rect 2994 54350 3108 54402
rect 2940 54348 3108 54350
rect 2940 54338 2996 54348
rect 2716 53506 2772 53518
rect 2716 53454 2718 53506
rect 2770 53454 2772 53506
rect 2716 53284 2772 53454
rect 2716 53218 2772 53228
rect 2604 53004 2772 53060
rect 2604 52834 2660 52846
rect 2604 52782 2606 52834
rect 2658 52782 2660 52834
rect 2604 52276 2660 52782
rect 2716 52388 2772 53004
rect 2940 52834 2996 52846
rect 2940 52782 2942 52834
rect 2994 52782 2996 52834
rect 2940 52612 2996 52782
rect 2940 52546 2996 52556
rect 2716 52332 2996 52388
rect 2604 52210 2660 52220
rect 2716 52052 2772 52062
rect 2716 51602 2772 51996
rect 2716 51550 2718 51602
rect 2770 51550 2772 51602
rect 2716 51538 2772 51550
rect 2828 51938 2884 51950
rect 2828 51886 2830 51938
rect 2882 51886 2884 51938
rect 2828 50036 2884 51886
rect 2716 49980 2884 50036
rect 2716 49028 2772 49980
rect 2716 48896 2772 48972
rect 2828 49810 2884 49822
rect 2828 49758 2830 49810
rect 2882 49758 2884 49810
rect 2828 49140 2884 49758
rect 2828 48692 2884 49084
rect 2380 48130 2548 48132
rect 2380 48078 2382 48130
rect 2434 48078 2548 48130
rect 2380 48076 2548 48078
rect 2716 48636 2884 48692
rect 1932 47404 2044 47460
rect 1932 46898 1988 47404
rect 2044 47328 2100 47404
rect 2156 47572 2212 47582
rect 1932 46846 1934 46898
rect 1986 46846 1988 46898
rect 1932 46834 1988 46846
rect 1932 46004 1988 46014
rect 1932 45910 1988 45948
rect 1932 44994 1988 45006
rect 1932 44942 1934 44994
rect 1986 44942 1988 44994
rect 1932 44436 1988 44942
rect 1932 44370 1988 44380
rect 2044 44996 2100 45006
rect 2044 44434 2100 44940
rect 2044 44382 2046 44434
rect 2098 44382 2100 44434
rect 2044 44370 2100 44382
rect 1820 43362 1876 43372
rect 1932 43426 1988 43438
rect 1932 43374 1934 43426
rect 1986 43374 1988 43426
rect 1932 43316 1988 43374
rect 1932 43250 1988 43260
rect 2156 43092 2212 47516
rect 2380 47460 2436 48076
rect 2268 47404 2436 47460
rect 2268 46900 2324 47404
rect 2380 47236 2436 47246
rect 2380 47234 2660 47236
rect 2380 47182 2382 47234
rect 2434 47182 2660 47234
rect 2380 47180 2660 47182
rect 2380 47170 2436 47180
rect 2268 46834 2324 46844
rect 2492 47012 2548 47022
rect 2268 46676 2324 46686
rect 2268 46674 2436 46676
rect 2268 46622 2270 46674
rect 2322 46622 2436 46674
rect 2268 46620 2436 46622
rect 2268 46610 2324 46620
rect 2380 43988 2436 46620
rect 2492 45778 2548 46956
rect 2604 46900 2660 47180
rect 2604 46834 2660 46844
rect 2604 46228 2660 46238
rect 2604 46002 2660 46172
rect 2604 45950 2606 46002
rect 2658 45950 2660 46002
rect 2604 45938 2660 45950
rect 2716 46004 2772 48636
rect 2940 48580 2996 52332
rect 3052 51268 3108 54348
rect 3388 54402 3556 54404
rect 3388 54350 3390 54402
rect 3442 54350 3556 54402
rect 3388 54348 3556 54350
rect 3388 54338 3444 54348
rect 3388 53844 3444 53854
rect 3164 53506 3220 53518
rect 3164 53454 3166 53506
rect 3218 53454 3220 53506
rect 3164 52836 3220 53454
rect 3164 51492 3220 52780
rect 3276 52164 3332 52174
rect 3276 52070 3332 52108
rect 3164 51436 3332 51492
rect 3052 51202 3108 51212
rect 3164 51266 3220 51278
rect 3164 51214 3166 51266
rect 3218 51214 3220 51266
rect 3052 50596 3108 50606
rect 3052 50502 3108 50540
rect 3164 50484 3220 51214
rect 3164 50418 3220 50428
rect 3164 49922 3220 49934
rect 3164 49870 3166 49922
rect 3218 49870 3220 49922
rect 3164 49700 3220 49870
rect 3164 49634 3220 49644
rect 3276 49252 3332 51436
rect 3388 49588 3444 53788
rect 3500 53732 3556 54348
rect 3836 54310 3892 54348
rect 3500 53666 3556 53676
rect 3612 53506 3668 53518
rect 3612 53454 3614 53506
rect 3666 53454 3668 53506
rect 3500 53284 3556 53294
rect 3500 53170 3556 53228
rect 3500 53118 3502 53170
rect 3554 53118 3556 53170
rect 3500 53106 3556 53118
rect 3612 53172 3668 53454
rect 3612 53106 3668 53116
rect 3948 53060 4004 54684
rect 4172 54404 4228 54414
rect 3724 53004 4004 53060
rect 4060 54402 4228 54404
rect 4060 54350 4174 54402
rect 4226 54350 4228 54402
rect 4060 54348 4228 54350
rect 4060 54290 4116 54348
rect 4172 54338 4228 54348
rect 4060 54238 4062 54290
rect 4114 54238 4116 54290
rect 4060 53506 4116 54238
rect 4060 53454 4062 53506
rect 4114 53454 4116 53506
rect 3724 52722 3780 53004
rect 3724 52670 3726 52722
rect 3778 52670 3780 52722
rect 3724 52658 3780 52670
rect 3948 52834 4004 52846
rect 3948 52782 3950 52834
rect 4002 52782 4004 52834
rect 3724 51938 3780 51950
rect 3724 51886 3726 51938
rect 3778 51886 3780 51938
rect 3612 51266 3668 51278
rect 3612 51214 3614 51266
rect 3666 51214 3668 51266
rect 3388 49522 3444 49532
rect 3500 51154 3556 51166
rect 3500 51102 3502 51154
rect 3554 51102 3556 51154
rect 3276 49186 3332 49196
rect 3052 48804 3108 48814
rect 3052 48710 3108 48748
rect 2940 48524 3332 48580
rect 3164 48356 3220 48366
rect 2940 48354 3220 48356
rect 2940 48302 3166 48354
rect 3218 48302 3220 48354
rect 2940 48300 3220 48302
rect 2828 48242 2884 48254
rect 2828 48190 2830 48242
rect 2882 48190 2884 48242
rect 2828 47908 2884 48190
rect 2828 47842 2884 47852
rect 2940 47684 2996 48300
rect 3164 48290 3220 48300
rect 2828 47628 2996 47684
rect 3052 47684 3108 47694
rect 2828 47236 2884 47628
rect 3052 47570 3108 47628
rect 3052 47518 3054 47570
rect 3106 47518 3108 47570
rect 3052 47506 3108 47518
rect 3164 47460 3220 47470
rect 3164 47366 3220 47404
rect 3052 47236 3108 47246
rect 2828 47180 2996 47236
rect 2828 46900 2884 46910
rect 2828 46806 2884 46844
rect 2940 46676 2996 47180
rect 3052 47142 3108 47180
rect 3164 46900 3220 46910
rect 3276 46900 3332 48524
rect 3500 47908 3556 51102
rect 3612 50932 3668 51214
rect 3612 50866 3668 50876
rect 3500 47842 3556 47852
rect 3612 50372 3668 50382
rect 3612 48802 3668 50316
rect 3724 50036 3780 51886
rect 3948 51044 4004 52782
rect 4060 51492 4116 53454
rect 4284 53170 4340 55020
rect 4620 55074 4676 55086
rect 4620 55022 4622 55074
rect 4674 55022 4676 55074
rect 4620 54290 4676 55022
rect 5180 54738 5236 55580
rect 5180 54686 5182 54738
rect 5234 54686 5236 54738
rect 5180 54674 5236 54686
rect 4620 54238 4622 54290
rect 4674 54238 4676 54290
rect 4620 54226 4676 54238
rect 4732 54402 4788 54414
rect 4732 54350 4734 54402
rect 4786 54350 4788 54402
rect 4732 54292 4788 54350
rect 4732 54236 5236 54292
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 5068 54068 5124 54078
rect 5068 53842 5124 54012
rect 5068 53790 5070 53842
rect 5122 53790 5124 53842
rect 5068 53778 5124 53790
rect 4508 53508 4564 53518
rect 5180 53508 5236 54236
rect 4508 53506 5012 53508
rect 4508 53454 4510 53506
rect 4562 53454 5012 53506
rect 4508 53452 5012 53454
rect 4508 53442 4564 53452
rect 4284 53118 4286 53170
rect 4338 53118 4340 53170
rect 4284 53060 4340 53118
rect 4284 52994 4340 53004
rect 4844 52834 4900 52846
rect 4844 52782 4846 52834
rect 4898 52782 4900 52834
rect 4172 52722 4228 52734
rect 4172 52670 4174 52722
rect 4226 52670 4228 52722
rect 4172 52388 4228 52670
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4172 52332 4564 52388
rect 4508 52274 4564 52332
rect 4508 52222 4510 52274
rect 4562 52222 4564 52274
rect 4508 52210 4564 52222
rect 4060 51426 4116 51436
rect 4172 51938 4228 51950
rect 4172 51886 4174 51938
rect 4226 51886 4228 51938
rect 4172 51604 4228 51886
rect 4844 51716 4900 52782
rect 4060 51266 4116 51278
rect 4060 51214 4062 51266
rect 4114 51214 4116 51266
rect 4060 51154 4116 51214
rect 4060 51102 4062 51154
rect 4114 51102 4116 51154
rect 4060 51090 4116 51102
rect 3948 50978 4004 50988
rect 3724 49970 3780 49980
rect 3948 50370 4004 50382
rect 3948 50318 3950 50370
rect 4002 50318 4004 50370
rect 3948 50036 4004 50318
rect 4172 50372 4228 51548
rect 4172 50306 4228 50316
rect 4284 51660 4900 51716
rect 4284 50260 4340 51660
rect 4844 51492 4900 51502
rect 4844 51398 4900 51436
rect 4620 51378 4676 51390
rect 4620 51326 4622 51378
rect 4674 51326 4676 51378
rect 4620 51156 4676 51326
rect 4956 51268 5012 53452
rect 5180 53442 5236 53452
rect 5404 52948 5460 55916
rect 5516 55748 5572 55758
rect 5516 54068 5572 55692
rect 5852 55410 5908 57148
rect 5852 55358 5854 55410
rect 5906 55358 5908 55410
rect 5852 55346 5908 55358
rect 5964 56196 6020 56206
rect 5516 54002 5572 54012
rect 5628 54402 5684 54414
rect 5628 54350 5630 54402
rect 5682 54350 5684 54402
rect 5628 53844 5684 54350
rect 5628 53778 5684 53788
rect 5740 53732 5796 53742
rect 5740 53638 5796 53676
rect 5964 53508 6020 56140
rect 6076 55972 6132 55982
rect 6076 55878 6132 55916
rect 6524 55972 6580 55982
rect 6524 55878 6580 55916
rect 6300 55074 6356 55086
rect 6300 55022 6302 55074
rect 6354 55022 6356 55074
rect 6300 54852 6356 55022
rect 6300 54786 6356 54796
rect 6076 54404 6132 54414
rect 6076 54402 6468 54404
rect 6076 54350 6078 54402
rect 6130 54350 6468 54402
rect 6076 54348 6468 54350
rect 6076 54338 6132 54348
rect 5740 53452 6020 53508
rect 6076 53732 6132 53742
rect 5628 53172 5684 53182
rect 5628 53078 5684 53116
rect 5404 52892 5684 52948
rect 5292 52834 5348 52846
rect 5292 52782 5294 52834
rect 5346 52782 5348 52834
rect 5180 52276 5236 52286
rect 4956 51202 5012 51212
rect 5068 52162 5124 52174
rect 5068 52110 5070 52162
rect 5122 52110 5124 52162
rect 5068 52052 5124 52110
rect 4620 51100 4900 51156
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4844 50820 4900 51100
rect 5068 51044 5124 51996
rect 5068 50978 5124 50988
rect 4844 50764 5124 50820
rect 4396 50594 4452 50606
rect 4396 50542 4398 50594
rect 4450 50542 4452 50594
rect 4396 50484 4452 50542
rect 4396 50418 4452 50428
rect 4620 50594 4676 50606
rect 4620 50542 4622 50594
rect 4674 50542 4676 50594
rect 4508 50372 4564 50382
rect 4508 50278 4564 50316
rect 4284 50194 4340 50204
rect 3948 49970 4004 49980
rect 4060 50036 4116 50046
rect 4060 50034 4452 50036
rect 4060 49982 4062 50034
rect 4114 49982 4452 50034
rect 4060 49980 4452 49982
rect 4060 49970 4116 49980
rect 3724 49810 3780 49822
rect 3724 49758 3726 49810
rect 3778 49758 3780 49810
rect 3724 49138 3780 49758
rect 3724 49086 3726 49138
rect 3778 49086 3780 49138
rect 3724 49074 3780 49086
rect 3948 49812 4004 49822
rect 3612 48750 3614 48802
rect 3666 48750 3668 48802
rect 3612 47068 3668 48750
rect 3164 46898 3332 46900
rect 3164 46846 3166 46898
rect 3218 46846 3332 46898
rect 3164 46844 3332 46846
rect 3500 47012 3668 47068
rect 3724 48804 3780 48814
rect 3164 46834 3220 46844
rect 3052 46788 3108 46798
rect 3052 46676 3108 46732
rect 3052 46620 3220 46676
rect 2940 46610 2996 46620
rect 2716 45948 2996 46004
rect 2492 45726 2494 45778
rect 2546 45726 2548 45778
rect 2492 45714 2548 45726
rect 2716 45778 2772 45790
rect 2716 45726 2718 45778
rect 2770 45726 2772 45778
rect 2716 45444 2772 45726
rect 2716 45378 2772 45388
rect 2828 45108 2884 45118
rect 2828 45014 2884 45052
rect 2492 44548 2548 44558
rect 2492 44434 2548 44492
rect 2492 44382 2494 44434
rect 2546 44382 2548 44434
rect 2492 44370 2548 44382
rect 2940 44324 2996 45948
rect 2940 44192 2996 44268
rect 3164 43988 3220 46620
rect 3500 46452 3556 47012
rect 3500 46386 3556 46396
rect 3612 46900 3668 46910
rect 3612 46114 3668 46844
rect 3724 46340 3780 48748
rect 3836 48804 3892 48814
rect 3948 48804 4004 49756
rect 4060 49810 4116 49822
rect 4284 49812 4340 49822
rect 4060 49758 4062 49810
rect 4114 49758 4116 49810
rect 4060 49700 4116 49758
rect 4060 49634 4116 49644
rect 4172 49810 4340 49812
rect 4172 49758 4286 49810
rect 4338 49758 4340 49810
rect 4172 49756 4340 49758
rect 4060 49476 4116 49486
rect 4060 48914 4116 49420
rect 4060 48862 4062 48914
rect 4114 48862 4116 48914
rect 4060 48850 4116 48862
rect 3836 48802 4004 48804
rect 3836 48750 3838 48802
rect 3890 48750 4004 48802
rect 3836 48748 4004 48750
rect 3836 48738 3892 48748
rect 4172 48580 4228 49756
rect 4284 49746 4340 49756
rect 4396 49588 4452 49980
rect 4060 48524 4228 48580
rect 4284 49532 4452 49588
rect 4620 49588 4676 50542
rect 4844 50596 4900 50606
rect 4844 50594 5012 50596
rect 4844 50542 4846 50594
rect 4898 50542 5012 50594
rect 4844 50540 5012 50542
rect 4844 50530 4900 50540
rect 4956 49812 5012 50540
rect 5068 50484 5124 50764
rect 5068 50418 5124 50428
rect 4956 49746 5012 49756
rect 3948 48020 4004 48030
rect 3948 47926 4004 47964
rect 3836 46676 3892 46686
rect 3836 46582 3892 46620
rect 3948 46676 4004 46686
rect 4060 46676 4116 48524
rect 4284 48468 4340 49532
rect 4620 49522 4676 49532
rect 5068 49698 5124 49710
rect 5068 49646 5070 49698
rect 5122 49646 5124 49698
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4844 49252 4900 49262
rect 4620 49250 4900 49252
rect 4620 49198 4846 49250
rect 4898 49198 4900 49250
rect 4620 49196 4900 49198
rect 4620 48804 4676 49196
rect 4844 49186 4900 49196
rect 4844 49028 4900 49038
rect 4732 48916 4788 48926
rect 4732 48822 4788 48860
rect 4844 48914 4900 48972
rect 4844 48862 4846 48914
rect 4898 48862 4900 48914
rect 4844 48850 4900 48862
rect 4620 48738 4676 48748
rect 5068 48692 5124 49646
rect 5068 48626 5124 48636
rect 4284 48402 4340 48412
rect 4844 48468 4900 48478
rect 4844 48374 4900 48412
rect 4172 48354 4228 48366
rect 4172 48302 4174 48354
rect 4226 48302 4228 48354
rect 4172 47012 4228 48302
rect 4284 48244 4340 48254
rect 4284 48130 4340 48188
rect 5068 48244 5124 48254
rect 5068 48150 5124 48188
rect 4284 48078 4286 48130
rect 4338 48078 4340 48130
rect 4284 48066 4340 48078
rect 4956 48130 5012 48142
rect 4956 48078 4958 48130
rect 5010 48078 5012 48130
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4508 47572 4564 47582
rect 4508 47478 4564 47516
rect 4732 47460 4788 47470
rect 4172 46956 4452 47012
rect 4284 46788 4340 46798
rect 4284 46694 4340 46732
rect 3948 46674 4116 46676
rect 3948 46622 3950 46674
rect 4002 46622 4116 46674
rect 3948 46620 4116 46622
rect 3724 46274 3780 46284
rect 3948 46228 4004 46620
rect 4396 46564 4452 46956
rect 4284 46508 4452 46564
rect 3948 46162 4004 46172
rect 4172 46452 4228 46462
rect 3612 46062 3614 46114
rect 3666 46062 3668 46114
rect 3388 45892 3444 45902
rect 3388 45798 3444 45836
rect 3612 45892 3668 46062
rect 3612 45826 3668 45836
rect 3836 46116 3892 46126
rect 3836 45890 3892 46060
rect 3836 45838 3838 45890
rect 3890 45838 3892 45890
rect 3836 45826 3892 45838
rect 4060 45780 4116 45790
rect 3724 45666 3780 45678
rect 3724 45614 3726 45666
rect 3778 45614 3780 45666
rect 2380 43932 3108 43988
rect 2716 43764 2772 43774
rect 1820 43036 2212 43092
rect 2268 43540 2324 43550
rect 1820 40964 1876 43036
rect 2268 42980 2324 43484
rect 2380 43428 2436 43438
rect 2380 43426 2548 43428
rect 2380 43374 2382 43426
rect 2434 43374 2548 43426
rect 2380 43372 2548 43374
rect 2380 43362 2436 43372
rect 2268 42924 2436 42980
rect 2268 42756 2324 42766
rect 2156 42644 2212 42682
rect 2156 42578 2212 42588
rect 2156 42420 2212 42430
rect 1932 41858 1988 41870
rect 1932 41806 1934 41858
rect 1986 41806 1988 41858
rect 1932 41748 1988 41806
rect 1932 41682 1988 41692
rect 1820 40898 1876 40908
rect 1820 40628 1876 40638
rect 1820 40534 1876 40572
rect 2156 40404 2212 42364
rect 2268 41298 2324 42700
rect 2380 42754 2436 42924
rect 2380 42702 2382 42754
rect 2434 42702 2436 42754
rect 2380 42690 2436 42702
rect 2380 41860 2436 41870
rect 2380 41766 2436 41804
rect 2268 41246 2270 41298
rect 2322 41246 2324 41298
rect 2268 41234 2324 41246
rect 2492 41300 2548 43372
rect 2604 42868 2660 42878
rect 2604 42774 2660 42812
rect 2716 42754 2772 43708
rect 2828 43652 2884 43662
rect 2828 43558 2884 43596
rect 2716 42702 2718 42754
rect 2770 42702 2772 42754
rect 2716 42690 2772 42702
rect 2940 43540 2996 43550
rect 2828 42644 2884 42654
rect 2828 42196 2884 42588
rect 2716 42140 2828 42196
rect 2492 41244 2660 41300
rect 2492 41074 2548 41086
rect 2492 41022 2494 41074
rect 2546 41022 2548 41074
rect 2268 40962 2324 40974
rect 2268 40910 2270 40962
rect 2322 40910 2324 40962
rect 2268 40628 2324 40910
rect 2268 40572 2436 40628
rect 2268 40404 2324 40414
rect 2156 40402 2324 40404
rect 2156 40350 2270 40402
rect 2322 40350 2324 40402
rect 2156 40348 2324 40350
rect 2268 40338 2324 40348
rect 2380 40292 2436 40572
rect 2380 40226 2436 40236
rect 2492 40516 2548 41022
rect 1708 39900 2212 39956
rect 1484 35858 1540 35868
rect 1596 39620 1652 39630
rect 1596 29428 1652 39564
rect 1932 39506 1988 39518
rect 1932 39454 1934 39506
rect 1986 39454 1988 39506
rect 1932 39060 1988 39454
rect 2156 39060 2212 39900
rect 1932 38994 1988 39004
rect 2044 39058 2212 39060
rect 2044 39006 2158 39058
rect 2210 39006 2212 39058
rect 2044 39004 2212 39006
rect 1820 38948 1876 38958
rect 1820 38668 1876 38892
rect 1932 38836 1988 38874
rect 1932 38770 1988 38780
rect 1820 38612 1988 38668
rect 1820 38274 1876 38286
rect 1820 38222 1822 38274
rect 1874 38222 1876 38274
rect 1708 37380 1764 37390
rect 1708 29652 1764 37324
rect 1820 37378 1876 38222
rect 1932 38162 1988 38612
rect 1932 38110 1934 38162
rect 1986 38110 1988 38162
rect 1932 38098 1988 38110
rect 1820 37326 1822 37378
rect 1874 37326 1876 37378
rect 1820 37314 1876 37326
rect 1932 36708 1988 36718
rect 1820 36596 1876 36606
rect 1820 36502 1876 36540
rect 1820 35924 1876 35934
rect 1932 35924 1988 36652
rect 1820 35922 1988 35924
rect 1820 35870 1822 35922
rect 1874 35870 1988 35922
rect 1820 35868 1988 35870
rect 1820 35858 1876 35868
rect 1820 34692 1876 34702
rect 1820 32788 1876 34636
rect 1932 34018 1988 34030
rect 1932 33966 1934 34018
rect 1986 33966 1988 34018
rect 1932 33684 1988 33966
rect 1932 33618 1988 33628
rect 1932 33460 1988 33470
rect 1932 33366 1988 33404
rect 1932 32788 1988 32798
rect 1820 32786 1988 32788
rect 1820 32734 1934 32786
rect 1986 32734 1988 32786
rect 1820 32732 1988 32734
rect 1820 31666 1876 32732
rect 1932 32722 1988 32732
rect 2044 31948 2100 39004
rect 2156 38994 2212 39004
rect 2156 38500 2212 38510
rect 2156 37490 2212 38444
rect 2156 37438 2158 37490
rect 2210 37438 2212 37490
rect 2156 37426 2212 37438
rect 2268 38274 2324 38286
rect 2268 38222 2270 38274
rect 2322 38222 2324 38274
rect 2268 36706 2324 38222
rect 2380 37940 2436 37950
rect 2380 37846 2436 37884
rect 2492 37828 2548 40460
rect 2604 39060 2660 41244
rect 2604 38994 2660 39004
rect 2716 38500 2772 42140
rect 2828 42102 2884 42140
rect 2940 40514 2996 43484
rect 3052 41188 3108 43932
rect 3164 42868 3220 43932
rect 3276 45108 3332 45118
rect 3276 44212 3332 45052
rect 3276 44098 3332 44156
rect 3276 44046 3278 44098
rect 3330 44046 3332 44098
rect 3276 43876 3332 44046
rect 3276 43820 3556 43876
rect 3276 43538 3332 43550
rect 3276 43486 3278 43538
rect 3330 43486 3332 43538
rect 3276 43092 3332 43486
rect 3276 43026 3332 43036
rect 3164 42812 3332 42868
rect 3164 42084 3220 42094
rect 3164 41990 3220 42028
rect 3052 41132 3220 41188
rect 3052 40964 3108 40974
rect 3052 40870 3108 40908
rect 2940 40462 2942 40514
rect 2994 40462 2996 40514
rect 2940 39732 2996 40462
rect 2828 39620 2884 39630
rect 2828 39526 2884 39564
rect 2828 38724 2884 38734
rect 2940 38724 2996 39676
rect 2828 38722 2996 38724
rect 2828 38670 2830 38722
rect 2882 38670 2996 38722
rect 2828 38668 2996 38670
rect 3052 40290 3108 40302
rect 3052 40238 3054 40290
rect 3106 40238 3108 40290
rect 2828 38658 2884 38668
rect 2716 38434 2772 38444
rect 2604 38276 2660 38286
rect 2604 38274 2884 38276
rect 2604 38222 2606 38274
rect 2658 38222 2884 38274
rect 2604 38220 2884 38222
rect 2604 38210 2660 38220
rect 2828 38050 2884 38220
rect 2828 37998 2830 38050
rect 2882 37998 2884 38050
rect 2828 37986 2884 37998
rect 2492 37772 2884 37828
rect 2716 37380 2772 37390
rect 2716 37266 2772 37324
rect 2716 37214 2718 37266
rect 2770 37214 2772 37266
rect 2716 37202 2772 37214
rect 2268 36654 2270 36706
rect 2322 36654 2324 36706
rect 2268 36642 2324 36654
rect 2380 36372 2436 36382
rect 2268 35924 2324 35934
rect 2268 35830 2324 35868
rect 2156 34916 2212 34926
rect 2156 34822 2212 34860
rect 2380 33908 2436 36316
rect 2380 33842 2436 33852
rect 2492 36148 2548 36158
rect 2380 33684 2436 33694
rect 2380 33458 2436 33628
rect 2380 33406 2382 33458
rect 2434 33406 2436 33458
rect 2380 33394 2436 33406
rect 2492 33236 2548 36092
rect 2716 35474 2772 35486
rect 2716 35422 2718 35474
rect 2770 35422 2772 35474
rect 2716 35140 2772 35422
rect 2828 35476 2884 37772
rect 2940 36372 2996 36382
rect 2940 36278 2996 36316
rect 3052 36148 3108 40238
rect 3164 39172 3220 41132
rect 3164 39106 3220 39116
rect 3052 36082 3108 36092
rect 3164 38836 3220 38846
rect 3052 35700 3108 35710
rect 3164 35700 3220 38780
rect 3276 38164 3332 42812
rect 3388 41300 3444 41310
rect 3388 41074 3444 41244
rect 3388 41022 3390 41074
rect 3442 41022 3444 41074
rect 3388 41010 3444 41022
rect 3500 40852 3556 43820
rect 3612 43650 3668 43662
rect 3612 43598 3614 43650
rect 3666 43598 3668 43650
rect 3612 43204 3668 43598
rect 3724 43316 3780 45614
rect 3948 45108 4004 45118
rect 3948 45014 4004 45052
rect 3948 44324 4004 44334
rect 3724 43250 3780 43260
rect 3836 44098 3892 44110
rect 3836 44046 3838 44098
rect 3890 44046 3892 44098
rect 3612 42980 3668 43148
rect 3612 42924 3780 42980
rect 3612 42756 3668 42766
rect 3612 42662 3668 42700
rect 3724 42644 3780 42924
rect 3836 42868 3892 44046
rect 3836 42736 3892 42812
rect 3724 42578 3780 42588
rect 3836 42308 3892 42318
rect 3836 42194 3892 42252
rect 3836 42142 3838 42194
rect 3890 42142 3892 42194
rect 3276 38032 3332 38108
rect 3388 40796 3556 40852
rect 3724 41300 3780 41310
rect 3276 37268 3332 37278
rect 3276 37174 3332 37212
rect 3276 36372 3332 36382
rect 3276 36278 3332 36316
rect 3052 35698 3332 35700
rect 3052 35646 3054 35698
rect 3106 35646 3332 35698
rect 3052 35644 3332 35646
rect 3052 35634 3108 35644
rect 3052 35476 3108 35486
rect 2828 35474 3108 35476
rect 2828 35422 3054 35474
rect 3106 35422 3108 35474
rect 2828 35420 3108 35422
rect 2716 35074 2772 35084
rect 2940 35252 2996 35262
rect 2604 34692 2660 34702
rect 2604 34598 2660 34636
rect 2940 34690 2996 35196
rect 2940 34638 2942 34690
rect 2994 34638 2996 34690
rect 2828 34132 2884 34142
rect 2380 33180 2548 33236
rect 2604 34130 2884 34132
rect 2604 34078 2830 34130
rect 2882 34078 2884 34130
rect 2604 34076 2884 34078
rect 2044 31892 2324 31948
rect 1820 31614 1822 31666
rect 1874 31614 1876 31666
rect 1820 31602 1876 31614
rect 2156 31666 2212 31678
rect 2156 31614 2158 31666
rect 2210 31614 2212 31666
rect 1932 31332 1988 31342
rect 1932 30436 1988 31276
rect 2044 31220 2100 31230
rect 2044 31126 2100 31164
rect 2156 30884 2212 31614
rect 2268 31332 2324 31892
rect 2268 31266 2324 31276
rect 2380 31108 2436 33180
rect 2380 31042 2436 31052
rect 2492 33012 2548 33022
rect 2492 30996 2548 32956
rect 2604 31108 2660 34076
rect 2828 34066 2884 34076
rect 2940 33796 2996 34638
rect 2940 33730 2996 33740
rect 2940 33346 2996 33358
rect 2940 33294 2942 33346
rect 2994 33294 2996 33346
rect 2716 32562 2772 32574
rect 2716 32510 2718 32562
rect 2770 32510 2772 32562
rect 2716 31668 2772 32510
rect 2940 32564 2996 33294
rect 3052 33012 3108 35420
rect 3164 35140 3220 35150
rect 3164 33684 3220 35084
rect 3164 33234 3220 33628
rect 3276 33460 3332 35644
rect 3276 33394 3332 33404
rect 3164 33182 3166 33234
rect 3218 33182 3220 33234
rect 3164 33170 3220 33182
rect 3276 33236 3332 33246
rect 3276 33012 3332 33180
rect 3052 32946 3108 32956
rect 3164 32956 3332 33012
rect 2828 31780 2884 31790
rect 2940 31780 2996 32508
rect 2828 31778 2996 31780
rect 2828 31726 2830 31778
rect 2882 31726 2996 31778
rect 2828 31724 2996 31726
rect 3052 31892 3108 31902
rect 2828 31714 2884 31724
rect 2716 31602 2772 31612
rect 3052 31666 3108 31836
rect 3052 31614 3054 31666
rect 3106 31614 3108 31666
rect 3052 31602 3108 31614
rect 3164 31444 3220 32956
rect 3388 32676 3444 40796
rect 3724 40628 3780 41244
rect 3724 40562 3780 40572
rect 3836 41188 3892 42142
rect 3836 40180 3892 41132
rect 3612 40124 3892 40180
rect 3948 40402 4004 44268
rect 4060 44212 4116 45724
rect 4172 45556 4228 46396
rect 4284 46004 4340 46508
rect 4732 46452 4788 47404
rect 4956 47124 5012 48078
rect 5180 47348 5236 52220
rect 5292 51828 5348 52782
rect 5628 51940 5684 52892
rect 5740 52052 5796 53452
rect 5964 52948 6020 52958
rect 5852 52276 5908 52286
rect 5852 52182 5908 52220
rect 5740 51996 5908 52052
rect 5628 51874 5684 51884
rect 5292 51762 5348 51772
rect 5628 51716 5684 51726
rect 5404 51604 5460 51614
rect 5404 51490 5460 51548
rect 5404 51438 5406 51490
rect 5458 51438 5460 51490
rect 5404 51426 5460 51438
rect 5292 51156 5348 51166
rect 5292 49700 5348 51100
rect 5628 50148 5684 51660
rect 5740 51604 5796 51614
rect 5740 51510 5796 51548
rect 5852 51492 5908 51996
rect 5852 51426 5908 51436
rect 5852 50820 5908 50830
rect 5964 50820 6020 52892
rect 5852 50818 6020 50820
rect 5852 50766 5854 50818
rect 5906 50766 6020 50818
rect 5852 50764 6020 50766
rect 5852 50754 5908 50764
rect 5964 50484 6020 50522
rect 5964 50418 6020 50428
rect 6076 50428 6132 53676
rect 6300 53506 6356 53518
rect 6300 53454 6302 53506
rect 6354 53454 6356 53506
rect 6188 53172 6244 53182
rect 6188 53078 6244 53116
rect 6300 52836 6356 53454
rect 6300 52770 6356 52780
rect 6412 50820 6468 54348
rect 6524 54402 6580 54414
rect 6524 54350 6526 54402
rect 6578 54350 6580 54402
rect 6524 54180 6580 54350
rect 6524 54114 6580 54124
rect 6524 53620 6580 53630
rect 6636 53620 6692 57260
rect 6748 56642 6804 59200
rect 10892 58212 10948 58222
rect 7532 57988 7588 57998
rect 6748 56590 6750 56642
rect 6802 56590 6804 56642
rect 6748 56578 6804 56590
rect 7420 57876 7476 57886
rect 7196 56082 7252 56094
rect 7196 56030 7198 56082
rect 7250 56030 7252 56082
rect 6860 55300 6916 55310
rect 6748 55076 6804 55086
rect 6748 54982 6804 55020
rect 6748 53620 6804 53630
rect 6636 53564 6748 53620
rect 6524 53170 6580 53564
rect 6748 53488 6804 53564
rect 6524 53118 6526 53170
rect 6578 53118 6580 53170
rect 6524 52276 6580 53118
rect 6524 52210 6580 52220
rect 6636 52052 6692 52062
rect 6524 51940 6580 51950
rect 6524 51602 6580 51884
rect 6524 51550 6526 51602
rect 6578 51550 6580 51602
rect 6524 51538 6580 51550
rect 6412 50754 6468 50764
rect 6636 50706 6692 51996
rect 6860 51940 6916 55244
rect 7196 55186 7252 56030
rect 7196 55134 7198 55186
rect 7250 55134 7252 55186
rect 7196 55122 7252 55134
rect 7420 54740 7476 57820
rect 7532 55298 7588 57932
rect 9324 57652 9380 57662
rect 7868 57540 7924 57550
rect 7644 56642 7700 56654
rect 7644 56590 7646 56642
rect 7698 56590 7700 56642
rect 7644 55970 7700 56590
rect 7644 55918 7646 55970
rect 7698 55918 7700 55970
rect 7644 55906 7700 55918
rect 7532 55246 7534 55298
rect 7586 55246 7588 55298
rect 7532 55234 7588 55246
rect 7420 54738 7812 54740
rect 7420 54686 7422 54738
rect 7474 54686 7812 54738
rect 7420 54684 7812 54686
rect 7420 54674 7476 54684
rect 6972 54402 7028 54414
rect 6972 54350 6974 54402
rect 7026 54350 7028 54402
rect 6972 53956 7028 54350
rect 6972 53890 7028 53900
rect 6972 53730 7028 53742
rect 6972 53678 6974 53730
rect 7026 53678 7028 53730
rect 6972 52948 7028 53678
rect 7756 53732 7812 54684
rect 7644 53620 7700 53630
rect 7644 53526 7700 53564
rect 7756 53618 7812 53676
rect 7756 53566 7758 53618
rect 7810 53566 7812 53618
rect 7756 53554 7812 53566
rect 7308 53058 7364 53070
rect 7308 53006 7310 53058
rect 7362 53006 7364 53058
rect 6972 52882 7028 52892
rect 7196 52948 7252 52958
rect 7308 52948 7364 53006
rect 7308 52892 7700 52948
rect 7196 52854 7252 52892
rect 7308 52722 7364 52734
rect 7308 52670 7310 52722
rect 7362 52670 7364 52722
rect 7196 52500 7252 52510
rect 6972 52276 7028 52286
rect 6972 52162 7028 52220
rect 7196 52164 7252 52444
rect 6972 52110 6974 52162
rect 7026 52110 7028 52162
rect 6972 52098 7028 52110
rect 7084 52162 7252 52164
rect 7084 52110 7198 52162
rect 7250 52110 7252 52162
rect 7084 52108 7252 52110
rect 6636 50654 6638 50706
rect 6690 50654 6692 50706
rect 5852 50372 5908 50382
rect 6076 50372 6244 50428
rect 5852 50278 5908 50316
rect 6188 50148 6244 50372
rect 5628 50092 5796 50148
rect 5740 50036 5796 50092
rect 6076 50092 6244 50148
rect 5852 50036 5908 50046
rect 5740 50034 5908 50036
rect 5740 49982 5854 50034
rect 5906 49982 5908 50034
rect 5740 49980 5908 49982
rect 5628 49924 5684 49934
rect 5404 49700 5460 49710
rect 5292 49698 5572 49700
rect 5292 49646 5406 49698
rect 5458 49646 5572 49698
rect 5292 49644 5572 49646
rect 5404 49634 5460 49644
rect 5404 48356 5460 48366
rect 5404 48242 5460 48300
rect 5404 48190 5406 48242
rect 5458 48190 5460 48242
rect 5404 48020 5460 48190
rect 5404 47954 5460 47964
rect 5180 47292 5348 47348
rect 5068 47236 5124 47246
rect 5068 47234 5236 47236
rect 5068 47182 5070 47234
rect 5122 47182 5236 47234
rect 5068 47180 5236 47182
rect 5068 47170 5124 47180
rect 4844 47068 5012 47124
rect 4844 47012 4900 47068
rect 4844 46946 4900 46956
rect 4956 46900 5012 46910
rect 4732 46396 4900 46452
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4620 46116 4676 46126
rect 4284 45938 4340 45948
rect 4508 46004 4564 46014
rect 4508 45910 4564 45948
rect 4172 45490 4228 45500
rect 4396 45892 4452 45902
rect 4284 45220 4340 45230
rect 4396 45220 4452 45836
rect 4620 45890 4676 46060
rect 4620 45838 4622 45890
rect 4674 45838 4676 45890
rect 4620 45826 4676 45838
rect 4284 45218 4452 45220
rect 4284 45166 4286 45218
rect 4338 45166 4452 45218
rect 4284 45164 4452 45166
rect 4508 45332 4564 45342
rect 4284 45154 4340 45164
rect 4172 44994 4228 45006
rect 4172 44942 4174 44994
rect 4226 44942 4228 44994
rect 4172 44884 4228 44942
rect 4508 44884 4564 45276
rect 4844 45220 4900 46396
rect 4956 45892 5012 46844
rect 5068 46564 5124 46574
rect 5068 46470 5124 46508
rect 5180 46450 5236 47180
rect 5180 46398 5182 46450
rect 5234 46398 5236 46450
rect 5180 46386 5236 46398
rect 5292 46116 5348 47292
rect 5404 47012 5460 47022
rect 5404 46898 5460 46956
rect 5404 46846 5406 46898
rect 5458 46846 5460 46898
rect 5404 46834 5460 46846
rect 5292 46050 5348 46060
rect 4956 45890 5348 45892
rect 4956 45838 4958 45890
rect 5010 45838 5348 45890
rect 4956 45836 5348 45838
rect 4956 45826 5012 45836
rect 5292 45330 5348 45836
rect 5292 45278 5294 45330
rect 5346 45278 5348 45330
rect 5292 45266 5348 45278
rect 5404 45780 5460 45790
rect 4844 45164 5012 45220
rect 4172 44818 4228 44828
rect 4284 44828 4564 44884
rect 4844 44994 4900 45006
rect 4844 44942 4846 44994
rect 4898 44942 4900 44994
rect 4844 44884 4900 44942
rect 4172 44212 4228 44222
rect 4060 44210 4228 44212
rect 4060 44158 4174 44210
rect 4226 44158 4228 44210
rect 4060 44156 4228 44158
rect 4172 44146 4228 44156
rect 4172 43540 4228 43550
rect 4172 43446 4228 43484
rect 4172 42082 4228 42094
rect 4172 42030 4174 42082
rect 4226 42030 4228 42082
rect 4172 41972 4228 42030
rect 4172 41906 4228 41916
rect 4060 41076 4116 41086
rect 4060 40982 4116 41020
rect 4284 40740 4340 44828
rect 4844 44818 4900 44828
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4508 44548 4564 44558
rect 4508 43762 4564 44492
rect 4508 43710 4510 43762
rect 4562 43710 4564 43762
rect 4508 43698 4564 43710
rect 4844 43204 4900 43214
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4508 42980 4564 42990
rect 4844 42980 4900 43148
rect 4508 42978 4900 42980
rect 4508 42926 4510 42978
rect 4562 42926 4900 42978
rect 4508 42924 4900 42926
rect 4508 42914 4564 42924
rect 4620 42754 4676 42766
rect 4620 42702 4622 42754
rect 4674 42702 4676 42754
rect 4620 41972 4676 42702
rect 4844 42084 4900 42094
rect 4620 41906 4676 41916
rect 4732 41970 4788 41982
rect 4732 41918 4734 41970
rect 4786 41918 4788 41970
rect 4732 41860 4788 41918
rect 4732 41794 4788 41804
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4620 41188 4676 41198
rect 4620 41094 4676 41132
rect 4732 41076 4788 41086
rect 4844 41076 4900 42028
rect 4956 41300 5012 45164
rect 5068 44098 5124 44110
rect 5068 44046 5070 44098
rect 5122 44046 5124 44098
rect 5068 41972 5124 44046
rect 5292 43764 5348 43774
rect 5180 43426 5236 43438
rect 5180 43374 5182 43426
rect 5234 43374 5236 43426
rect 5180 43314 5236 43374
rect 5180 43262 5182 43314
rect 5234 43262 5236 43314
rect 5180 43250 5236 43262
rect 5068 41916 5236 41972
rect 4956 41234 5012 41244
rect 5068 41748 5124 41758
rect 4788 41020 4900 41076
rect 4732 41010 4788 41020
rect 4284 40674 4340 40684
rect 4508 40964 4564 40974
rect 3948 40350 3950 40402
rect 4002 40350 4004 40402
rect 3500 39620 3556 39630
rect 3500 37380 3556 39564
rect 3500 37314 3556 37324
rect 3612 35810 3668 40124
rect 3724 39844 3780 39854
rect 3724 39730 3780 39788
rect 3724 39678 3726 39730
rect 3778 39678 3780 39730
rect 3724 37492 3780 39678
rect 3836 39732 3892 39742
rect 3836 39618 3892 39676
rect 3836 39566 3838 39618
rect 3890 39566 3892 39618
rect 3836 39554 3892 39566
rect 3948 39620 4004 40350
rect 4508 40402 4564 40908
rect 4508 40350 4510 40402
rect 4562 40350 4564 40402
rect 4508 40338 4564 40350
rect 4284 40292 4340 40302
rect 3948 39554 4004 39564
rect 4172 39732 4228 39742
rect 4172 39618 4228 39676
rect 4172 39566 4174 39618
rect 4226 39566 4228 39618
rect 4172 39554 4228 39566
rect 3836 39172 3892 39182
rect 3836 38948 3892 39116
rect 3836 38854 3892 38892
rect 4172 39060 4228 39070
rect 4172 38164 4228 39004
rect 4284 38836 4340 40236
rect 4844 40068 4900 41020
rect 4956 41076 5012 41086
rect 4956 40982 5012 41020
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4844 40002 4900 40012
rect 4956 40740 5012 40750
rect 4476 39946 4740 39956
rect 4956 39844 5012 40684
rect 4284 38722 4340 38780
rect 4284 38670 4286 38722
rect 4338 38670 4340 38722
rect 4284 38658 4340 38670
rect 4844 39788 5012 39844
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4172 38108 4452 38164
rect 4284 37938 4340 37950
rect 4284 37886 4286 37938
rect 4338 37886 4340 37938
rect 3948 37828 4004 37838
rect 3948 37734 4004 37772
rect 3836 37492 3892 37502
rect 3724 37490 3892 37492
rect 3724 37438 3838 37490
rect 3890 37438 3892 37490
rect 3724 37436 3892 37438
rect 3836 37426 3892 37436
rect 4284 37268 4340 37886
rect 4396 37490 4452 38108
rect 4844 37492 4900 39788
rect 4956 39394 5012 39406
rect 4956 39342 4958 39394
rect 5010 39342 5012 39394
rect 4956 39284 5012 39342
rect 4956 39218 5012 39228
rect 5068 39060 5124 41692
rect 5180 39732 5236 41916
rect 5180 39666 5236 39676
rect 4396 37438 4398 37490
rect 4450 37438 4452 37490
rect 4396 37426 4452 37438
rect 4732 37436 4900 37492
rect 4956 39004 5124 39060
rect 5180 39508 5236 39518
rect 4956 37828 5012 39004
rect 5180 38948 5236 39452
rect 5068 38892 5236 38948
rect 5068 38162 5124 38892
rect 5180 38724 5236 38762
rect 5180 38658 5236 38668
rect 5068 38110 5070 38162
rect 5122 38110 5124 38162
rect 5068 38098 5124 38110
rect 5180 38500 5236 38510
rect 4956 37492 5012 37772
rect 5180 37828 5236 38444
rect 4956 37436 5124 37492
rect 4172 37266 4340 37268
rect 4172 37214 4286 37266
rect 4338 37214 4340 37266
rect 4172 37212 4340 37214
rect 4060 36708 4116 36718
rect 4060 36614 4116 36652
rect 4172 36372 4228 37212
rect 4284 37202 4340 37212
rect 4508 37268 4564 37278
rect 4508 37174 4564 37212
rect 4732 37044 4788 37436
rect 3948 36260 4004 36270
rect 3948 35922 4004 36204
rect 3948 35870 3950 35922
rect 4002 35870 4004 35922
rect 3948 35858 4004 35870
rect 3612 35758 3614 35810
rect 3666 35758 3668 35810
rect 3500 35028 3556 35038
rect 3500 34690 3556 34972
rect 3500 34638 3502 34690
rect 3554 34638 3556 34690
rect 3500 33012 3556 34638
rect 3612 34356 3668 35758
rect 4172 35810 4228 36316
rect 4172 35758 4174 35810
rect 4226 35758 4228 35810
rect 4172 35746 4228 35758
rect 4284 36988 4788 37044
rect 4844 37266 4900 37278
rect 4844 37214 4846 37266
rect 4898 37214 4900 37266
rect 3836 35698 3892 35710
rect 3836 35646 3838 35698
rect 3890 35646 3892 35698
rect 3836 34916 3892 35646
rect 3612 33348 3668 34300
rect 3724 34914 3892 34916
rect 3724 34862 3838 34914
rect 3890 34862 3892 34914
rect 3724 34860 3892 34862
rect 3724 34130 3780 34860
rect 3836 34850 3892 34860
rect 3724 34078 3726 34130
rect 3778 34078 3780 34130
rect 3724 33570 3780 34078
rect 3948 34242 4004 34254
rect 3948 34190 3950 34242
rect 4002 34190 4004 34242
rect 3948 34020 4004 34190
rect 3948 33954 4004 33964
rect 4172 34132 4228 34142
rect 3724 33518 3726 33570
rect 3778 33518 3780 33570
rect 3724 33506 3780 33518
rect 3612 33282 3668 33292
rect 4060 33460 4116 33470
rect 3836 33236 3892 33246
rect 3836 33234 4004 33236
rect 3836 33182 3838 33234
rect 3890 33182 4004 33234
rect 3836 33180 4004 33182
rect 3836 33170 3892 33180
rect 3500 32956 3892 33012
rect 3612 32676 3668 32686
rect 3388 32620 3556 32676
rect 3276 32564 3332 32574
rect 3276 32470 3332 32508
rect 3052 31388 3220 31444
rect 3388 32452 3444 32462
rect 2940 31108 2996 31118
rect 2604 31052 2772 31108
rect 2492 30930 2548 30940
rect 2380 30884 2436 30894
rect 2156 30882 2436 30884
rect 2156 30830 2382 30882
rect 2434 30830 2436 30882
rect 2156 30828 2436 30830
rect 1932 30380 2212 30436
rect 1932 30212 1988 30222
rect 1932 30118 1988 30156
rect 1708 29586 1764 29596
rect 1596 29362 1652 29372
rect 1932 29316 1988 29326
rect 2044 29316 2100 29326
rect 1932 29314 2044 29316
rect 1932 29262 1934 29314
rect 1986 29262 2044 29314
rect 1932 29260 2044 29262
rect 1932 29250 1988 29260
rect 1260 28130 1316 28140
rect 1932 27746 1988 27758
rect 1932 27694 1934 27746
rect 1986 27694 1988 27746
rect 1932 27636 1988 27694
rect 1932 27570 1988 27580
rect 1932 22260 1988 22270
rect 1932 22166 1988 22204
rect 2044 20188 2100 29260
rect 2156 28644 2212 30380
rect 2268 29876 2324 30828
rect 2380 30818 2436 30828
rect 2716 30436 2772 31052
rect 2380 30380 2772 30436
rect 2828 30884 2884 30894
rect 2380 30098 2436 30380
rect 2380 30046 2382 30098
rect 2434 30046 2436 30098
rect 2380 30034 2436 30046
rect 2716 30098 2772 30110
rect 2716 30046 2718 30098
rect 2770 30046 2772 30098
rect 2716 29988 2772 30046
rect 2716 29922 2772 29932
rect 2268 29820 2436 29876
rect 2268 29314 2324 29326
rect 2268 29262 2270 29314
rect 2322 29262 2324 29314
rect 2268 29202 2324 29262
rect 2268 29150 2270 29202
rect 2322 29150 2324 29202
rect 2268 29138 2324 29150
rect 2156 28588 2324 28644
rect 2156 28420 2212 28430
rect 2156 28326 2212 28364
rect 2156 27188 2212 27198
rect 2268 27188 2324 28588
rect 2380 28084 2436 29820
rect 2828 29650 2884 30828
rect 2828 29598 2830 29650
rect 2882 29598 2884 29650
rect 2828 29586 2884 29598
rect 2604 28756 2660 28766
rect 2604 28662 2660 28700
rect 2380 28018 2436 28028
rect 2156 27186 2324 27188
rect 2156 27134 2158 27186
rect 2210 27134 2324 27186
rect 2156 27132 2324 27134
rect 2156 27122 2212 27132
rect 2940 24948 2996 31052
rect 3052 29202 3108 31388
rect 3164 31220 3220 31230
rect 3164 31126 3220 31164
rect 3276 29988 3332 29998
rect 3276 29894 3332 29932
rect 3276 29652 3332 29662
rect 3276 29558 3332 29596
rect 3052 29150 3054 29202
rect 3106 29150 3108 29202
rect 3052 28754 3108 29150
rect 3388 29202 3444 32396
rect 3388 29150 3390 29202
rect 3442 29150 3444 29202
rect 3388 29138 3444 29150
rect 3500 28866 3556 32620
rect 3612 32452 3668 32620
rect 3612 32386 3668 32396
rect 3612 31668 3668 31678
rect 3612 31218 3668 31612
rect 3612 31166 3614 31218
rect 3666 31166 3668 31218
rect 3612 30770 3668 31166
rect 3612 30718 3614 30770
rect 3666 30718 3668 30770
rect 3612 30706 3668 30718
rect 3724 30434 3780 30446
rect 3724 30382 3726 30434
rect 3778 30382 3780 30434
rect 3724 30322 3780 30382
rect 3724 30270 3726 30322
rect 3778 30270 3780 30322
rect 3724 30212 3780 30270
rect 3724 30146 3780 30156
rect 3500 28814 3502 28866
rect 3554 28814 3556 28866
rect 3500 28802 3556 28814
rect 3612 29652 3668 29662
rect 3052 28702 3054 28754
rect 3106 28702 3108 28754
rect 3052 28690 3108 28702
rect 3612 28754 3668 29596
rect 3836 29540 3892 32956
rect 3948 32674 4004 33180
rect 3948 32622 3950 32674
rect 4002 32622 4004 32674
rect 3948 32564 4004 32622
rect 3948 32498 4004 32508
rect 3948 31668 4004 31678
rect 4060 31668 4116 33404
rect 3948 31666 4116 31668
rect 3948 31614 3950 31666
rect 4002 31614 4116 31666
rect 3948 31612 4116 31614
rect 3948 30434 4004 31612
rect 4172 31108 4228 34076
rect 4284 32788 4340 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4508 36482 4564 36494
rect 4508 36430 4510 36482
rect 4562 36430 4564 36482
rect 4508 36372 4564 36430
rect 4732 36484 4788 36494
rect 4844 36484 4900 37214
rect 4732 36482 4900 36484
rect 4732 36430 4734 36482
rect 4786 36430 4900 36482
rect 4732 36428 4900 36430
rect 4732 36418 4788 36428
rect 4508 36306 4564 36316
rect 4732 35924 4788 35934
rect 4732 35830 4788 35868
rect 4844 35364 4900 36428
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4844 35298 4900 35308
rect 4956 37268 5012 37278
rect 4956 36482 5012 37212
rect 4956 36430 4958 36482
rect 5010 36430 5012 36482
rect 4476 35242 4740 35252
rect 4732 34916 4788 34926
rect 4956 34916 5012 36430
rect 5068 35252 5124 37436
rect 5068 35186 5124 35196
rect 4396 34356 4452 34366
rect 4396 34262 4452 34300
rect 4732 33908 4788 34860
rect 4844 34860 5012 34916
rect 4844 34132 4900 34860
rect 4956 34690 5012 34702
rect 4956 34638 4958 34690
rect 5010 34638 5012 34690
rect 4956 34580 5012 34638
rect 4956 34514 5012 34524
rect 5180 34468 5236 37772
rect 5292 36148 5348 43708
rect 5404 42980 5460 45724
rect 5516 45668 5572 49644
rect 5628 49364 5684 49868
rect 5628 47570 5684 49308
rect 5628 47518 5630 47570
rect 5682 47518 5684 47570
rect 5628 47506 5684 47518
rect 5740 47682 5796 47694
rect 5740 47630 5742 47682
rect 5794 47630 5796 47682
rect 5628 47348 5684 47358
rect 5628 47124 5684 47292
rect 5628 47058 5684 47068
rect 5516 45602 5572 45612
rect 5628 46788 5684 46798
rect 5628 45444 5684 46732
rect 5740 46676 5796 47630
rect 5852 46788 5908 49980
rect 5964 49140 6020 49150
rect 5964 49046 6020 49084
rect 5852 46732 6020 46788
rect 5740 46610 5796 46620
rect 5852 46562 5908 46574
rect 5852 46510 5854 46562
rect 5906 46510 5908 46562
rect 5740 46450 5796 46462
rect 5740 46398 5742 46450
rect 5794 46398 5796 46450
rect 5740 45668 5796 46398
rect 5852 46116 5908 46510
rect 5964 46340 6020 46732
rect 5964 46274 6020 46284
rect 5852 46060 6020 46116
rect 5852 45668 5908 45678
rect 5740 45666 5908 45668
rect 5740 45614 5854 45666
rect 5906 45614 5908 45666
rect 5740 45612 5908 45614
rect 5740 45444 5796 45454
rect 5628 45388 5740 45444
rect 5628 45106 5684 45118
rect 5628 45054 5630 45106
rect 5682 45054 5684 45106
rect 5628 44100 5684 45054
rect 5628 44034 5684 44044
rect 5740 44210 5796 45388
rect 5740 44158 5742 44210
rect 5794 44158 5796 44210
rect 5516 43428 5572 43438
rect 5516 43334 5572 43372
rect 5404 42868 5460 42924
rect 5628 42868 5684 42878
rect 5404 42866 5684 42868
rect 5404 42814 5630 42866
rect 5682 42814 5684 42866
rect 5404 42812 5684 42814
rect 5628 42802 5684 42812
rect 5516 42084 5572 42122
rect 5516 42018 5572 42028
rect 5292 36082 5348 36092
rect 5516 41860 5572 41870
rect 5180 34402 5236 34412
rect 5292 35812 5348 35822
rect 5516 35812 5572 41804
rect 5740 41748 5796 44158
rect 5852 43764 5908 45612
rect 5964 44772 6020 46060
rect 6076 45108 6132 50092
rect 6188 49252 6244 49262
rect 6188 47570 6244 49196
rect 6524 49026 6580 49038
rect 6524 48974 6526 49026
rect 6578 48974 6580 49026
rect 6412 48356 6468 48366
rect 6412 48262 6468 48300
rect 6300 48242 6356 48254
rect 6300 48190 6302 48242
rect 6354 48190 6356 48242
rect 6300 47682 6356 48190
rect 6300 47630 6302 47682
rect 6354 47630 6356 47682
rect 6300 47618 6356 47630
rect 6188 47518 6190 47570
rect 6242 47518 6244 47570
rect 6188 47506 6244 47518
rect 6412 47460 6468 47470
rect 6412 46900 6468 47404
rect 6524 47236 6580 48974
rect 6636 48468 6692 50654
rect 6636 48402 6692 48412
rect 6748 51884 6916 51940
rect 6636 48244 6692 48254
rect 6636 48150 6692 48188
rect 6636 47236 6692 47246
rect 6524 47234 6692 47236
rect 6524 47182 6638 47234
rect 6690 47182 6692 47234
rect 6524 47180 6692 47182
rect 6636 47124 6692 47180
rect 6636 47058 6692 47068
rect 6300 46844 6468 46900
rect 6076 45042 6132 45052
rect 6188 46116 6244 46126
rect 5964 44706 6020 44716
rect 6076 44882 6132 44894
rect 6076 44830 6078 44882
rect 6130 44830 6132 44882
rect 5964 44100 6020 44110
rect 5964 44006 6020 44044
rect 5852 43698 5908 43708
rect 6076 43652 6132 44830
rect 5964 43596 6132 43652
rect 6188 44210 6244 46060
rect 6300 45890 6356 46844
rect 6524 46788 6580 46798
rect 6524 46694 6580 46732
rect 6412 46676 6468 46686
rect 6412 46582 6468 46620
rect 6524 46452 6580 46462
rect 6636 46452 6692 46462
rect 6524 46450 6636 46452
rect 6524 46398 6526 46450
rect 6578 46398 6636 46450
rect 6524 46396 6636 46398
rect 6748 46452 6804 51884
rect 6860 51716 6916 51726
rect 6860 51602 6916 51660
rect 6860 51550 6862 51602
rect 6914 51550 6916 51602
rect 6860 51538 6916 51550
rect 7084 50708 7140 52108
rect 7196 52098 7252 52108
rect 7308 51604 7364 52670
rect 7532 52164 7588 52174
rect 7420 52052 7476 52062
rect 7532 52052 7588 52108
rect 7420 52050 7588 52052
rect 7420 51998 7422 52050
rect 7474 51998 7588 52050
rect 7420 51996 7588 51998
rect 7420 51986 7476 51996
rect 7644 51940 7700 52892
rect 7644 51874 7700 51884
rect 7756 52836 7812 52846
rect 7308 51538 7364 51548
rect 7420 51492 7476 51502
rect 7084 50652 7252 50708
rect 7084 50372 7140 50382
rect 7084 50278 7140 50316
rect 6860 49924 6916 49934
rect 6860 49810 6916 49868
rect 6860 49758 6862 49810
rect 6914 49758 6916 49810
rect 6860 49252 6916 49758
rect 7084 49812 7140 49822
rect 6972 49586 7028 49598
rect 6972 49534 6974 49586
rect 7026 49534 7028 49586
rect 6972 49476 7028 49534
rect 6972 49410 7028 49420
rect 6860 49186 6916 49196
rect 6972 49026 7028 49038
rect 6972 48974 6974 49026
rect 7026 48974 7028 49026
rect 6860 48580 6916 48590
rect 6860 48354 6916 48524
rect 6860 48302 6862 48354
rect 6914 48302 6916 48354
rect 6860 47460 6916 48302
rect 6972 48356 7028 48974
rect 7084 49028 7140 49756
rect 7084 48962 7140 48972
rect 6972 48290 7028 48300
rect 7196 48020 7252 50652
rect 7420 50484 7476 51436
rect 7420 50418 7476 50428
rect 7644 51044 7700 51054
rect 7532 50372 7588 50382
rect 7532 49812 7588 50316
rect 7532 49718 7588 49756
rect 7644 49252 7700 50988
rect 7644 49186 7700 49196
rect 7644 49028 7700 49038
rect 7644 48934 7700 48972
rect 7756 48466 7812 52780
rect 7868 51490 7924 57484
rect 9212 56308 9268 56318
rect 8988 55970 9044 55982
rect 8988 55918 8990 55970
rect 9042 55918 9044 55970
rect 8988 55860 9044 55918
rect 8988 55794 9044 55804
rect 8092 55074 8148 55086
rect 8092 55022 8094 55074
rect 8146 55022 8148 55074
rect 7980 54402 8036 54414
rect 7980 54350 7982 54402
rect 8034 54350 8036 54402
rect 7980 54068 8036 54350
rect 7980 54002 8036 54012
rect 7980 53508 8036 53518
rect 7980 53414 8036 53452
rect 8092 53172 8148 55022
rect 8540 55074 8596 55086
rect 8540 55022 8542 55074
rect 8594 55022 8596 55074
rect 8540 54740 8596 55022
rect 8876 55074 8932 55086
rect 8876 55022 8878 55074
rect 8930 55022 8932 55074
rect 8540 54674 8596 54684
rect 8652 54964 8708 54974
rect 8652 54738 8708 54908
rect 8876 54852 8932 55022
rect 8876 54786 8932 54796
rect 8652 54686 8654 54738
rect 8706 54686 8708 54738
rect 8652 54674 8708 54686
rect 8428 54514 8484 54526
rect 8428 54462 8430 54514
rect 8482 54462 8484 54514
rect 8092 53106 8148 53116
rect 8204 54404 8260 54414
rect 8092 52948 8148 52958
rect 8204 52948 8260 54348
rect 8428 53844 8484 54462
rect 9100 54514 9156 54526
rect 9100 54462 9102 54514
rect 9154 54462 9156 54514
rect 8428 53778 8484 53788
rect 8540 54402 8596 54414
rect 8540 54350 8542 54402
rect 8594 54350 8596 54402
rect 8540 53620 8596 54350
rect 9100 54404 9156 54462
rect 9100 54338 9156 54348
rect 9100 53844 9156 53854
rect 9100 53750 9156 53788
rect 8428 53564 8596 53620
rect 8428 53508 8484 53564
rect 8652 53508 8708 53518
rect 8092 52946 8204 52948
rect 8092 52894 8094 52946
rect 8146 52894 8204 52946
rect 8092 52892 8204 52894
rect 8092 52882 8148 52892
rect 8204 52816 8260 52892
rect 8316 53452 8484 53508
rect 8540 53506 8708 53508
rect 8540 53454 8654 53506
rect 8706 53454 8708 53506
rect 8540 53452 8708 53454
rect 8204 52388 8260 52398
rect 8092 52164 8148 52174
rect 7868 51438 7870 51490
rect 7922 51438 7924 51490
rect 7868 51426 7924 51438
rect 7980 51492 8036 51502
rect 7980 51398 8036 51436
rect 8092 51490 8148 52108
rect 8204 52162 8260 52332
rect 8204 52110 8206 52162
rect 8258 52110 8260 52162
rect 8204 52052 8260 52110
rect 8204 51986 8260 51996
rect 8316 52050 8372 53452
rect 8540 52724 8596 53452
rect 8652 53442 8708 53452
rect 8876 53508 8932 53518
rect 8540 52658 8596 52668
rect 8652 52834 8708 52846
rect 8652 52782 8654 52834
rect 8706 52782 8708 52834
rect 8316 51998 8318 52050
rect 8370 51998 8372 52050
rect 8316 51986 8372 51998
rect 8652 51940 8708 52782
rect 8876 52162 8932 53452
rect 8876 52110 8878 52162
rect 8930 52110 8932 52162
rect 8876 52098 8932 52110
rect 9100 52834 9156 52846
rect 9100 52782 9102 52834
rect 9154 52782 9156 52834
rect 9100 52164 9156 52782
rect 9100 52098 9156 52108
rect 8092 51438 8094 51490
rect 8146 51438 8148 51490
rect 8092 51426 8148 51438
rect 8428 51884 8708 51940
rect 8764 52050 8820 52062
rect 8764 51998 8766 52050
rect 8818 51998 8820 52050
rect 8316 51380 8372 51390
rect 8428 51380 8484 51884
rect 8540 51604 8596 51614
rect 8764 51604 8820 51998
rect 9100 51940 9156 51950
rect 9212 51940 9268 56252
rect 9100 51938 9268 51940
rect 9100 51886 9102 51938
rect 9154 51886 9268 51938
rect 9100 51884 9268 51886
rect 9324 53620 9380 57596
rect 10444 56084 10500 56094
rect 9772 55970 9828 55982
rect 9772 55918 9774 55970
rect 9826 55918 9828 55970
rect 9772 55524 9828 55918
rect 10220 55972 10276 55982
rect 10220 55878 10276 55916
rect 9772 55458 9828 55468
rect 10444 55300 10500 56028
rect 10668 56084 10724 56094
rect 10668 55970 10724 56028
rect 10668 55918 10670 55970
rect 10722 55918 10724 55970
rect 10668 55748 10724 55918
rect 10668 55682 10724 55692
rect 10444 55244 10836 55300
rect 9436 55188 9492 55198
rect 9436 55094 9492 55132
rect 9884 55188 9940 55198
rect 9772 55074 9828 55086
rect 9772 55022 9774 55074
rect 9826 55022 9828 55074
rect 9772 54964 9828 55022
rect 9772 54898 9828 54908
rect 9884 54626 9940 55132
rect 9884 54574 9886 54626
rect 9938 54574 9940 54626
rect 9772 54404 9828 54414
rect 9436 53956 9492 53966
rect 9436 53862 9492 53900
rect 9772 53732 9828 54348
rect 9884 54068 9940 54574
rect 9884 54002 9940 54012
rect 10108 55076 10164 55086
rect 9884 53732 9940 53742
rect 9772 53730 9940 53732
rect 9772 53678 9886 53730
rect 9938 53678 9940 53730
rect 9772 53676 9940 53678
rect 9884 53666 9940 53676
rect 9324 53618 9828 53620
rect 9324 53566 9326 53618
rect 9378 53566 9828 53618
rect 9324 53564 9828 53566
rect 9100 51874 9156 51884
rect 9212 51716 9268 51726
rect 9324 51716 9380 53564
rect 9772 53170 9828 53564
rect 10108 53618 10164 55020
rect 10332 54628 10388 54638
rect 10332 54534 10388 54572
rect 10444 54626 10500 55244
rect 10668 55076 10724 55086
rect 10444 54574 10446 54626
rect 10498 54574 10500 54626
rect 10444 54562 10500 54574
rect 10556 55074 10724 55076
rect 10556 55022 10670 55074
rect 10722 55022 10724 55074
rect 10556 55020 10724 55022
rect 10220 54514 10276 54526
rect 10220 54462 10222 54514
rect 10274 54462 10276 54514
rect 10220 53844 10276 54462
rect 10556 54404 10612 55020
rect 10668 55010 10724 55020
rect 10444 54348 10612 54404
rect 10444 53844 10500 54348
rect 10220 53788 10500 53844
rect 10108 53566 10110 53618
rect 10162 53566 10164 53618
rect 10108 53554 10164 53566
rect 10220 53618 10276 53630
rect 10220 53566 10222 53618
rect 10274 53566 10276 53618
rect 9772 53118 9774 53170
rect 9826 53118 9828 53170
rect 9772 53106 9828 53118
rect 10220 52836 10276 53566
rect 10220 52770 10276 52780
rect 10332 52834 10388 52846
rect 10332 52782 10334 52834
rect 10386 52782 10388 52834
rect 9996 52612 10052 52622
rect 9996 52162 10052 52556
rect 9996 52110 9998 52162
rect 10050 52110 10052 52162
rect 9996 51828 10052 52110
rect 9996 51762 10052 51772
rect 8540 51602 8820 51604
rect 8540 51550 8542 51602
rect 8594 51550 8820 51602
rect 8540 51548 8820 51550
rect 8988 51660 9212 51716
rect 9268 51660 9380 51716
rect 8988 51602 9044 51660
rect 8988 51550 8990 51602
rect 9042 51550 9044 51602
rect 9212 51584 9268 51660
rect 9884 51604 9940 51614
rect 8540 51538 8596 51548
rect 8988 51538 9044 51550
rect 9884 51510 9940 51548
rect 9996 51380 10052 51390
rect 8428 51324 8596 51380
rect 8316 51268 8372 51324
rect 8316 51212 8484 51268
rect 7980 51156 8036 51166
rect 7756 48414 7758 48466
rect 7810 48414 7812 48466
rect 7756 48402 7812 48414
rect 7868 50370 7924 50382
rect 7868 50318 7870 50370
rect 7922 50318 7924 50370
rect 7420 48356 7476 48366
rect 7420 48262 7476 48300
rect 6860 47394 6916 47404
rect 6972 47964 7252 48020
rect 6972 47346 7028 47964
rect 7868 47460 7924 50318
rect 7980 49140 8036 51100
rect 8204 50820 8260 50830
rect 8204 50706 8260 50764
rect 8204 50654 8206 50706
rect 8258 50654 8260 50706
rect 8204 50642 8260 50654
rect 8092 50484 8148 50494
rect 8092 49810 8148 50428
rect 8092 49758 8094 49810
rect 8146 49758 8148 49810
rect 8092 49746 8148 49758
rect 7980 49074 8036 49084
rect 8204 49252 8260 49262
rect 7980 48914 8036 48926
rect 7980 48862 7982 48914
rect 8034 48862 8036 48914
rect 7980 47908 8036 48862
rect 7980 47842 8036 47852
rect 7756 47404 7924 47460
rect 7980 47460 8036 47470
rect 6972 47294 6974 47346
rect 7026 47294 7028 47346
rect 6972 47282 7028 47294
rect 7308 47348 7364 47358
rect 6748 46396 7140 46452
rect 6524 46386 6580 46396
rect 6300 45838 6302 45890
rect 6354 45838 6356 45890
rect 6300 45332 6356 45838
rect 6300 45266 6356 45276
rect 6412 46228 6468 46238
rect 6300 44994 6356 45006
rect 6300 44942 6302 44994
rect 6354 44942 6356 44994
rect 6300 44882 6356 44942
rect 6300 44830 6302 44882
rect 6354 44830 6356 44882
rect 6300 44818 6356 44830
rect 6300 44660 6356 44670
rect 6300 44546 6356 44604
rect 6300 44494 6302 44546
rect 6354 44494 6356 44546
rect 6300 44482 6356 44494
rect 6412 44324 6468 46172
rect 6188 44158 6190 44210
rect 6242 44158 6244 44210
rect 5740 41682 5796 41692
rect 5852 43540 5908 43550
rect 5852 41076 5908 43484
rect 5964 42196 6020 43596
rect 6076 43428 6132 43438
rect 6076 43334 6132 43372
rect 5964 42140 6132 42196
rect 5964 41970 6020 41982
rect 5964 41918 5966 41970
rect 6018 41918 6020 41970
rect 5964 41860 6020 41918
rect 5964 41794 6020 41804
rect 6076 41524 6132 42140
rect 6188 41860 6244 44158
rect 6300 44268 6468 44324
rect 6636 44324 6692 46396
rect 6860 46228 6916 46238
rect 6860 45890 6916 46172
rect 6860 45838 6862 45890
rect 6914 45838 6916 45890
rect 6860 45826 6916 45838
rect 6748 45666 6804 45678
rect 6748 45614 6750 45666
rect 6802 45614 6804 45666
rect 6748 45556 6804 45614
rect 6972 45668 7028 45678
rect 6972 45574 7028 45612
rect 6748 45490 6804 45500
rect 6300 42532 6356 44268
rect 6636 44258 6692 44268
rect 6748 45220 6804 45230
rect 6748 43876 6804 45164
rect 6972 45220 7028 45230
rect 6972 45126 7028 45164
rect 6860 45108 6916 45118
rect 6860 44660 6916 45052
rect 7084 45108 7140 46396
rect 7308 46004 7364 47292
rect 7196 45948 7364 46004
rect 7420 46564 7476 46574
rect 7196 45556 7252 45948
rect 7196 45490 7252 45500
rect 7308 45668 7364 45678
rect 7084 45106 7252 45108
rect 7084 45054 7086 45106
rect 7138 45054 7252 45106
rect 7084 45052 7252 45054
rect 7084 45042 7140 45052
rect 6860 44594 6916 44604
rect 6860 44436 6916 44446
rect 6860 44342 6916 44380
rect 6972 44322 7028 44334
rect 6972 44270 6974 44322
rect 7026 44270 7028 44322
rect 6972 43988 7028 44270
rect 6972 43922 7028 43932
rect 6748 43810 6804 43820
rect 6524 43426 6580 43438
rect 6524 43374 6526 43426
rect 6578 43374 6580 43426
rect 6524 42980 6580 43374
rect 6972 43426 7028 43438
rect 6972 43374 6974 43426
rect 7026 43374 7028 43426
rect 6636 43314 6692 43326
rect 6636 43262 6638 43314
rect 6690 43262 6692 43314
rect 6636 42980 6692 43262
rect 6748 42980 6804 42990
rect 6636 42924 6748 42980
rect 6524 42914 6580 42924
rect 6748 42914 6804 42924
rect 6412 42868 6468 42878
rect 6412 42754 6468 42812
rect 6412 42702 6414 42754
rect 6466 42702 6468 42754
rect 6412 42690 6468 42702
rect 6748 42756 6804 42766
rect 6524 42642 6580 42654
rect 6524 42590 6526 42642
rect 6578 42590 6580 42642
rect 6300 42530 6468 42532
rect 6300 42478 6302 42530
rect 6354 42478 6468 42530
rect 6300 42476 6468 42478
rect 6300 42466 6356 42476
rect 6300 41972 6356 41982
rect 6300 41878 6356 41916
rect 6188 41794 6244 41804
rect 6076 41458 6132 41468
rect 5964 41300 6020 41310
rect 5964 41206 6020 41244
rect 5852 41020 6020 41076
rect 5852 40402 5908 40414
rect 5852 40350 5854 40402
rect 5906 40350 5908 40402
rect 5740 38836 5796 38874
rect 5852 38836 5908 40350
rect 5796 38780 5908 38836
rect 5740 38770 5796 38780
rect 5852 38050 5908 38780
rect 5964 39730 6020 41020
rect 6412 40516 6468 42476
rect 6524 41636 6580 42590
rect 6636 42644 6692 42682
rect 6748 42662 6804 42700
rect 6636 42578 6692 42588
rect 6524 41570 6580 41580
rect 6860 42082 6916 42094
rect 6860 42030 6862 42082
rect 6914 42030 6916 42082
rect 6860 41300 6916 42030
rect 6412 40450 6468 40460
rect 6636 41188 6692 41198
rect 5964 39678 5966 39730
rect 6018 39678 6020 39730
rect 5964 38388 6020 39678
rect 6524 39394 6580 39406
rect 6524 39342 6526 39394
rect 6578 39342 6580 39394
rect 5964 38322 6020 38332
rect 6076 38946 6132 38958
rect 6076 38894 6078 38946
rect 6130 38894 6132 38946
rect 6076 38612 6132 38894
rect 6300 38836 6356 38846
rect 6524 38836 6580 39342
rect 6300 38834 6580 38836
rect 6300 38782 6302 38834
rect 6354 38782 6580 38834
rect 6300 38780 6580 38782
rect 6300 38668 6356 38780
rect 6300 38612 6468 38668
rect 5852 37998 5854 38050
rect 5906 37998 5908 38050
rect 5852 37986 5908 37998
rect 5740 37940 5796 37950
rect 5740 37266 5796 37884
rect 5852 37828 5908 37838
rect 5852 37734 5908 37772
rect 5740 37214 5742 37266
rect 5794 37214 5796 37266
rect 5740 37202 5796 37214
rect 6076 36932 6132 38556
rect 6412 37938 6468 38612
rect 6412 37886 6414 37938
rect 6466 37886 6468 37938
rect 6076 36866 6132 36876
rect 6300 37266 6356 37278
rect 6300 37214 6302 37266
rect 6354 37214 6356 37266
rect 6076 36596 6132 36606
rect 6076 36502 6132 36540
rect 6300 36372 6356 37214
rect 6412 36484 6468 37886
rect 6412 36418 6468 36428
rect 6300 36306 6356 36316
rect 6412 36260 6468 36270
rect 6412 36258 6580 36260
rect 6412 36206 6414 36258
rect 6466 36206 6580 36258
rect 6412 36204 6580 36206
rect 6412 36194 6468 36204
rect 5292 35810 5572 35812
rect 5292 35758 5294 35810
rect 5346 35758 5572 35810
rect 5292 35756 5572 35758
rect 6524 35812 6580 36204
rect 4956 34356 5012 34366
rect 4956 34262 5012 34300
rect 4844 34076 5012 34132
rect 4732 33852 4900 33908
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4620 33460 4676 33470
rect 4620 33366 4676 33404
rect 4284 32732 4452 32788
rect 4284 32564 4340 32574
rect 4284 32470 4340 32508
rect 4396 32340 4452 32732
rect 4284 32284 4452 32340
rect 4284 31220 4340 32284
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4732 31780 4788 31790
rect 4844 31780 4900 33852
rect 4956 33684 5012 34076
rect 4956 33628 5124 33684
rect 4956 33460 5012 33470
rect 4956 32674 5012 33404
rect 4956 32622 4958 32674
rect 5010 32622 5012 32674
rect 4956 32610 5012 32622
rect 5068 32340 5124 33628
rect 5180 32340 5236 32350
rect 5068 32338 5236 32340
rect 5068 32286 5182 32338
rect 5234 32286 5236 32338
rect 5068 32284 5236 32286
rect 5292 32340 5348 35756
rect 6524 35746 6580 35756
rect 5628 35700 5684 35710
rect 6300 35700 6356 35710
rect 5628 35698 6468 35700
rect 5628 35646 5630 35698
rect 5682 35646 6302 35698
rect 6354 35646 6468 35698
rect 5628 35644 6468 35646
rect 5628 35634 5684 35644
rect 6300 35634 6356 35644
rect 5628 35476 5684 35486
rect 5516 35252 5572 35262
rect 5516 34468 5572 35196
rect 5628 35026 5684 35420
rect 5628 34974 5630 35026
rect 5682 34974 5684 35026
rect 5628 34962 5684 34974
rect 5852 34916 5908 34926
rect 5516 34402 5572 34412
rect 5740 34692 5796 34702
rect 5404 34356 5460 34366
rect 5404 34262 5460 34300
rect 5740 34354 5796 34636
rect 5740 34302 5742 34354
rect 5794 34302 5796 34354
rect 5740 34290 5796 34302
rect 5516 34244 5572 34254
rect 5404 32564 5460 32574
rect 5404 32470 5460 32508
rect 5292 32284 5460 32340
rect 5180 32004 5236 32284
rect 5180 31938 5236 31948
rect 4732 31778 4900 31780
rect 4732 31726 4734 31778
rect 4786 31726 4900 31778
rect 4732 31724 4900 31726
rect 4284 31164 4676 31220
rect 4172 31052 4340 31108
rect 3948 30382 3950 30434
rect 4002 30382 4004 30434
rect 3948 30370 4004 30382
rect 4172 30882 4228 30894
rect 4172 30830 4174 30882
rect 4226 30830 4228 30882
rect 4172 30770 4228 30830
rect 4172 30718 4174 30770
rect 4226 30718 4228 30770
rect 4172 30212 4228 30718
rect 4284 30436 4340 31052
rect 4620 30772 4676 31164
rect 4732 31218 4788 31724
rect 4956 31668 5012 31678
rect 4956 31574 5012 31612
rect 4732 31166 4734 31218
rect 4786 31166 4788 31218
rect 4732 31154 4788 31166
rect 4956 31444 5012 31454
rect 4620 30716 4900 30772
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4284 30380 4788 30436
rect 4172 30146 4228 30156
rect 4284 29986 4340 29998
rect 4284 29934 4286 29986
rect 4338 29934 4340 29986
rect 4284 29764 4340 29934
rect 4284 29698 4340 29708
rect 4620 29986 4676 29998
rect 4620 29934 4622 29986
rect 4674 29934 4676 29986
rect 4284 29540 4340 29550
rect 3836 29538 4340 29540
rect 3836 29486 4286 29538
rect 4338 29486 4340 29538
rect 3836 29484 4340 29486
rect 4284 29474 4340 29484
rect 3612 28702 3614 28754
rect 3666 28702 3668 28754
rect 3612 28690 3668 28702
rect 3724 29428 3780 29438
rect 3724 29314 3780 29372
rect 4620 29428 4676 29934
rect 4732 29650 4788 30380
rect 4732 29598 4734 29650
rect 4786 29598 4788 29650
rect 4732 29586 4788 29598
rect 4844 29652 4900 30716
rect 4844 29586 4900 29596
rect 4956 29428 5012 31388
rect 5068 30996 5124 31006
rect 5068 30902 5124 30940
rect 4620 29372 5012 29428
rect 5068 29988 5124 29998
rect 4620 29316 4676 29372
rect 3724 29262 3726 29314
rect 3778 29262 3780 29314
rect 3276 28644 3332 28654
rect 3052 28084 3108 28094
rect 3052 27858 3108 28028
rect 3052 27806 3054 27858
rect 3106 27806 3108 27858
rect 3052 27794 3108 27806
rect 3276 25172 3332 28588
rect 3500 28084 3556 28094
rect 3500 27990 3556 28028
rect 3276 25106 3332 25116
rect 2940 24882 2996 24892
rect 2828 22372 2884 22382
rect 2380 22370 2884 22372
rect 2380 22318 2830 22370
rect 2882 22318 2884 22370
rect 2380 22316 2884 22318
rect 2380 20690 2436 22316
rect 2828 22306 2884 22316
rect 2380 20638 2382 20690
rect 2434 20638 2436 20690
rect 2380 20626 2436 20638
rect 2716 20690 2772 20702
rect 2716 20638 2718 20690
rect 2770 20638 2772 20690
rect 2716 20580 2772 20638
rect 2716 20514 2772 20524
rect 3276 20580 3332 20590
rect 3276 20486 3332 20524
rect 2044 20132 2324 20188
rect 1932 17554 1988 17566
rect 1932 17502 1934 17554
rect 1986 17502 1988 17554
rect 1932 16884 1988 17502
rect 1932 16818 1988 16828
rect 1932 11282 1988 11294
rect 1932 11230 1934 11282
rect 1986 11230 1988 11282
rect 1932 10836 1988 11230
rect 1932 10770 1988 10780
rect 2268 9716 2324 20132
rect 2828 17668 2884 17678
rect 2380 17666 2884 17668
rect 2380 17614 2830 17666
rect 2882 17614 2884 17666
rect 2380 17612 2884 17614
rect 2380 17106 2436 17612
rect 2828 17602 2884 17612
rect 2380 17054 2382 17106
rect 2434 17054 2436 17106
rect 2380 17042 2436 17054
rect 2716 17108 2772 17118
rect 2716 16994 2772 17052
rect 3276 17108 3332 17118
rect 3276 17014 3332 17052
rect 2716 16942 2718 16994
rect 2770 16942 2772 16994
rect 2716 16930 2772 16942
rect 2716 12404 2772 12414
rect 2716 12310 2772 12348
rect 3724 12404 3780 29262
rect 4284 29260 4676 29316
rect 4060 28866 4116 28878
rect 4060 28814 4062 28866
rect 4114 28814 4116 28866
rect 4060 28754 4116 28814
rect 4060 28702 4062 28754
rect 4114 28702 4116 28754
rect 4060 28690 4116 28702
rect 4060 28084 4116 28094
rect 4284 28084 4340 29260
rect 4956 29202 5012 29214
rect 4956 29150 4958 29202
rect 5010 29150 5012 29202
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4508 28644 4564 28654
rect 4508 28550 4564 28588
rect 4956 28642 5012 29150
rect 4956 28590 4958 28642
rect 5010 28590 5012 28642
rect 4060 28082 4340 28084
rect 4060 28030 4062 28082
rect 4114 28030 4340 28082
rect 4060 28028 4340 28030
rect 4060 28018 4116 28028
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4956 23492 5012 28590
rect 5068 24388 5124 29932
rect 5180 29540 5236 29550
rect 5180 28756 5236 29484
rect 5404 29202 5460 32284
rect 5516 31556 5572 34188
rect 5740 33460 5796 33470
rect 5852 33460 5908 34860
rect 6188 34916 6244 34926
rect 6188 34822 6244 34860
rect 5740 33458 5908 33460
rect 5740 33406 5742 33458
rect 5794 33406 5908 33458
rect 5740 33404 5908 33406
rect 6188 34468 6244 34478
rect 5740 33394 5796 33404
rect 5852 33236 5908 33246
rect 5628 32338 5684 32350
rect 5628 32286 5630 32338
rect 5682 32286 5684 32338
rect 5628 32228 5684 32286
rect 5628 32162 5684 32172
rect 5740 31556 5796 31566
rect 5516 31554 5796 31556
rect 5516 31502 5742 31554
rect 5794 31502 5796 31554
rect 5516 31500 5796 31502
rect 5404 29150 5406 29202
rect 5458 29150 5460 29202
rect 5404 29138 5460 29150
rect 5516 30996 5572 31006
rect 5516 30882 5572 30940
rect 5516 30830 5518 30882
rect 5570 30830 5572 30882
rect 5180 28690 5236 28700
rect 5516 28084 5572 30830
rect 5628 29764 5684 31500
rect 5740 31490 5796 31500
rect 5740 30212 5796 30222
rect 5852 30212 5908 33180
rect 6076 32900 6132 32910
rect 6076 32786 6132 32844
rect 6076 32734 6078 32786
rect 6130 32734 6132 32786
rect 6076 32722 6132 32734
rect 5964 32564 6020 32574
rect 5964 31778 6020 32508
rect 5964 31726 5966 31778
rect 6018 31726 6020 31778
rect 5964 31668 6020 31726
rect 5964 31602 6020 31612
rect 5740 30210 5908 30212
rect 5740 30158 5742 30210
rect 5794 30158 5908 30210
rect 5740 30156 5908 30158
rect 5740 30146 5796 30156
rect 5628 29698 5684 29708
rect 6076 29652 6132 29662
rect 6188 29652 6244 34412
rect 6300 34356 6356 34366
rect 6300 34262 6356 34300
rect 6412 33572 6468 35644
rect 6636 35026 6692 41132
rect 6860 40964 6916 41244
rect 6860 40898 6916 40908
rect 6860 39844 6916 39854
rect 6748 39732 6804 39742
rect 6748 38834 6804 39676
rect 6860 39506 6916 39788
rect 6860 39454 6862 39506
rect 6914 39454 6916 39506
rect 6860 39442 6916 39454
rect 6748 38782 6750 38834
rect 6802 38782 6804 38834
rect 6748 37268 6804 38782
rect 6972 37492 7028 43374
rect 7084 42082 7140 42094
rect 7084 42030 7086 42082
rect 7138 42030 7140 42082
rect 7084 41860 7140 42030
rect 7196 41860 7252 45052
rect 7308 43316 7364 45612
rect 7420 45666 7476 46508
rect 7420 45614 7422 45666
rect 7474 45614 7476 45666
rect 7420 45556 7476 45614
rect 7420 45490 7476 45500
rect 7532 46562 7588 46574
rect 7532 46510 7534 46562
rect 7586 46510 7588 46562
rect 7532 45332 7588 46510
rect 7532 45266 7588 45276
rect 7532 45108 7588 45118
rect 7532 45014 7588 45052
rect 7532 44772 7588 44782
rect 7532 44324 7588 44716
rect 7756 44772 7812 47404
rect 7868 47234 7924 47246
rect 7868 47182 7870 47234
rect 7922 47182 7924 47234
rect 7868 45668 7924 47182
rect 7980 46786 8036 47404
rect 7980 46734 7982 46786
rect 8034 46734 8036 46786
rect 8092 47348 8148 47358
rect 8092 46900 8148 47292
rect 8092 46768 8148 46844
rect 7980 46722 8036 46734
rect 8092 46452 8148 46462
rect 8092 46358 8148 46396
rect 7980 46004 8036 46014
rect 7980 45890 8036 45948
rect 7980 45838 7982 45890
rect 8034 45838 8036 45890
rect 7980 45826 8036 45838
rect 7868 45602 7924 45612
rect 8204 45220 8260 49196
rect 8316 49028 8372 49038
rect 8316 47570 8372 48972
rect 8316 47518 8318 47570
rect 8370 47518 8372 47570
rect 8316 47506 8372 47518
rect 8428 47460 8484 51212
rect 8428 47394 8484 47404
rect 8540 46116 8596 51324
rect 9884 51378 10052 51380
rect 9884 51326 9998 51378
rect 10050 51326 10052 51378
rect 9884 51324 10052 51326
rect 8876 51268 8932 51278
rect 8876 50596 8932 51212
rect 9660 50932 9716 50942
rect 9660 50818 9716 50876
rect 9660 50766 9662 50818
rect 9714 50766 9716 50818
rect 9660 50754 9716 50766
rect 8876 50540 9044 50596
rect 8988 50484 9044 50540
rect 9100 50484 9156 50494
rect 8988 50482 9156 50484
rect 8988 50430 9102 50482
rect 9154 50430 9156 50482
rect 8988 50428 9156 50430
rect 8652 50370 8708 50382
rect 8652 50318 8654 50370
rect 8706 50318 8708 50370
rect 8652 50260 8708 50318
rect 8652 50194 8708 50204
rect 8652 49810 8708 49822
rect 8652 49758 8654 49810
rect 8706 49758 8708 49810
rect 8652 49700 8708 49758
rect 8652 49476 8708 49644
rect 9100 49700 9156 50428
rect 9436 50372 9492 50382
rect 9100 49634 9156 49644
rect 9324 49924 9380 49934
rect 8652 49410 8708 49420
rect 8988 49140 9044 49150
rect 8988 49046 9044 49084
rect 8652 48354 8708 48366
rect 8652 48302 8654 48354
rect 8706 48302 8708 48354
rect 8652 48244 8708 48302
rect 8652 48178 8708 48188
rect 8988 48242 9044 48254
rect 8988 48190 8990 48242
rect 9042 48190 9044 48242
rect 8764 48132 8820 48142
rect 8764 47460 8820 48076
rect 8428 45892 8484 45902
rect 8428 45798 8484 45836
rect 8204 45088 8260 45164
rect 8428 45106 8484 45118
rect 8428 45054 8430 45106
rect 8482 45054 8484 45106
rect 7756 44706 7812 44716
rect 8204 44772 8260 44782
rect 7980 44436 8036 44446
rect 7532 44322 7812 44324
rect 7532 44270 7534 44322
rect 7586 44270 7812 44322
rect 7532 44268 7812 44270
rect 7532 44258 7588 44268
rect 7532 44100 7588 44110
rect 7420 43540 7476 43550
rect 7420 43446 7476 43484
rect 7308 43260 7476 43316
rect 7308 42644 7364 42654
rect 7308 42194 7364 42588
rect 7308 42142 7310 42194
rect 7362 42142 7364 42194
rect 7308 42130 7364 42142
rect 7420 42084 7476 43260
rect 7420 41990 7476 42028
rect 7532 42754 7588 44044
rect 7532 42702 7534 42754
rect 7586 42702 7588 42754
rect 7196 41804 7476 41860
rect 7084 41794 7140 41804
rect 7308 41188 7364 41198
rect 7308 41074 7364 41132
rect 7308 41022 7310 41074
rect 7362 41022 7364 41074
rect 7308 41010 7364 41022
rect 7084 40516 7140 40526
rect 7084 40422 7140 40460
rect 7196 40292 7252 40302
rect 7196 40198 7252 40236
rect 7308 40180 7364 40190
rect 7308 40086 7364 40124
rect 7420 39956 7476 41804
rect 7532 41186 7588 42702
rect 7532 41134 7534 41186
rect 7586 41134 7588 41186
rect 7532 41076 7588 41134
rect 7644 43988 7700 43998
rect 7756 43988 7812 44268
rect 7868 43988 7924 43998
rect 7756 43932 7868 43988
rect 7644 43650 7700 43932
rect 7868 43922 7924 43932
rect 7644 43598 7646 43650
rect 7698 43598 7700 43650
rect 7644 41188 7700 43598
rect 7868 43762 7924 43774
rect 7868 43710 7870 43762
rect 7922 43710 7924 43762
rect 7868 43540 7924 43710
rect 7980 43650 8036 44380
rect 8092 44210 8148 44222
rect 8092 44158 8094 44210
rect 8146 44158 8148 44210
rect 8092 43876 8148 44158
rect 8092 43810 8148 43820
rect 7980 43598 7982 43650
rect 8034 43598 8036 43650
rect 7980 43586 8036 43598
rect 8092 43652 8148 43662
rect 7868 43474 7924 43484
rect 7756 43428 7812 43438
rect 7756 42642 7812 43372
rect 7756 42590 7758 42642
rect 7810 42590 7812 42642
rect 7756 42308 7812 42590
rect 7756 42242 7812 42252
rect 7644 41122 7700 41132
rect 7756 42084 7812 42094
rect 7532 41010 7588 41020
rect 7756 40964 7812 42028
rect 7980 41300 8036 41310
rect 7980 41206 8036 41244
rect 7196 39900 7476 39956
rect 7644 40908 7812 40964
rect 7084 39620 7140 39630
rect 7084 39060 7140 39564
rect 7084 38994 7140 39004
rect 7084 38052 7140 38062
rect 7084 37958 7140 37996
rect 7196 37604 7252 39900
rect 7532 39842 7588 39854
rect 7532 39790 7534 39842
rect 7586 39790 7588 39842
rect 7532 39730 7588 39790
rect 7532 39678 7534 39730
rect 7586 39678 7588 39730
rect 7532 39666 7588 39678
rect 7420 38834 7476 38846
rect 7420 38782 7422 38834
rect 7474 38782 7476 38834
rect 7420 38612 7476 38782
rect 7644 38668 7700 40908
rect 8092 39956 8148 43596
rect 8204 42196 8260 44716
rect 8428 44660 8484 45054
rect 8540 44884 8596 46060
rect 8652 47458 8820 47460
rect 8652 47406 8766 47458
rect 8818 47406 8820 47458
rect 8652 47404 8820 47406
rect 8652 45892 8708 47404
rect 8764 47394 8820 47404
rect 8876 47684 8932 47694
rect 8876 47068 8932 47628
rect 8988 47348 9044 48190
rect 9212 47684 9268 47694
rect 9212 47570 9268 47628
rect 9212 47518 9214 47570
rect 9266 47518 9268 47570
rect 9212 47506 9268 47518
rect 8988 47216 9044 47292
rect 9212 47348 9268 47358
rect 8764 47012 8932 47068
rect 8764 46786 8820 47012
rect 8764 46734 8766 46786
rect 8818 46734 8820 46786
rect 8764 46722 8820 46734
rect 8876 46900 8932 46910
rect 8876 46004 8932 46844
rect 8652 45826 8708 45836
rect 8764 45948 8932 46004
rect 9100 46674 9156 46686
rect 9100 46622 9102 46674
rect 9154 46622 9156 46674
rect 8764 45780 8820 45948
rect 8988 45892 9044 45902
rect 8988 45798 9044 45836
rect 8764 45724 8932 45780
rect 8652 45668 8708 45678
rect 8708 45612 8820 45668
rect 8652 45602 8708 45612
rect 8652 45108 8708 45118
rect 8652 45014 8708 45052
rect 8540 44828 8708 44884
rect 8428 44594 8484 44604
rect 8428 44324 8484 44334
rect 8428 44230 8484 44268
rect 8540 43652 8596 43662
rect 8540 43558 8596 43596
rect 8316 43428 8372 43438
rect 8316 42532 8372 43372
rect 8316 42466 8372 42476
rect 8428 43316 8484 43326
rect 8428 42308 8484 43260
rect 8540 42532 8596 42542
rect 8540 42438 8596 42476
rect 8428 42252 8596 42308
rect 8204 42084 8260 42140
rect 8316 42084 8372 42094
rect 8204 42082 8372 42084
rect 8204 42030 8318 42082
rect 8370 42030 8372 42082
rect 8204 42028 8372 42030
rect 8316 42018 8372 42028
rect 8428 41524 8484 41534
rect 8428 41186 8484 41468
rect 8428 41134 8430 41186
rect 8482 41134 8484 41186
rect 8428 40740 8484 41134
rect 8428 40674 8484 40684
rect 8540 40628 8596 42252
rect 8652 42194 8708 44828
rect 8764 42868 8820 45612
rect 8876 45218 8932 45724
rect 8876 45166 8878 45218
rect 8930 45166 8932 45218
rect 8876 45154 8932 45166
rect 9100 45108 9156 46622
rect 9212 45444 9268 47292
rect 9212 45378 9268 45388
rect 9212 45108 9268 45118
rect 9100 45052 9212 45108
rect 9212 45042 9268 45052
rect 8988 44996 9044 45006
rect 8988 44994 9156 44996
rect 8988 44942 8990 44994
rect 9042 44942 9156 44994
rect 8988 44940 9156 44942
rect 8988 44930 9044 44940
rect 8988 44212 9044 44222
rect 8988 43876 9044 44156
rect 8988 43810 9044 43820
rect 8988 43428 9044 43438
rect 8988 43334 9044 43372
rect 8988 42868 9044 42878
rect 8764 42866 9044 42868
rect 8764 42814 8990 42866
rect 9042 42814 9044 42866
rect 8764 42812 9044 42814
rect 8652 42142 8654 42194
rect 8706 42142 8708 42194
rect 8652 42130 8708 42142
rect 8988 41860 9044 42812
rect 8988 41794 9044 41804
rect 9100 41188 9156 44940
rect 9212 44322 9268 44334
rect 9212 44270 9214 44322
rect 9266 44270 9268 44322
rect 9212 44100 9268 44270
rect 9212 44034 9268 44044
rect 9212 43428 9268 43438
rect 9212 41300 9268 43372
rect 9324 42084 9380 49868
rect 9436 49252 9492 50316
rect 9772 50036 9828 50046
rect 9436 49026 9492 49196
rect 9436 48974 9438 49026
rect 9490 48974 9492 49026
rect 9436 48962 9492 48974
rect 9548 49700 9604 49710
rect 9436 47460 9492 47470
rect 9436 47366 9492 47404
rect 9548 47124 9604 49644
rect 9772 48914 9828 49980
rect 9772 48862 9774 48914
rect 9826 48862 9828 48914
rect 9772 48850 9828 48862
rect 9548 45890 9604 47068
rect 9772 48356 9828 48366
rect 9660 46900 9716 46910
rect 9660 46806 9716 46844
rect 9772 46898 9828 48300
rect 9884 47684 9940 51324
rect 9996 51314 10052 51324
rect 10220 51378 10276 51390
rect 10220 51326 10222 51378
rect 10274 51326 10276 51378
rect 10108 51268 10164 51278
rect 10108 51174 10164 51212
rect 10220 50932 10276 51326
rect 9996 50876 10276 50932
rect 9996 50818 10052 50876
rect 9996 50766 9998 50818
rect 10050 50766 10052 50818
rect 9996 50754 10052 50766
rect 9996 50596 10052 50606
rect 9996 50594 10164 50596
rect 9996 50542 9998 50594
rect 10050 50542 10164 50594
rect 9996 50540 10164 50542
rect 9996 50530 10052 50540
rect 10108 50484 10164 50540
rect 10332 50428 10388 52782
rect 10444 51380 10500 53788
rect 10444 51286 10500 51324
rect 10556 54068 10612 54078
rect 10556 51268 10612 54012
rect 10780 53844 10836 55244
rect 10780 53778 10836 53788
rect 10668 53730 10724 53742
rect 10668 53678 10670 53730
rect 10722 53678 10724 53730
rect 10668 53170 10724 53678
rect 10668 53118 10670 53170
rect 10722 53118 10724 53170
rect 10668 53106 10724 53118
rect 10892 53170 10948 58156
rect 11116 55972 11172 55982
rect 11116 55878 11172 55916
rect 12124 55970 12180 59200
rect 13356 58436 13412 58446
rect 13244 57764 13300 57774
rect 12796 56756 12852 56766
rect 12796 56082 12852 56700
rect 12796 56030 12798 56082
rect 12850 56030 12852 56082
rect 12796 56018 12852 56030
rect 12124 55918 12126 55970
rect 12178 55918 12180 55970
rect 12124 55906 12180 55918
rect 12908 55412 12964 55422
rect 12964 55356 13076 55412
rect 12908 55318 12964 55356
rect 12124 55188 12180 55198
rect 12124 55094 12180 55132
rect 12572 55188 12628 55198
rect 12572 55186 12964 55188
rect 12572 55134 12574 55186
rect 12626 55134 12964 55186
rect 12572 55132 12964 55134
rect 12572 55122 12628 55132
rect 11004 55076 11060 55086
rect 11004 55074 11172 55076
rect 11004 55022 11006 55074
rect 11058 55022 11172 55074
rect 11004 55020 11172 55022
rect 11004 55010 11060 55020
rect 11004 54628 11060 54638
rect 11004 54514 11060 54572
rect 11004 54462 11006 54514
rect 11058 54462 11060 54514
rect 11004 54450 11060 54462
rect 11116 54404 11172 55020
rect 11116 54338 11172 54348
rect 11676 55074 11732 55086
rect 11676 55022 11678 55074
rect 11730 55022 11732 55074
rect 11116 53508 11172 53518
rect 10892 53118 10894 53170
rect 10946 53118 10948 53170
rect 10892 52276 10948 53118
rect 11004 53506 11172 53508
rect 11004 53454 11118 53506
rect 11170 53454 11172 53506
rect 11004 53452 11172 53454
rect 11004 52946 11060 53452
rect 11116 53442 11172 53452
rect 11228 53506 11284 53518
rect 11228 53454 11230 53506
rect 11282 53454 11284 53506
rect 11004 52894 11006 52946
rect 11058 52894 11060 52946
rect 11004 52276 11060 52894
rect 11228 52948 11284 53454
rect 11340 53508 11396 53518
rect 11340 53506 11620 53508
rect 11340 53454 11342 53506
rect 11394 53454 11620 53506
rect 11340 53452 11620 53454
rect 11340 53442 11396 53452
rect 11228 52882 11284 52892
rect 11004 52220 11396 52276
rect 10892 52210 10948 52220
rect 11116 52052 11172 52062
rect 10780 52050 11172 52052
rect 10780 51998 11118 52050
rect 11170 51998 11172 52050
rect 10780 51996 11172 51998
rect 10668 51268 10724 51278
rect 10556 51266 10724 51268
rect 10556 51214 10670 51266
rect 10722 51214 10724 51266
rect 10556 51212 10724 51214
rect 10668 51202 10724 51212
rect 10108 50418 10164 50428
rect 10220 50372 10388 50428
rect 10444 50820 10500 50830
rect 9996 49700 10052 49710
rect 9996 49606 10052 49644
rect 9996 48356 10052 48366
rect 9996 48262 10052 48300
rect 9884 47618 9940 47628
rect 10108 47796 10164 47806
rect 9996 47572 10052 47582
rect 9996 47478 10052 47516
rect 9772 46846 9774 46898
rect 9826 46846 9828 46898
rect 9772 46676 9828 46846
rect 9548 45838 9550 45890
rect 9602 45838 9604 45890
rect 9548 45826 9604 45838
rect 9660 46620 9828 46676
rect 9884 47460 9940 47470
rect 9660 44548 9716 46620
rect 9884 46564 9940 47404
rect 10108 46788 10164 47740
rect 10220 47124 10276 50372
rect 10332 50036 10388 50046
rect 10444 50036 10500 50764
rect 10388 49980 10500 50036
rect 10332 49140 10388 49980
rect 10780 49924 10836 51996
rect 11116 51986 11172 51996
rect 11228 51938 11284 51950
rect 11228 51886 11230 51938
rect 11282 51886 11284 51938
rect 11228 51828 11284 51886
rect 11228 51762 11284 51772
rect 11340 51716 11396 52220
rect 11452 52162 11508 52174
rect 11452 52110 11454 52162
rect 11506 52110 11508 52162
rect 11452 52052 11508 52110
rect 11452 51986 11508 51996
rect 11340 51604 11396 51660
rect 11228 51548 11396 51604
rect 11004 51380 11060 51390
rect 10332 49074 10388 49084
rect 10444 49868 10836 49924
rect 10892 51378 11060 51380
rect 10892 51326 11006 51378
rect 11058 51326 11060 51378
rect 10892 51324 11060 51326
rect 10892 51266 10948 51324
rect 11004 51314 11060 51324
rect 10892 51214 10894 51266
rect 10946 51214 10948 51266
rect 10444 49698 10500 49868
rect 10444 49646 10446 49698
rect 10498 49646 10500 49698
rect 10332 48356 10388 48366
rect 10332 48262 10388 48300
rect 10332 47348 10388 47358
rect 10332 47254 10388 47292
rect 10220 47068 10388 47124
rect 10220 46788 10276 46798
rect 10108 46786 10276 46788
rect 10108 46734 10222 46786
rect 10274 46734 10276 46786
rect 10108 46732 10276 46734
rect 9772 46508 9940 46564
rect 9996 46674 10052 46686
rect 9996 46622 9998 46674
rect 10050 46622 10052 46674
rect 9772 45780 9828 46508
rect 9996 46340 10052 46622
rect 9996 46274 10052 46284
rect 9884 46004 9940 46014
rect 9884 46002 10052 46004
rect 9884 45950 9886 46002
rect 9938 45950 10052 46002
rect 9884 45948 10052 45950
rect 9884 45938 9940 45948
rect 9772 45724 9940 45780
rect 9884 45332 9940 45724
rect 9996 45444 10052 45948
rect 10108 45780 10164 45790
rect 10108 45686 10164 45724
rect 10220 45444 10276 46732
rect 10332 46340 10388 47068
rect 10444 46450 10500 49646
rect 10668 49700 10724 49710
rect 10668 49606 10724 49644
rect 10892 49252 10948 51214
rect 11004 50706 11060 50718
rect 11004 50654 11006 50706
rect 11058 50654 11060 50706
rect 11004 50034 11060 50654
rect 11004 49982 11006 50034
rect 11058 49982 11060 50034
rect 11004 49970 11060 49982
rect 10892 49196 11172 49252
rect 10780 49140 10836 49150
rect 10836 49084 10948 49140
rect 10780 49074 10836 49084
rect 10556 48916 10612 48926
rect 10556 48822 10612 48860
rect 10892 48914 10948 49084
rect 10892 48862 10894 48914
rect 10946 48862 10948 48914
rect 10892 48850 10948 48862
rect 10780 48804 10836 48814
rect 10444 46398 10446 46450
rect 10498 46398 10500 46450
rect 10444 46386 10500 46398
rect 10556 47572 10612 47582
rect 10332 46274 10388 46284
rect 9996 45388 10164 45444
rect 9884 45276 10052 45332
rect 9772 45220 9828 45230
rect 9772 45126 9828 45164
rect 9660 44492 9940 44548
rect 9660 44324 9716 44334
rect 9660 44230 9716 44268
rect 9772 44322 9828 44334
rect 9772 44270 9774 44322
rect 9826 44270 9828 44322
rect 9436 44212 9492 44222
rect 9436 44118 9492 44156
rect 9772 44212 9828 44270
rect 9772 44146 9828 44156
rect 9772 43876 9828 43886
rect 9772 43762 9828 43820
rect 9772 43710 9774 43762
rect 9826 43710 9828 43762
rect 9772 43698 9828 43710
rect 9548 43092 9604 43102
rect 9884 43092 9940 44492
rect 9548 42642 9604 43036
rect 9548 42590 9550 42642
rect 9602 42590 9604 42642
rect 9548 42196 9604 42590
rect 9548 42130 9604 42140
rect 9660 43036 9940 43092
rect 9324 42018 9380 42028
rect 9660 41748 9716 43036
rect 9884 42866 9940 42878
rect 9884 42814 9886 42866
rect 9938 42814 9940 42866
rect 9884 42756 9940 42814
rect 9884 42690 9940 42700
rect 9772 42530 9828 42542
rect 9772 42478 9774 42530
rect 9826 42478 9828 42530
rect 9772 41972 9828 42478
rect 9772 41906 9828 41916
rect 9884 41858 9940 41870
rect 9884 41806 9886 41858
rect 9938 41806 9940 41858
rect 9884 41748 9940 41806
rect 9660 41746 9940 41748
rect 9660 41694 9886 41746
rect 9938 41694 9940 41746
rect 9660 41692 9940 41694
rect 9884 41616 9940 41692
rect 9548 41356 9828 41412
rect 9548 41300 9604 41356
rect 9212 41244 9604 41300
rect 9660 41188 9716 41198
rect 9100 41186 9716 41188
rect 9100 41134 9662 41186
rect 9714 41134 9716 41186
rect 9100 41132 9716 41134
rect 9660 41122 9716 41132
rect 9772 41188 9828 41356
rect 9772 41122 9828 41132
rect 9884 41186 9940 41198
rect 9884 41134 9886 41186
rect 9938 41134 9940 41186
rect 8764 40628 8820 40638
rect 8540 40626 8820 40628
rect 8540 40574 8766 40626
rect 8818 40574 8820 40626
rect 8540 40572 8820 40574
rect 8764 40562 8820 40572
rect 8876 40628 8932 40666
rect 8876 40562 8932 40572
rect 9884 40628 9940 41134
rect 9884 40562 9940 40572
rect 7756 39900 8148 39956
rect 8428 40514 8484 40526
rect 8428 40462 8430 40514
rect 8482 40462 8484 40514
rect 7756 39842 7812 39900
rect 7756 39790 7758 39842
rect 7810 39790 7812 39842
rect 7756 39778 7812 39790
rect 7980 39620 8036 39630
rect 7980 39526 8036 39564
rect 8316 39506 8372 39518
rect 8316 39454 8318 39506
rect 8370 39454 8372 39506
rect 8204 39396 8260 39406
rect 8316 39396 8372 39454
rect 8260 39340 8372 39396
rect 8428 39396 8484 40462
rect 8204 39330 8260 39340
rect 8428 39330 8484 39340
rect 8540 40402 8596 40414
rect 8540 40350 8542 40402
rect 8594 40350 8596 40402
rect 7756 39284 7812 39294
rect 7756 39058 7812 39228
rect 7756 39006 7758 39058
rect 7810 39006 7812 39058
rect 7756 38994 7812 39006
rect 8092 39060 8148 39070
rect 8092 38966 8148 39004
rect 7980 38946 8036 38958
rect 7980 38894 7982 38946
rect 8034 38894 8036 38946
rect 7644 38612 7812 38668
rect 7420 38546 7476 38556
rect 6972 37426 7028 37436
rect 7084 37548 7252 37604
rect 7308 38276 7364 38286
rect 6972 37268 7028 37278
rect 6804 37266 7028 37268
rect 6804 37214 6974 37266
rect 7026 37214 7028 37266
rect 6804 37212 7028 37214
rect 6748 37136 6804 37212
rect 6972 37202 7028 37212
rect 6860 37044 6916 37054
rect 7084 37044 7140 37548
rect 7196 37380 7252 37390
rect 7196 37286 7252 37324
rect 7308 37156 7364 38220
rect 7420 38164 7476 38174
rect 7420 37266 7476 38108
rect 7532 38052 7588 38062
rect 7532 37958 7588 37996
rect 7420 37214 7422 37266
rect 7474 37214 7476 37266
rect 7420 37202 7476 37214
rect 6860 37042 7140 37044
rect 6860 36990 6862 37042
rect 6914 36990 7140 37042
rect 6860 36988 7140 36990
rect 7196 37100 7364 37156
rect 6860 36708 6916 36988
rect 6860 36642 6916 36652
rect 6972 36820 7028 36830
rect 6972 36594 7028 36764
rect 6972 36542 6974 36594
rect 7026 36542 7028 36594
rect 6972 36530 7028 36542
rect 6748 36484 6804 36494
rect 6748 35698 6804 36428
rect 6748 35646 6750 35698
rect 6802 35646 6804 35698
rect 6748 35634 6804 35646
rect 7196 35586 7252 37100
rect 7644 37044 7700 37054
rect 7532 37042 7700 37044
rect 7532 36990 7646 37042
rect 7698 36990 7700 37042
rect 7532 36988 7700 36990
rect 7420 36932 7476 36942
rect 7420 36482 7476 36876
rect 7420 36430 7422 36482
rect 7474 36430 7476 36482
rect 7420 36418 7476 36430
rect 7532 36596 7588 36988
rect 7644 36978 7700 36988
rect 7196 35534 7198 35586
rect 7250 35534 7252 35586
rect 7196 35474 7252 35534
rect 7196 35422 7198 35474
rect 7250 35422 7252 35474
rect 7196 35410 7252 35422
rect 6636 34974 6638 35026
rect 6690 34974 6692 35026
rect 6636 34962 6692 34974
rect 7308 35140 7364 35150
rect 7308 35026 7364 35084
rect 7308 34974 7310 35026
rect 7362 34974 7364 35026
rect 7308 34962 7364 34974
rect 6860 34692 6916 34702
rect 6860 34130 6916 34636
rect 6860 34078 6862 34130
rect 6914 34078 6916 34130
rect 6860 34066 6916 34078
rect 6636 33908 6692 33918
rect 6636 33814 6692 33852
rect 7308 33908 7364 33918
rect 6636 33572 6692 33582
rect 6412 33570 6692 33572
rect 6412 33518 6638 33570
rect 6690 33518 6692 33570
rect 6412 33516 6692 33518
rect 6636 33506 6692 33516
rect 6748 33236 6804 33246
rect 6748 33142 6804 33180
rect 7308 33234 7364 33852
rect 7308 33182 7310 33234
rect 7362 33182 7364 33234
rect 6412 32788 6468 32798
rect 6412 32694 6468 32732
rect 7196 32788 7252 32798
rect 7196 32694 7252 32732
rect 6412 32228 6468 32238
rect 6412 31218 6468 32172
rect 6860 31778 6916 31790
rect 6860 31726 6862 31778
rect 6914 31726 6916 31778
rect 6636 31554 6692 31566
rect 6636 31502 6638 31554
rect 6690 31502 6692 31554
rect 6636 31444 6692 31502
rect 6636 31378 6692 31388
rect 6412 31166 6414 31218
rect 6466 31166 6468 31218
rect 6412 31154 6468 31166
rect 6748 30996 6804 31006
rect 6860 30996 6916 31726
rect 7308 31218 7364 33182
rect 7420 33236 7476 33246
rect 7420 32562 7476 33180
rect 7420 32510 7422 32562
rect 7474 32510 7476 32562
rect 7420 31668 7476 32510
rect 7420 31602 7476 31612
rect 7308 31166 7310 31218
rect 7362 31166 7364 31218
rect 7308 31154 7364 31166
rect 6748 30994 6916 30996
rect 6748 30942 6750 30994
rect 6802 30942 6916 30994
rect 6748 30940 6916 30942
rect 6748 30884 6804 30940
rect 6748 30818 6804 30828
rect 7308 30212 7364 30222
rect 7308 30118 7364 30156
rect 6412 30100 6468 30110
rect 6412 30006 6468 30044
rect 6636 30100 6692 30110
rect 6076 29650 6244 29652
rect 6076 29598 6078 29650
rect 6130 29598 6244 29650
rect 6076 29596 6244 29598
rect 6636 29650 6692 30044
rect 7532 29876 7588 36540
rect 7644 35586 7700 35598
rect 7644 35534 7646 35586
rect 7698 35534 7700 35586
rect 7644 35140 7700 35534
rect 7644 35074 7700 35084
rect 7644 34244 7700 34254
rect 7756 34244 7812 38612
rect 7980 38500 8036 38894
rect 7980 38434 8036 38444
rect 8204 38388 8260 38398
rect 8204 38164 8260 38332
rect 7980 36594 8036 36606
rect 7980 36542 7982 36594
rect 8034 36542 8036 36594
rect 7980 35588 8036 36542
rect 8092 36484 8148 36494
rect 8092 36390 8148 36428
rect 8204 35922 8260 38108
rect 8540 38052 8596 40350
rect 8876 40404 8932 40414
rect 8876 40292 8932 40348
rect 8764 40236 8932 40292
rect 8988 40402 9044 40414
rect 8988 40350 8990 40402
rect 9042 40350 9044 40402
rect 8652 38836 8708 38846
rect 8652 38742 8708 38780
rect 8764 38668 8820 40236
rect 8988 39730 9044 40350
rect 9772 40404 9828 40414
rect 9772 40310 9828 40348
rect 8988 39678 8990 39730
rect 9042 39678 9044 39730
rect 8988 39666 9044 39678
rect 9100 40180 9156 40190
rect 9996 40180 10052 45276
rect 10108 45106 10164 45388
rect 10220 45378 10276 45388
rect 10444 45780 10500 45790
rect 10108 45054 10110 45106
rect 10162 45054 10164 45106
rect 10108 45042 10164 45054
rect 10332 44994 10388 45006
rect 10332 44942 10334 44994
rect 10386 44942 10388 44994
rect 10220 43426 10276 43438
rect 10220 43374 10222 43426
rect 10274 43374 10276 43426
rect 10220 42868 10276 43374
rect 10220 42802 10276 42812
rect 10108 42420 10164 42430
rect 10108 40626 10164 42364
rect 10332 42196 10388 44942
rect 10444 43988 10500 45724
rect 10556 44436 10612 47516
rect 10668 47012 10724 47022
rect 10668 46898 10724 46956
rect 10668 46846 10670 46898
rect 10722 46846 10724 46898
rect 10668 46834 10724 46846
rect 10780 45780 10836 48748
rect 10892 48242 10948 48254
rect 10892 48190 10894 48242
rect 10946 48190 10948 48242
rect 10892 47572 10948 48190
rect 11116 48244 11172 49196
rect 11228 48356 11284 51548
rect 11340 51378 11396 51390
rect 11340 51326 11342 51378
rect 11394 51326 11396 51378
rect 11340 50932 11396 51326
rect 11340 50866 11396 50876
rect 11452 51266 11508 51278
rect 11452 51214 11454 51266
rect 11506 51214 11508 51266
rect 11340 50594 11396 50606
rect 11340 50542 11342 50594
rect 11394 50542 11396 50594
rect 11340 49364 11396 50542
rect 11452 50596 11508 51214
rect 11564 51156 11620 53452
rect 11676 51604 11732 55022
rect 12796 54964 12852 54974
rect 12236 54740 12292 54750
rect 12236 54516 12292 54684
rect 12460 54628 12516 54638
rect 12460 54534 12516 54572
rect 12796 54626 12852 54908
rect 12796 54574 12798 54626
rect 12850 54574 12852 54626
rect 12012 54514 12292 54516
rect 12012 54462 12238 54514
rect 12290 54462 12292 54514
rect 12012 54460 12292 54462
rect 11900 53508 11956 53518
rect 11676 51538 11732 51548
rect 11788 53506 11956 53508
rect 11788 53454 11902 53506
rect 11954 53454 11956 53506
rect 11788 53452 11956 53454
rect 11564 51090 11620 51100
rect 11676 51378 11732 51390
rect 11676 51326 11678 51378
rect 11730 51326 11732 51378
rect 11564 50596 11620 50606
rect 11452 50594 11620 50596
rect 11452 50542 11566 50594
rect 11618 50542 11620 50594
rect 11452 50540 11620 50542
rect 11564 50530 11620 50540
rect 11340 49140 11396 49308
rect 11340 48804 11396 49084
rect 11452 50260 11508 50270
rect 11452 48916 11508 50204
rect 11676 50260 11732 51326
rect 11564 49810 11620 49822
rect 11564 49758 11566 49810
rect 11618 49758 11620 49810
rect 11564 49700 11620 49758
rect 11564 49634 11620 49644
rect 11564 49252 11620 49262
rect 11676 49252 11732 50204
rect 11564 49250 11732 49252
rect 11564 49198 11566 49250
rect 11618 49198 11732 49250
rect 11564 49196 11732 49198
rect 11564 49186 11620 49196
rect 11564 48916 11620 48926
rect 11452 48914 11620 48916
rect 11452 48862 11566 48914
rect 11618 48862 11620 48914
rect 11452 48860 11620 48862
rect 11564 48850 11620 48860
rect 11676 48916 11732 48954
rect 11676 48850 11732 48860
rect 11340 48748 11508 48804
rect 11228 48290 11284 48300
rect 11116 48150 11172 48188
rect 10892 47506 10948 47516
rect 11004 48132 11060 48142
rect 10892 47348 10948 47358
rect 11004 47348 11060 48076
rect 11340 48018 11396 48030
rect 11340 47966 11342 48018
rect 11394 47966 11396 48018
rect 10892 47346 11060 47348
rect 10892 47294 10894 47346
rect 10946 47294 11060 47346
rect 10892 47292 11060 47294
rect 11116 47458 11172 47470
rect 11116 47406 11118 47458
rect 11170 47406 11172 47458
rect 10892 47282 10948 47292
rect 11004 46450 11060 46462
rect 11004 46398 11006 46450
rect 11058 46398 11060 46450
rect 10780 45714 10836 45724
rect 10892 46340 10948 46350
rect 10892 45106 10948 46284
rect 11004 45890 11060 46398
rect 11004 45838 11006 45890
rect 11058 45838 11060 45890
rect 11004 45826 11060 45838
rect 10892 45054 10894 45106
rect 10946 45054 10948 45106
rect 10780 44546 10836 44558
rect 10780 44494 10782 44546
rect 10834 44494 10836 44546
rect 10780 44436 10836 44494
rect 10556 44434 10836 44436
rect 10556 44382 10782 44434
rect 10834 44382 10836 44434
rect 10556 44380 10836 44382
rect 10780 44370 10836 44380
rect 10444 43932 10724 43988
rect 10668 43764 10724 43932
rect 10780 43764 10836 43774
rect 10668 43762 10836 43764
rect 10668 43710 10782 43762
rect 10834 43710 10836 43762
rect 10668 43708 10836 43710
rect 10780 43698 10836 43708
rect 10780 43428 10836 43438
rect 10668 42754 10724 42766
rect 10668 42702 10670 42754
rect 10722 42702 10724 42754
rect 10444 42644 10500 42654
rect 10444 42550 10500 42588
rect 10332 42140 10500 42196
rect 10332 41972 10388 41982
rect 10332 41878 10388 41916
rect 10108 40574 10110 40626
rect 10162 40574 10164 40626
rect 10108 40562 10164 40574
rect 10220 41746 10276 41758
rect 10444 41748 10500 42140
rect 10668 41972 10724 42702
rect 10668 41906 10724 41916
rect 10780 42420 10836 43372
rect 10892 43092 10948 45054
rect 11116 43708 11172 47406
rect 11340 47236 11396 47966
rect 11340 47170 11396 47180
rect 11228 46676 11284 46686
rect 11228 46582 11284 46620
rect 11452 46450 11508 48748
rect 11676 48692 11732 48702
rect 11676 48466 11732 48636
rect 11676 48414 11678 48466
rect 11730 48414 11732 48466
rect 11676 48402 11732 48414
rect 11676 48244 11732 48254
rect 11676 48150 11732 48188
rect 11788 46676 11844 53452
rect 11900 53442 11956 53452
rect 11900 52946 11956 52958
rect 11900 52894 11902 52946
rect 11954 52894 11956 52946
rect 11900 52388 11956 52894
rect 11900 52322 11956 52332
rect 12012 52500 12068 54460
rect 12236 54450 12292 54460
rect 12684 54402 12740 54414
rect 12684 54350 12686 54402
rect 12738 54350 12740 54402
rect 12572 53508 12628 53518
rect 12572 53414 12628 53452
rect 12684 53058 12740 54350
rect 12684 53006 12686 53058
rect 12738 53006 12740 53058
rect 12684 52994 12740 53006
rect 12572 52948 12628 52958
rect 12572 52854 12628 52892
rect 12012 52444 12292 52500
rect 12012 52386 12068 52444
rect 12012 52334 12014 52386
rect 12066 52334 12068 52386
rect 12012 52322 12068 52334
rect 12124 52276 12180 52286
rect 11900 52164 11956 52174
rect 12124 52164 12180 52220
rect 11900 52162 12180 52164
rect 11900 52110 11902 52162
rect 11954 52110 12180 52162
rect 11900 52108 12180 52110
rect 11900 52098 11956 52108
rect 12124 51940 12180 51950
rect 12236 51940 12292 52444
rect 12796 52388 12852 54574
rect 12908 52724 12964 55132
rect 13020 54292 13076 55356
rect 13132 54964 13188 54974
rect 13132 54740 13188 54908
rect 13132 54674 13188 54684
rect 13132 54514 13188 54526
rect 13132 54462 13134 54514
rect 13186 54462 13188 54514
rect 13132 54404 13188 54462
rect 13132 54338 13188 54348
rect 13020 54226 13076 54236
rect 13020 53506 13076 53518
rect 13020 53454 13022 53506
rect 13074 53454 13076 53506
rect 13020 53060 13076 53454
rect 13020 52994 13076 53004
rect 13132 52948 13188 52958
rect 13132 52854 13188 52892
rect 12908 52668 13188 52724
rect 12796 52322 12852 52332
rect 13020 52388 13076 52398
rect 12684 52276 12740 52286
rect 12684 52164 12740 52220
rect 12908 52276 12964 52286
rect 12908 52182 12964 52220
rect 12796 52164 12852 52174
rect 12684 52162 12852 52164
rect 12684 52110 12798 52162
rect 12850 52110 12852 52162
rect 12684 52108 12852 52110
rect 12796 52098 12852 52108
rect 12572 52052 12628 52062
rect 12572 51958 12628 51996
rect 12180 51884 12292 51940
rect 12348 51940 12404 51950
rect 12124 51874 12180 51884
rect 12348 51846 12404 51884
rect 12236 51492 12292 51502
rect 12236 51398 12292 51436
rect 12124 51380 12180 51390
rect 12124 51286 12180 51324
rect 12460 51380 12516 51390
rect 12460 51286 12516 51324
rect 12796 51380 12852 51390
rect 13020 51380 13076 52332
rect 12796 51378 13076 51380
rect 12796 51326 12798 51378
rect 12850 51326 13076 51378
rect 12796 51324 13076 51326
rect 12796 51314 12852 51324
rect 12236 51268 12292 51278
rect 12124 50932 12180 50942
rect 12012 50708 12068 50718
rect 12012 50594 12068 50652
rect 12012 50542 12014 50594
rect 12066 50542 12068 50594
rect 11900 49922 11956 49934
rect 11900 49870 11902 49922
rect 11954 49870 11956 49922
rect 11900 49476 11956 49870
rect 11900 49410 11956 49420
rect 12012 47572 12068 50542
rect 12124 48132 12180 50876
rect 12236 50594 12292 51212
rect 13020 51156 13076 51166
rect 12236 50542 12238 50594
rect 12290 50542 12292 50594
rect 12236 50530 12292 50542
rect 12460 50818 12516 50830
rect 12460 50766 12462 50818
rect 12514 50766 12516 50818
rect 12348 50148 12404 50158
rect 12348 50034 12404 50092
rect 12348 49982 12350 50034
rect 12402 49982 12404 50034
rect 12348 49970 12404 49982
rect 12124 48038 12180 48076
rect 12236 48802 12292 48814
rect 12236 48750 12238 48802
rect 12290 48750 12292 48802
rect 12012 47478 12068 47516
rect 12236 47348 12292 48750
rect 12460 48804 12516 50766
rect 13020 50708 13076 51100
rect 12908 49812 12964 49822
rect 12908 49718 12964 49756
rect 12908 49140 12964 49150
rect 13020 49140 13076 50652
rect 12908 49138 13076 49140
rect 12908 49086 12910 49138
rect 12962 49086 13076 49138
rect 12908 49084 13076 49086
rect 12908 49074 12964 49084
rect 12460 48738 12516 48748
rect 12796 48468 12852 48478
rect 12236 47282 12292 47292
rect 12460 48244 12516 48254
rect 12460 46788 12516 48188
rect 12684 48242 12740 48254
rect 12684 48190 12686 48242
rect 12738 48190 12740 48242
rect 12460 46722 12516 46732
rect 12572 47346 12628 47358
rect 12572 47294 12574 47346
rect 12626 47294 12628 47346
rect 12572 47124 12628 47294
rect 12684 47236 12740 48190
rect 12796 47570 12852 48412
rect 12908 48356 12964 48366
rect 13132 48356 13188 52668
rect 13244 52612 13300 57708
rect 13356 53396 13412 58380
rect 13692 57876 13748 57886
rect 13468 57316 13524 57326
rect 13468 56532 13524 57260
rect 13692 57316 13748 57820
rect 16380 57876 16436 57886
rect 13692 57250 13748 57260
rect 13916 57428 13972 57438
rect 13468 56466 13524 56476
rect 13692 55972 13748 55982
rect 13692 55970 13860 55972
rect 13692 55918 13694 55970
rect 13746 55918 13860 55970
rect 13692 55916 13860 55918
rect 13692 55906 13748 55916
rect 13692 55074 13748 55086
rect 13692 55022 13694 55074
rect 13746 55022 13748 55074
rect 13692 54180 13748 55022
rect 13804 54404 13860 55916
rect 13804 54338 13860 54348
rect 13916 54738 13972 57372
rect 14924 57428 14980 57438
rect 14812 57204 14868 57214
rect 14924 57204 14980 57372
rect 15036 57204 15092 57214
rect 14924 57148 15036 57204
rect 14140 56196 14196 56206
rect 13916 54686 13918 54738
rect 13970 54686 13972 54738
rect 13692 54114 13748 54124
rect 13804 53620 13860 53630
rect 13804 53526 13860 53564
rect 13356 53340 13524 53396
rect 13356 53172 13412 53182
rect 13356 52946 13412 53116
rect 13356 52894 13358 52946
rect 13410 52894 13412 52946
rect 13356 52882 13412 52894
rect 13468 52724 13524 53340
rect 13692 53060 13748 53070
rect 13916 53060 13972 54686
rect 13692 53058 13972 53060
rect 13692 53006 13694 53058
rect 13746 53006 13972 53058
rect 13692 53004 13972 53006
rect 14028 56084 14084 56094
rect 13692 52994 13748 53004
rect 13244 52388 13300 52556
rect 13244 52322 13300 52332
rect 13356 52668 13524 52724
rect 13356 51156 13412 52668
rect 14028 52050 14084 56028
rect 14140 55860 14196 56140
rect 14588 55970 14644 55982
rect 14588 55918 14590 55970
rect 14642 55918 14644 55970
rect 14140 55794 14196 55804
rect 14364 55858 14420 55870
rect 14364 55806 14366 55858
rect 14418 55806 14420 55858
rect 14140 55076 14196 55086
rect 14140 54516 14196 55020
rect 14140 54450 14196 54460
rect 14252 54290 14308 54302
rect 14252 54238 14254 54290
rect 14306 54238 14308 54290
rect 14140 53508 14196 53518
rect 14140 53414 14196 53452
rect 14028 51998 14030 52050
rect 14082 51998 14084 52050
rect 13692 51938 13748 51950
rect 13692 51886 13694 51938
rect 13746 51886 13748 51938
rect 13692 51828 13748 51886
rect 13356 51090 13412 51100
rect 13580 51772 13692 51828
rect 13468 51044 13524 51054
rect 13244 50932 13300 50942
rect 13244 50034 13300 50876
rect 13244 49982 13246 50034
rect 13298 49982 13300 50034
rect 13244 49970 13300 49982
rect 13356 49812 13412 49822
rect 13244 48356 13300 48366
rect 12908 48262 12964 48300
rect 13020 48300 13244 48356
rect 13020 47796 13076 48300
rect 13244 48224 13300 48300
rect 13020 47730 13076 47740
rect 13132 48130 13188 48142
rect 13132 48078 13134 48130
rect 13186 48078 13188 48130
rect 13132 47684 13188 48078
rect 13356 47796 13412 49756
rect 13356 47730 13412 47740
rect 13132 47618 13188 47628
rect 12796 47518 12798 47570
rect 12850 47518 12852 47570
rect 12796 47506 12852 47518
rect 12796 47236 12852 47246
rect 12684 47180 12796 47236
rect 12796 47142 12852 47180
rect 12124 46676 12180 46686
rect 11788 46620 11956 46676
rect 11564 46564 11620 46574
rect 11564 46470 11620 46508
rect 11452 46398 11454 46450
rect 11506 46398 11508 46450
rect 11340 46116 11396 46126
rect 11340 45890 11396 46060
rect 11340 45838 11342 45890
rect 11394 45838 11396 45890
rect 11228 45780 11284 45790
rect 11228 45686 11284 45724
rect 11340 44772 11396 45838
rect 11340 44706 11396 44716
rect 11452 45218 11508 46398
rect 11900 45332 11956 46620
rect 12124 46582 12180 46620
rect 12460 46562 12516 46574
rect 12460 46510 12462 46562
rect 12514 46510 12516 46562
rect 12460 45780 12516 46510
rect 12460 45714 12516 45724
rect 12124 45668 12180 45678
rect 12124 45666 12292 45668
rect 12124 45614 12126 45666
rect 12178 45614 12292 45666
rect 12124 45612 12292 45614
rect 12124 45602 12180 45612
rect 11900 45276 12068 45332
rect 11452 45166 11454 45218
rect 11506 45166 11508 45218
rect 11452 44324 11508 45166
rect 11676 45106 11732 45118
rect 11676 45054 11678 45106
rect 11730 45054 11732 45106
rect 11452 44258 11508 44268
rect 11564 44546 11620 44558
rect 11564 44494 11566 44546
rect 11618 44494 11620 44546
rect 11340 44100 11396 44110
rect 11340 44098 11508 44100
rect 11340 44046 11342 44098
rect 11394 44046 11508 44098
rect 11340 44044 11508 44046
rect 11340 44034 11396 44044
rect 11116 43652 11284 43708
rect 10892 43026 10948 43036
rect 11004 43540 11060 43550
rect 11004 42868 11060 43484
rect 10780 42194 10836 42364
rect 10780 42142 10782 42194
rect 10834 42142 10836 42194
rect 10220 41694 10222 41746
rect 10274 41694 10276 41746
rect 9100 39508 9156 40124
rect 9660 40124 10052 40180
rect 9548 39620 9604 39630
rect 9548 39526 9604 39564
rect 9100 39414 9156 39452
rect 8876 39394 8932 39406
rect 8876 39342 8878 39394
rect 8930 39342 8932 39394
rect 8876 39284 8932 39342
rect 8876 39218 8932 39228
rect 9100 38722 9156 38734
rect 9100 38670 9102 38722
rect 9154 38670 9156 38722
rect 9100 38668 9156 38670
rect 8764 38612 8932 38668
rect 9100 38612 9268 38668
rect 8540 37986 8596 37996
rect 8764 37266 8820 37278
rect 8764 37214 8766 37266
rect 8818 37214 8820 37266
rect 8316 36484 8372 36494
rect 8316 36370 8372 36428
rect 8316 36318 8318 36370
rect 8370 36318 8372 36370
rect 8316 36306 8372 36318
rect 8204 35870 8206 35922
rect 8258 35870 8260 35922
rect 8204 35858 8260 35870
rect 7700 34188 7812 34244
rect 7868 35474 7924 35486
rect 7868 35422 7870 35474
rect 7922 35422 7924 35474
rect 7868 34802 7924 35422
rect 7868 34750 7870 34802
rect 7922 34750 7924 34802
rect 7644 34150 7700 34188
rect 7756 33908 7812 33918
rect 7644 33122 7700 33134
rect 7644 33070 7646 33122
rect 7698 33070 7700 33122
rect 7644 33012 7700 33070
rect 7644 32946 7700 32956
rect 7756 31890 7812 33852
rect 7756 31838 7758 31890
rect 7810 31838 7812 31890
rect 7756 31826 7812 31838
rect 7868 31444 7924 34750
rect 7980 34130 8036 35532
rect 8428 35812 8484 35822
rect 7980 34078 7982 34130
rect 8034 34078 8036 34130
rect 7980 32900 8036 34078
rect 8092 35140 8148 35150
rect 8092 33458 8148 35084
rect 8204 34804 8260 34814
rect 8204 34710 8260 34748
rect 8428 34354 8484 35756
rect 8652 35700 8708 35710
rect 8652 35606 8708 35644
rect 8764 35698 8820 37214
rect 8764 35646 8766 35698
rect 8818 35646 8820 35698
rect 8876 35812 8932 38612
rect 9100 38500 9156 38510
rect 9100 38050 9156 38444
rect 9100 37998 9102 38050
rect 9154 37998 9156 38050
rect 9100 37986 9156 37998
rect 9212 37940 9268 38612
rect 9212 37874 9268 37884
rect 8988 37380 9044 37390
rect 8988 37286 9044 37324
rect 9212 36596 9268 36606
rect 9212 36502 9268 36540
rect 8876 35680 8932 35756
rect 9548 35812 9604 35822
rect 9100 35700 9156 35710
rect 8764 35588 8820 35646
rect 8764 35522 8820 35532
rect 8876 35476 8932 35486
rect 8764 34804 8820 34814
rect 8876 34804 8932 35420
rect 8764 34802 8932 34804
rect 8764 34750 8766 34802
rect 8818 34750 8932 34802
rect 8764 34748 8932 34750
rect 8988 35140 9044 35150
rect 8764 34738 8820 34748
rect 8428 34302 8430 34354
rect 8482 34302 8484 34354
rect 8428 34290 8484 34302
rect 8876 34018 8932 34030
rect 8876 33966 8878 34018
rect 8930 33966 8932 34018
rect 8876 33908 8932 33966
rect 8876 33842 8932 33852
rect 8092 33406 8094 33458
rect 8146 33406 8148 33458
rect 8092 33394 8148 33406
rect 8876 33346 8932 33358
rect 8876 33294 8878 33346
rect 8930 33294 8932 33346
rect 7980 32844 8148 32900
rect 7868 31378 7924 31388
rect 7980 32676 8036 32686
rect 7644 30994 7700 31006
rect 7644 30942 7646 30994
rect 7698 30942 7700 30994
rect 7644 30884 7700 30942
rect 7644 30818 7700 30828
rect 7980 30210 8036 32620
rect 8092 32340 8148 32844
rect 8876 32788 8932 33294
rect 8988 33234 9044 35084
rect 9100 35138 9156 35644
rect 9100 35086 9102 35138
rect 9154 35086 9156 35138
rect 9100 34804 9156 35086
rect 9324 35140 9380 35150
rect 9324 35026 9380 35084
rect 9324 34974 9326 35026
rect 9378 34974 9380 35026
rect 9324 34962 9380 34974
rect 9100 34738 9156 34748
rect 8988 33182 8990 33234
rect 9042 33182 9044 33234
rect 8988 33170 9044 33182
rect 9436 33572 9492 33582
rect 8652 32732 8932 32788
rect 8652 32676 8708 32732
rect 8428 32620 8708 32676
rect 8428 32562 8484 32620
rect 8428 32510 8430 32562
rect 8482 32510 8484 32562
rect 8428 32498 8484 32510
rect 8540 32452 8596 32462
rect 8540 32358 8596 32396
rect 8092 32284 8484 32340
rect 8428 31666 8484 32284
rect 8652 32228 8708 32620
rect 8652 32162 8708 32172
rect 8764 32562 8820 32574
rect 8764 32510 8766 32562
rect 8818 32510 8820 32562
rect 8764 31892 8820 32510
rect 8988 32564 9044 32574
rect 8988 32470 9044 32508
rect 8764 31826 8820 31836
rect 8428 31614 8430 31666
rect 8482 31614 8484 31666
rect 8428 31602 8484 31614
rect 8764 31666 8820 31678
rect 8764 31614 8766 31666
rect 8818 31614 8820 31666
rect 8764 31556 8820 31614
rect 8540 31444 8596 31454
rect 8092 31332 8148 31342
rect 8092 31218 8148 31276
rect 8092 31166 8094 31218
rect 8146 31166 8148 31218
rect 8092 31154 8148 31166
rect 8540 31218 8596 31388
rect 8540 31166 8542 31218
rect 8594 31166 8596 31218
rect 8540 31154 8596 31166
rect 7980 30158 7982 30210
rect 8034 30158 8036 30210
rect 7980 30100 8036 30158
rect 8316 30212 8372 30222
rect 7980 30034 8036 30044
rect 8204 30098 8260 30110
rect 8204 30046 8206 30098
rect 8258 30046 8260 30098
rect 7532 29810 7588 29820
rect 8204 29876 8260 30046
rect 8204 29810 8260 29820
rect 6636 29598 6638 29650
rect 6690 29598 6692 29650
rect 6076 29540 6132 29596
rect 6076 29474 6132 29484
rect 5740 29314 5796 29326
rect 5740 29262 5742 29314
rect 5794 29262 5796 29314
rect 5740 29202 5796 29262
rect 5740 29150 5742 29202
rect 5794 29150 5796 29202
rect 5740 29138 5796 29150
rect 5516 28018 5572 28028
rect 5068 24322 5124 24332
rect 4956 23426 5012 23436
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 6636 20916 6692 29598
rect 7196 29652 7252 29662
rect 7196 29558 7252 29596
rect 7644 29652 7700 29662
rect 7644 29558 7700 29596
rect 8316 29650 8372 30156
rect 8316 29598 8318 29650
rect 8370 29598 8372 29650
rect 8316 29586 8372 29598
rect 8652 30100 8708 30110
rect 8652 29650 8708 30044
rect 8764 30098 8820 31500
rect 9100 30996 9156 31006
rect 9100 30902 9156 30940
rect 9212 30660 9268 30670
rect 8764 30046 8766 30098
rect 8818 30046 8820 30098
rect 8764 30034 8820 30046
rect 9100 30100 9156 30110
rect 8652 29598 8654 29650
rect 8706 29598 8708 29650
rect 8652 29586 8708 29598
rect 9100 29540 9156 30044
rect 9100 29474 9156 29484
rect 6636 20850 6692 20860
rect 7532 26516 7588 26526
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 7532 17108 7588 26460
rect 7532 17042 7588 17052
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 6972 14308 7028 14318
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 3724 12338 3780 12348
rect 2492 12178 2548 12190
rect 2492 12126 2494 12178
rect 2546 12126 2548 12178
rect 2492 12068 2548 12126
rect 2492 12002 2548 12012
rect 3164 12068 3220 12078
rect 3164 11974 3220 12012
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 2828 11396 2884 11406
rect 2380 11394 2884 11396
rect 2380 11342 2830 11394
rect 2882 11342 2884 11394
rect 2380 11340 2884 11342
rect 2380 10834 2436 11340
rect 2828 11330 2884 11340
rect 2380 10782 2382 10834
rect 2434 10782 2436 10834
rect 2380 10770 2436 10782
rect 2716 10836 2772 10846
rect 2716 10722 2772 10780
rect 3276 10836 3332 10846
rect 3276 10742 3332 10780
rect 2716 10670 2718 10722
rect 2770 10670 2772 10722
rect 2716 10658 2772 10670
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 2380 9716 2436 9726
rect 2268 9714 2436 9716
rect 2268 9662 2382 9714
rect 2434 9662 2436 9714
rect 2268 9660 2436 9662
rect 2380 9650 2436 9660
rect 2716 9716 2772 9726
rect 2716 9622 2772 9660
rect 3276 9716 3332 9726
rect 3276 9622 3332 9660
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 2716 6578 2772 6590
rect 2716 6526 2718 6578
rect 2770 6526 2772 6578
rect 2380 6466 2436 6478
rect 2380 6414 2382 6466
rect 2434 6414 2436 6466
rect 2380 5908 2436 6414
rect 2716 6468 2772 6526
rect 3164 6468 3220 6478
rect 2716 6466 3220 6468
rect 2716 6414 3166 6466
rect 3218 6414 3220 6466
rect 2716 6412 3220 6414
rect 2828 5908 2884 5918
rect 2380 5906 2884 5908
rect 2380 5854 2830 5906
rect 2882 5854 2884 5906
rect 2380 5852 2884 5854
rect 2828 5842 2884 5852
rect 1932 5794 1988 5806
rect 1932 5742 1934 5794
rect 1986 5742 1988 5794
rect 1932 5460 1988 5742
rect 1932 5394 1988 5404
rect 2716 4564 2772 4574
rect 2380 4450 2436 4462
rect 2380 4398 2382 4450
rect 2434 4398 2436 4450
rect 2380 3556 2436 4398
rect 2716 4450 2772 4508
rect 2716 4398 2718 4450
rect 2770 4398 2772 4450
rect 2716 4386 2772 4398
rect 2828 3556 2884 3566
rect 2380 3554 2884 3556
rect 2380 3502 2830 3554
rect 2882 3502 2884 3554
rect 2380 3500 2884 3502
rect 2828 3490 2884 3500
rect 1932 3442 1988 3454
rect 1932 3390 1934 3442
rect 1986 3390 1988 3442
rect 28 1876 84 1886
rect 28 800 84 1820
rect 1932 1876 1988 3390
rect 3164 2660 3220 6412
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 3276 4564 3332 4574
rect 3276 4470 3332 4508
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 6972 3666 7028 14252
rect 9212 4564 9268 30604
rect 9436 30100 9492 33516
rect 9548 33570 9604 35756
rect 9660 35588 9716 40124
rect 9996 39844 10052 39854
rect 9996 39618 10052 39788
rect 9996 39566 9998 39618
rect 10050 39566 10052 39618
rect 9996 39554 10052 39566
rect 10220 39618 10276 41694
rect 10220 39566 10222 39618
rect 10274 39566 10276 39618
rect 10220 39508 10276 39566
rect 10220 39442 10276 39452
rect 10332 41692 10500 41748
rect 10668 41748 10724 41758
rect 10780 41748 10836 42142
rect 10892 42812 11060 42868
rect 11116 43538 11172 43550
rect 11116 43486 11118 43538
rect 11170 43486 11172 43538
rect 10892 42194 10948 42812
rect 10892 42142 10894 42194
rect 10946 42142 10948 42194
rect 10892 42130 10948 42142
rect 11004 42084 11060 42094
rect 11116 42084 11172 43486
rect 11228 42756 11284 43652
rect 11228 42690 11284 42700
rect 11340 42754 11396 42766
rect 11340 42702 11342 42754
rect 11394 42702 11396 42754
rect 11340 42644 11396 42702
rect 11340 42578 11396 42588
rect 11452 42196 11508 44044
rect 11564 42420 11620 44494
rect 11676 44212 11732 45054
rect 12012 45106 12068 45276
rect 12012 45054 12014 45106
rect 12066 45054 12068 45106
rect 11900 44996 11956 45006
rect 11900 44902 11956 44940
rect 11676 44146 11732 44156
rect 11788 44884 11844 44894
rect 11788 44212 11844 44828
rect 12012 44548 12068 45054
rect 12236 44884 12292 45612
rect 12572 45220 12628 47068
rect 13468 46900 13524 50988
rect 13580 50932 13636 51772
rect 13692 51762 13748 51772
rect 13804 51938 13860 51950
rect 13804 51886 13806 51938
rect 13858 51886 13860 51938
rect 13692 51380 13748 51390
rect 13692 51286 13748 51324
rect 13804 51268 13860 51886
rect 13916 51938 13972 51950
rect 13916 51886 13918 51938
rect 13970 51886 13972 51938
rect 13916 51716 13972 51886
rect 13916 51650 13972 51660
rect 14028 51828 14084 51998
rect 13916 51268 13972 51278
rect 13804 51266 13972 51268
rect 13804 51214 13918 51266
rect 13970 51214 13972 51266
rect 13804 51212 13972 51214
rect 13916 51202 13972 51212
rect 13580 50596 13636 50876
rect 13804 50820 13860 50830
rect 13692 50596 13748 50606
rect 13580 50594 13748 50596
rect 13580 50542 13694 50594
rect 13746 50542 13748 50594
rect 13580 50540 13748 50542
rect 13692 48244 13748 50540
rect 13804 50428 13860 50764
rect 13916 50596 13972 50606
rect 14028 50596 14084 51772
rect 14252 50706 14308 54238
rect 14364 53172 14420 55806
rect 14364 53106 14420 53116
rect 14476 53508 14532 53518
rect 14364 52836 14420 52846
rect 14364 52742 14420 52780
rect 14476 52162 14532 53452
rect 14588 53396 14644 55918
rect 14700 55186 14756 55198
rect 14700 55134 14702 55186
rect 14754 55134 14756 55186
rect 14700 54740 14756 55134
rect 14700 54674 14756 54684
rect 14812 55076 14868 57148
rect 15036 57138 15092 57148
rect 14812 54626 14868 55020
rect 14812 54574 14814 54626
rect 14866 54574 14868 54626
rect 14812 54562 14868 54574
rect 14924 56644 14980 56654
rect 14924 55188 14980 56588
rect 16380 56306 16436 57820
rect 16380 56254 16382 56306
rect 16434 56254 16436 56306
rect 15036 55970 15092 55982
rect 15036 55918 15038 55970
rect 15090 55918 15092 55970
rect 15036 55858 15092 55918
rect 15036 55806 15038 55858
rect 15090 55806 15092 55858
rect 15036 55794 15092 55806
rect 15484 55970 15540 55982
rect 15484 55918 15486 55970
rect 15538 55918 15540 55970
rect 14924 54514 14980 55132
rect 14924 54462 14926 54514
rect 14978 54462 14980 54514
rect 14812 54404 14868 54414
rect 14700 53732 14756 53742
rect 14700 53638 14756 53676
rect 14588 53330 14644 53340
rect 14812 53506 14868 54348
rect 14812 53454 14814 53506
rect 14866 53454 14868 53506
rect 14476 52110 14478 52162
rect 14530 52110 14532 52162
rect 14476 52098 14532 52110
rect 14588 53060 14644 53070
rect 14364 51268 14420 51278
rect 14364 51174 14420 51212
rect 14252 50654 14254 50706
rect 14306 50654 14308 50706
rect 14252 50642 14308 50654
rect 14364 50820 14420 50830
rect 13916 50594 14084 50596
rect 13916 50542 13918 50594
rect 13970 50542 14084 50594
rect 13916 50540 14084 50542
rect 13916 50530 13972 50540
rect 14140 50482 14196 50494
rect 14140 50430 14142 50482
rect 14194 50430 14196 50482
rect 13804 50372 13972 50428
rect 13916 49250 13972 50372
rect 14140 49924 14196 50430
rect 14252 50484 14308 50522
rect 14252 50418 14308 50428
rect 14028 49700 14084 49710
rect 14028 49606 14084 49644
rect 14140 49364 14196 49868
rect 14140 49298 14196 49308
rect 13916 49198 13918 49250
rect 13970 49198 13972 49250
rect 13916 49186 13972 49198
rect 14252 49252 14308 49262
rect 14252 49158 14308 49196
rect 14364 49140 14420 50764
rect 14588 50484 14644 53004
rect 14700 52948 14756 52958
rect 14700 52854 14756 52892
rect 14812 52612 14868 53454
rect 14812 52546 14868 52556
rect 14588 50418 14644 50428
rect 14700 52164 14756 52174
rect 14364 49074 14420 49084
rect 14476 49698 14532 49710
rect 14476 49646 14478 49698
rect 14530 49646 14532 49698
rect 13804 49026 13860 49038
rect 13804 48974 13806 49026
rect 13858 48974 13860 49026
rect 13804 48468 13860 48974
rect 14140 49028 14196 49038
rect 14140 48934 14196 48972
rect 13804 48402 13860 48412
rect 14364 48916 14420 48926
rect 13804 48244 13860 48254
rect 13692 48242 13860 48244
rect 13692 48190 13806 48242
rect 13858 48190 13860 48242
rect 13692 48188 13860 48190
rect 13804 48178 13860 48188
rect 14140 48020 14196 48030
rect 14028 47684 14084 47694
rect 14028 47590 14084 47628
rect 14140 47682 14196 47964
rect 14140 47630 14142 47682
rect 14194 47630 14196 47682
rect 14140 47618 14196 47630
rect 14364 47682 14420 48860
rect 14364 47630 14366 47682
rect 14418 47630 14420 47682
rect 14364 47618 14420 47630
rect 14476 47684 14532 49646
rect 14476 47618 14532 47628
rect 14588 49586 14644 49598
rect 14588 49534 14590 49586
rect 14642 49534 14644 49586
rect 14476 47460 14532 47470
rect 14476 47366 14532 47404
rect 13916 46900 13972 46910
rect 13468 46834 13524 46844
rect 13580 46898 13972 46900
rect 13580 46846 13918 46898
rect 13970 46846 13972 46898
rect 13580 46844 13972 46846
rect 13468 46676 13524 46686
rect 13468 46582 13524 46620
rect 12908 46562 12964 46574
rect 12908 46510 12910 46562
rect 12962 46510 12964 46562
rect 12908 46450 12964 46510
rect 12908 46398 12910 46450
rect 12962 46398 12964 46450
rect 12908 46386 12964 46398
rect 13468 46116 13524 46126
rect 12684 46004 12740 46014
rect 12684 45890 12740 45948
rect 12684 45838 12686 45890
rect 12738 45838 12740 45890
rect 12684 45826 12740 45838
rect 12796 45666 12852 45678
rect 12796 45614 12798 45666
rect 12850 45614 12852 45666
rect 12796 45556 12852 45614
rect 12796 45490 12852 45500
rect 13020 45666 13076 45678
rect 13020 45614 13022 45666
rect 13074 45614 13076 45666
rect 13020 45332 13076 45614
rect 13020 45266 13076 45276
rect 13468 45332 13524 46060
rect 13580 45892 13636 46844
rect 13916 46834 13972 46844
rect 14028 46900 14084 46910
rect 13692 46676 13748 46686
rect 14028 46676 14084 46844
rect 13692 46674 13860 46676
rect 13692 46622 13694 46674
rect 13746 46622 13860 46674
rect 13692 46620 13860 46622
rect 13692 46610 13748 46620
rect 13804 46004 13860 46620
rect 14028 46610 14084 46620
rect 14140 46788 14196 46798
rect 14028 46450 14084 46462
rect 14028 46398 14030 46450
rect 14082 46398 14084 46450
rect 14028 46004 14084 46398
rect 13804 45948 13972 46004
rect 13692 45892 13748 45902
rect 13580 45890 13748 45892
rect 13580 45838 13694 45890
rect 13746 45838 13748 45890
rect 13580 45836 13748 45838
rect 13580 45332 13636 45342
rect 13468 45330 13636 45332
rect 13468 45278 13582 45330
rect 13634 45278 13636 45330
rect 13468 45276 13636 45278
rect 12236 44818 12292 44828
rect 12460 45164 12628 45220
rect 13468 45220 13524 45276
rect 13580 45266 13636 45276
rect 13692 45330 13748 45836
rect 13916 45890 13972 45948
rect 14028 45938 14084 45948
rect 13916 45838 13918 45890
rect 13970 45838 13972 45890
rect 13692 45278 13694 45330
rect 13746 45278 13748 45330
rect 13692 45266 13748 45278
rect 13804 45780 13860 45790
rect 12012 44482 12068 44492
rect 12460 44546 12516 45164
rect 13468 45154 13524 45164
rect 13020 45108 13076 45118
rect 12684 45106 13076 45108
rect 12684 45054 13022 45106
rect 13074 45054 13076 45106
rect 12684 45052 13076 45054
rect 12460 44494 12462 44546
rect 12514 44494 12516 44546
rect 12012 44322 12068 44334
rect 12012 44270 12014 44322
rect 12066 44270 12068 44322
rect 11788 44210 11956 44212
rect 11788 44158 11790 44210
rect 11842 44158 11956 44210
rect 11788 44156 11956 44158
rect 11788 44146 11844 44156
rect 11788 43988 11844 43998
rect 11788 43316 11844 43932
rect 11900 43538 11956 44156
rect 12012 43652 12068 44270
rect 12236 44324 12292 44334
rect 12236 44322 12404 44324
rect 12236 44270 12238 44322
rect 12290 44270 12404 44322
rect 12236 44268 12404 44270
rect 12236 44258 12292 44268
rect 12348 43876 12404 44268
rect 12460 43988 12516 44494
rect 12572 44994 12628 45006
rect 12572 44942 12574 44994
rect 12626 44942 12628 44994
rect 12572 44548 12628 44942
rect 12572 44482 12628 44492
rect 12460 43922 12516 43932
rect 12348 43764 12404 43820
rect 12572 43764 12628 43774
rect 12348 43762 12628 43764
rect 12348 43710 12574 43762
rect 12626 43710 12628 43762
rect 12348 43708 12628 43710
rect 12572 43698 12628 43708
rect 12684 43708 12740 45052
rect 13020 45042 13076 45052
rect 13356 45106 13412 45118
rect 13356 45054 13358 45106
rect 13410 45054 13412 45106
rect 12796 44884 12852 44894
rect 12796 44324 12852 44828
rect 12908 44548 12964 44558
rect 13356 44548 13412 45054
rect 12908 44546 13412 44548
rect 12908 44494 12910 44546
rect 12962 44494 13412 44546
rect 12908 44492 13412 44494
rect 13468 44548 13524 44558
rect 12908 44482 12964 44492
rect 12796 44268 13076 44324
rect 12236 43652 12292 43662
rect 12684 43652 12852 43708
rect 12012 43596 12236 43652
rect 11900 43486 11902 43538
rect 11954 43486 11956 43538
rect 11900 43474 11956 43486
rect 12236 43540 12292 43596
rect 12348 43540 12404 43550
rect 12236 43538 12404 43540
rect 12236 43486 12350 43538
rect 12402 43486 12404 43538
rect 12236 43484 12404 43486
rect 12124 43426 12180 43438
rect 12124 43374 12126 43426
rect 12178 43374 12180 43426
rect 12124 43316 12180 43374
rect 11788 43260 12180 43316
rect 11564 42354 11620 42364
rect 11900 42980 11956 42990
rect 11900 42756 11956 42924
rect 12012 42756 12068 42766
rect 11900 42754 12068 42756
rect 11900 42702 12014 42754
rect 12066 42702 12068 42754
rect 11900 42700 12068 42702
rect 11452 42140 11732 42196
rect 11004 42082 11396 42084
rect 11004 42030 11006 42082
rect 11058 42030 11396 42082
rect 11004 42028 11396 42030
rect 11004 42018 11060 42028
rect 10780 41692 11284 41748
rect 9884 39340 10164 39396
rect 9884 38948 9940 39340
rect 10108 39284 10164 39340
rect 10108 39218 10164 39228
rect 9996 39172 10052 39182
rect 9996 39058 10052 39116
rect 9996 39006 9998 39058
rect 10050 39006 10052 39058
rect 9996 38994 10052 39006
rect 9884 38882 9940 38892
rect 10108 38948 10164 38958
rect 10108 38854 10164 38892
rect 9884 38724 9940 38762
rect 9884 37716 9940 38668
rect 9996 38612 10052 38622
rect 9996 38162 10052 38556
rect 9996 38110 9998 38162
rect 10050 38110 10052 38162
rect 9996 38098 10052 38110
rect 10108 37938 10164 37950
rect 10108 37886 10110 37938
rect 10162 37886 10164 37938
rect 10108 37828 10164 37886
rect 10108 37762 10164 37772
rect 9884 37650 9940 37660
rect 9884 37492 9940 37502
rect 9940 37436 10052 37492
rect 9884 37398 9940 37436
rect 9996 36820 10052 37436
rect 9996 36764 10164 36820
rect 9884 36708 9940 36718
rect 9884 36706 10052 36708
rect 9884 36654 9886 36706
rect 9938 36654 10052 36706
rect 9884 36652 10052 36654
rect 9884 36642 9940 36652
rect 9772 36370 9828 36382
rect 9772 36318 9774 36370
rect 9826 36318 9828 36370
rect 9772 35812 9828 36318
rect 9772 35746 9828 35756
rect 9884 36258 9940 36270
rect 9884 36206 9886 36258
rect 9938 36206 9940 36258
rect 9772 35588 9828 35598
rect 9660 35586 9828 35588
rect 9660 35534 9774 35586
rect 9826 35534 9828 35586
rect 9660 35532 9828 35534
rect 9660 35476 9716 35532
rect 9772 35522 9828 35532
rect 9660 35410 9716 35420
rect 9884 35140 9940 36206
rect 9996 35924 10052 36652
rect 9996 35858 10052 35868
rect 10108 35700 10164 36764
rect 9884 35074 9940 35084
rect 9996 35644 10164 35700
rect 10220 36484 10276 36494
rect 9884 34356 9940 34366
rect 9884 34262 9940 34300
rect 9548 33518 9550 33570
rect 9602 33518 9604 33570
rect 9548 32788 9604 33518
rect 9884 33572 9940 33582
rect 9996 33572 10052 35644
rect 10220 35252 10276 36428
rect 10332 35924 10388 41692
rect 10668 41298 10724 41692
rect 10668 41246 10670 41298
rect 10722 41246 10724 41298
rect 10668 41234 10724 41246
rect 10780 41186 10836 41198
rect 10780 41134 10782 41186
rect 10834 41134 10836 41186
rect 10668 41076 10724 41086
rect 10668 40626 10724 41020
rect 10668 40574 10670 40626
rect 10722 40574 10724 40626
rect 10668 40562 10724 40574
rect 10780 40292 10836 41134
rect 11116 41074 11172 41086
rect 11116 41022 11118 41074
rect 11170 41022 11172 41074
rect 11116 40628 11172 41022
rect 11116 40562 11172 40572
rect 11228 40402 11284 41692
rect 11228 40350 11230 40402
rect 11282 40350 11284 40402
rect 11228 40338 11284 40350
rect 10780 40226 10836 40236
rect 11116 40178 11172 40190
rect 11116 40126 11118 40178
rect 11170 40126 11172 40178
rect 11116 39844 11172 40126
rect 11340 39956 11396 42028
rect 11452 41860 11508 41870
rect 11452 41524 11508 41804
rect 11452 41458 11508 41468
rect 11564 40964 11620 40974
rect 11564 40516 11620 40908
rect 11564 40402 11620 40460
rect 11564 40350 11566 40402
rect 11618 40350 11620 40402
rect 11564 40338 11620 40350
rect 11452 40180 11508 40190
rect 11452 40178 11620 40180
rect 11452 40126 11454 40178
rect 11506 40126 11620 40178
rect 11452 40124 11620 40126
rect 11452 40114 11508 40124
rect 11564 40068 11620 40124
rect 11564 40002 11620 40012
rect 11340 39900 11508 39956
rect 11116 39788 11396 39844
rect 10444 39732 10500 39742
rect 10444 39730 11172 39732
rect 10444 39678 10446 39730
rect 10498 39678 11172 39730
rect 10444 39676 11172 39678
rect 10444 39666 10500 39676
rect 11116 39618 11172 39676
rect 11116 39566 11118 39618
rect 11170 39566 11172 39618
rect 11116 39554 11172 39566
rect 11340 39618 11396 39788
rect 11340 39566 11342 39618
rect 11394 39566 11396 39618
rect 11340 39554 11396 39566
rect 10444 39508 10500 39518
rect 10444 39172 10500 39452
rect 10444 37380 10500 39116
rect 10556 39506 10612 39518
rect 10556 39454 10558 39506
rect 10610 39454 10612 39506
rect 10556 39284 10612 39454
rect 10556 38668 10612 39228
rect 10780 39508 10836 39518
rect 10780 38946 10836 39452
rect 11228 39394 11284 39406
rect 11228 39342 11230 39394
rect 11282 39342 11284 39394
rect 11228 39284 11284 39342
rect 11228 39218 11284 39228
rect 10780 38894 10782 38946
rect 10834 38894 10836 38946
rect 10556 38612 10724 38668
rect 10444 36148 10500 37324
rect 10556 37378 10612 37390
rect 10556 37326 10558 37378
rect 10610 37326 10612 37378
rect 10556 37156 10612 37326
rect 10556 37090 10612 37100
rect 10668 36932 10724 38612
rect 10668 36866 10724 36876
rect 10556 36484 10612 36494
rect 10556 36390 10612 36428
rect 10668 36372 10724 36382
rect 10668 36278 10724 36316
rect 10444 36092 10724 36148
rect 10332 35868 10500 35924
rect 10220 34356 10276 35196
rect 10332 35698 10388 35710
rect 10332 35646 10334 35698
rect 10386 35646 10388 35698
rect 10332 35364 10388 35646
rect 10332 34914 10388 35308
rect 10332 34862 10334 34914
rect 10386 34862 10388 34914
rect 10332 34850 10388 34862
rect 10332 34356 10388 34366
rect 10220 34354 10388 34356
rect 10220 34302 10334 34354
rect 10386 34302 10388 34354
rect 10220 34300 10388 34302
rect 10332 34290 10388 34300
rect 9884 33570 10052 33572
rect 9884 33518 9886 33570
rect 9938 33518 10052 33570
rect 9884 33516 10052 33518
rect 9884 33506 9940 33516
rect 9548 32722 9604 32732
rect 9996 32564 10052 32574
rect 9996 32470 10052 32508
rect 9884 32338 9940 32350
rect 9884 32286 9886 32338
rect 9938 32286 9940 32338
rect 9884 32228 9940 32286
rect 9884 32162 9940 32172
rect 10220 32338 10276 32350
rect 10220 32286 10222 32338
rect 10274 32286 10276 32338
rect 9996 31892 10052 31902
rect 9548 31666 9604 31678
rect 9548 31614 9550 31666
rect 9602 31614 9604 31666
rect 9548 31444 9604 31614
rect 9884 31668 9940 31678
rect 9772 31556 9828 31566
rect 9772 31462 9828 31500
rect 9548 31378 9604 31388
rect 9884 31220 9940 31612
rect 9996 31666 10052 31836
rect 10220 31892 10276 32286
rect 10332 32340 10388 32350
rect 10332 32246 10388 32284
rect 10108 31780 10164 31790
rect 10108 31686 10164 31724
rect 9996 31614 9998 31666
rect 10050 31614 10052 31666
rect 9996 31602 10052 31614
rect 9996 31220 10052 31230
rect 9884 31218 10052 31220
rect 9884 31166 9998 31218
rect 10050 31166 10052 31218
rect 9884 31164 10052 31166
rect 9996 31154 10052 31164
rect 9436 30034 9492 30044
rect 9996 30772 10052 30782
rect 9660 29988 9716 29998
rect 9660 29894 9716 29932
rect 9660 29540 9716 29550
rect 9660 28308 9716 29484
rect 9660 28242 9716 28252
rect 9996 24164 10052 30716
rect 10220 30098 10276 31836
rect 10332 30996 10388 31006
rect 10332 30902 10388 30940
rect 10220 30046 10222 30098
rect 10274 30046 10276 30098
rect 10220 30034 10276 30046
rect 10444 29876 10500 35868
rect 10556 34804 10612 34814
rect 10556 34710 10612 34748
rect 10556 33460 10612 33470
rect 10668 33460 10724 36092
rect 10780 35308 10836 38894
rect 11116 38948 11172 38958
rect 11116 38854 11172 38892
rect 11452 38668 11508 39900
rect 11676 39844 11732 42140
rect 11788 41972 11844 41982
rect 11788 41186 11844 41916
rect 11788 41134 11790 41186
rect 11842 41134 11844 41186
rect 11788 41122 11844 41134
rect 11676 39778 11732 39788
rect 11116 38612 11508 38668
rect 11676 39618 11732 39630
rect 11676 39566 11678 39618
rect 11730 39566 11732 39618
rect 11676 38668 11732 39566
rect 11676 38612 11844 38668
rect 10892 37266 10948 37278
rect 10892 37214 10894 37266
rect 10946 37214 10948 37266
rect 10892 36594 10948 37214
rect 10892 36542 10894 36594
rect 10946 36542 10948 36594
rect 10892 36530 10948 36542
rect 11004 35812 11060 35822
rect 11004 35718 11060 35756
rect 10780 35252 11060 35308
rect 10780 34916 10836 34926
rect 10780 34354 10836 34860
rect 10780 34302 10782 34354
rect 10834 34302 10836 34354
rect 10780 34290 10836 34302
rect 10556 33458 10724 33460
rect 10556 33406 10558 33458
rect 10610 33406 10724 33458
rect 10556 33404 10724 33406
rect 11004 33458 11060 35252
rect 11116 34916 11172 38612
rect 11788 38052 11844 38612
rect 11788 37958 11844 37996
rect 11676 37940 11732 37950
rect 11228 37826 11284 37838
rect 11228 37774 11230 37826
rect 11282 37774 11284 37826
rect 11228 37716 11284 37774
rect 11228 37650 11284 37660
rect 11564 37716 11620 37726
rect 11452 35700 11508 35710
rect 11340 35588 11396 35598
rect 11340 35494 11396 35532
rect 11452 35308 11508 35644
rect 11564 35364 11620 37660
rect 11676 36482 11732 37884
rect 11900 36596 11956 42700
rect 12012 42690 12068 42700
rect 12124 42756 12180 42766
rect 12124 42662 12180 42700
rect 12124 42420 12180 42430
rect 12124 42194 12180 42364
rect 12124 42142 12126 42194
rect 12178 42142 12180 42194
rect 12124 42130 12180 42142
rect 12236 42194 12292 43484
rect 12348 43474 12404 43484
rect 12460 43540 12516 43550
rect 12796 43540 12852 43652
rect 12460 43538 12852 43540
rect 12460 43486 12462 43538
rect 12514 43486 12852 43538
rect 12460 43484 12852 43486
rect 12460 43474 12516 43484
rect 12236 42142 12238 42194
rect 12290 42142 12292 42194
rect 12236 42130 12292 42142
rect 12684 42978 12740 42990
rect 12684 42926 12686 42978
rect 12738 42926 12740 42978
rect 12684 42084 12740 42926
rect 12684 42018 12740 42028
rect 13020 41972 13076 44268
rect 13468 44100 13524 44492
rect 13692 44212 13748 44222
rect 13692 44118 13748 44156
rect 13356 43540 13412 43550
rect 13356 43446 13412 43484
rect 13468 43316 13524 44044
rect 13692 43764 13748 43774
rect 13580 43652 13636 43662
rect 13580 43558 13636 43596
rect 13692 43650 13748 43708
rect 13692 43598 13694 43650
rect 13746 43598 13748 43650
rect 13692 43586 13748 43598
rect 13356 43260 13524 43316
rect 13132 42532 13188 42542
rect 13132 42308 13188 42476
rect 13132 42194 13188 42252
rect 13132 42142 13134 42194
rect 13186 42142 13188 42194
rect 13132 42130 13188 42142
rect 13020 41906 13076 41916
rect 12348 41746 12404 41758
rect 12348 41694 12350 41746
rect 12402 41694 12404 41746
rect 12348 41636 12404 41694
rect 12908 41748 12964 41758
rect 13244 41748 13300 41758
rect 12908 41746 13076 41748
rect 12908 41694 12910 41746
rect 12962 41694 13076 41746
rect 12908 41692 13076 41694
rect 12908 41682 12964 41692
rect 12012 41580 12404 41636
rect 12012 41188 12068 41580
rect 12012 41074 12068 41132
rect 12012 41022 12014 41074
rect 12066 41022 12068 41074
rect 12012 40964 12068 41022
rect 12012 40898 12068 40908
rect 12124 41412 12180 41422
rect 12124 41186 12180 41356
rect 12124 41134 12126 41186
rect 12178 41134 12180 41186
rect 12012 38724 12068 38762
rect 12012 38658 12068 38668
rect 11900 36530 11956 36540
rect 11676 36430 11678 36482
rect 11730 36430 11732 36482
rect 11676 36036 11732 36430
rect 11676 35970 11732 35980
rect 12012 36036 12068 36046
rect 11900 35812 11956 35822
rect 11900 35718 11956 35756
rect 11564 35308 11732 35364
rect 11116 34822 11172 34860
rect 11228 35252 11508 35308
rect 11228 34354 11284 35252
rect 11564 35138 11620 35150
rect 11564 35086 11566 35138
rect 11618 35086 11620 35138
rect 11452 35026 11508 35038
rect 11452 34974 11454 35026
rect 11506 34974 11508 35026
rect 11228 34302 11230 34354
rect 11282 34302 11284 34354
rect 11228 33570 11284 34302
rect 11228 33518 11230 33570
rect 11282 33518 11284 33570
rect 11004 33406 11006 33458
rect 11058 33406 11060 33458
rect 10556 33394 10612 33404
rect 11004 33394 11060 33406
rect 11116 33460 11172 33470
rect 11004 32788 11060 32798
rect 10668 32786 11060 32788
rect 10668 32734 11006 32786
rect 11058 32734 11060 32786
rect 10668 32732 11060 32734
rect 10668 31892 10724 32732
rect 11004 32722 11060 32732
rect 10668 31826 10724 31836
rect 10892 32562 10948 32574
rect 10892 32510 10894 32562
rect 10946 32510 10948 32562
rect 10780 31780 10836 31790
rect 10892 31780 10948 32510
rect 11116 32228 11172 33404
rect 11228 32786 11284 33518
rect 11340 34916 11396 34926
rect 11340 33460 11396 34860
rect 11452 34804 11508 34974
rect 11452 34738 11508 34748
rect 11564 34132 11620 35086
rect 11676 34916 11732 35308
rect 11676 34850 11732 34860
rect 11676 34468 11732 34478
rect 11676 34354 11732 34412
rect 11676 34302 11678 34354
rect 11730 34302 11732 34354
rect 11676 34290 11732 34302
rect 12012 34356 12068 35980
rect 12124 35700 12180 41134
rect 12908 40964 12964 40974
rect 12796 40962 12964 40964
rect 12796 40910 12910 40962
rect 12962 40910 12964 40962
rect 12796 40908 12964 40910
rect 12236 40852 12292 40862
rect 12236 40626 12292 40796
rect 12236 40574 12238 40626
rect 12290 40574 12292 40626
rect 12236 40562 12292 40574
rect 12796 40402 12852 40908
rect 12908 40898 12964 40908
rect 12908 40516 12964 40526
rect 12908 40422 12964 40460
rect 12796 40350 12798 40402
rect 12850 40350 12852 40402
rect 12460 40068 12516 40078
rect 12460 39730 12516 40012
rect 12460 39678 12462 39730
rect 12514 39678 12516 39730
rect 12348 39396 12404 39406
rect 12348 39058 12404 39340
rect 12348 39006 12350 39058
rect 12402 39006 12404 39058
rect 12348 38994 12404 39006
rect 12236 38052 12292 38062
rect 12236 37266 12292 37996
rect 12348 37828 12404 37838
rect 12348 37734 12404 37772
rect 12236 37214 12238 37266
rect 12290 37214 12292 37266
rect 12236 37202 12292 37214
rect 12124 35634 12180 35644
rect 12236 36596 12292 36606
rect 12124 34356 12180 34366
rect 12012 34354 12180 34356
rect 12012 34302 12126 34354
rect 12178 34302 12180 34354
rect 12012 34300 12180 34302
rect 11452 33460 11508 33470
rect 11340 33458 11508 33460
rect 11340 33406 11454 33458
rect 11506 33406 11508 33458
rect 11340 33404 11508 33406
rect 11452 33394 11508 33404
rect 11564 33236 11620 34076
rect 11228 32734 11230 32786
rect 11282 32734 11284 32786
rect 11228 32722 11284 32734
rect 11340 33180 11620 33236
rect 11676 33684 11732 33694
rect 10780 31778 10948 31780
rect 10780 31726 10782 31778
rect 10834 31726 10948 31778
rect 10780 31724 10948 31726
rect 11004 32172 11172 32228
rect 10556 31668 10612 31678
rect 10556 31574 10612 31612
rect 10780 31556 10836 31724
rect 10780 31490 10836 31500
rect 10556 30996 10612 31006
rect 10556 30098 10612 30940
rect 10892 30882 10948 30894
rect 10892 30830 10894 30882
rect 10946 30830 10948 30882
rect 10892 30212 10948 30830
rect 10892 30146 10948 30156
rect 10556 30046 10558 30098
rect 10610 30046 10612 30098
rect 10556 29988 10612 30046
rect 11004 29988 11060 32172
rect 11116 32004 11172 32014
rect 11116 31910 11172 31948
rect 11340 31220 11396 33180
rect 11676 33012 11732 33628
rect 11452 32956 11732 33012
rect 11788 33570 11844 33582
rect 11788 33518 11790 33570
rect 11842 33518 11844 33570
rect 11452 31556 11508 32956
rect 11676 32788 11732 32798
rect 11676 32694 11732 32732
rect 11676 31892 11732 31902
rect 11676 31666 11732 31836
rect 11788 31780 11844 33518
rect 11900 33460 11956 33470
rect 12012 33460 12068 34300
rect 12124 34290 12180 34300
rect 11900 33458 12068 33460
rect 11900 33406 11902 33458
rect 11954 33406 12068 33458
rect 11900 33404 12068 33406
rect 11900 33394 11956 33404
rect 12236 33348 12292 36540
rect 12348 36482 12404 36494
rect 12348 36430 12350 36482
rect 12402 36430 12404 36482
rect 12348 35924 12404 36430
rect 12460 36148 12516 39678
rect 12572 39172 12628 39182
rect 12572 39058 12628 39116
rect 12572 39006 12574 39058
rect 12626 39006 12628 39058
rect 12572 38994 12628 39006
rect 12684 38836 12740 38846
rect 12684 38388 12740 38780
rect 12684 38322 12740 38332
rect 12796 38164 12852 40350
rect 12908 39732 12964 39742
rect 12908 39638 12964 39676
rect 12796 38098 12852 38108
rect 12684 37938 12740 37950
rect 12684 37886 12686 37938
rect 12738 37886 12740 37938
rect 12572 37492 12628 37502
rect 12572 36706 12628 37436
rect 12572 36654 12574 36706
rect 12626 36654 12628 36706
rect 12572 36642 12628 36654
rect 12460 36082 12516 36092
rect 12348 35868 12628 35924
rect 12572 35812 12628 35868
rect 12684 35812 12740 37886
rect 13020 37492 13076 41692
rect 13244 41654 13300 41692
rect 13132 41300 13188 41310
rect 13132 40626 13188 41244
rect 13132 40574 13134 40626
rect 13186 40574 13188 40626
rect 13132 40562 13188 40574
rect 13356 40292 13412 43260
rect 13692 42644 13748 42654
rect 13804 42644 13860 45724
rect 13916 45332 13972 45838
rect 14028 45780 14084 45790
rect 14140 45780 14196 46732
rect 14476 46562 14532 46574
rect 14476 46510 14478 46562
rect 14530 46510 14532 46562
rect 14476 46452 14532 46510
rect 14476 46386 14532 46396
rect 14028 45778 14196 45780
rect 14028 45726 14030 45778
rect 14082 45726 14196 45778
rect 14028 45724 14196 45726
rect 14028 45714 14084 45724
rect 14476 45666 14532 45678
rect 14476 45614 14478 45666
rect 14530 45614 14532 45666
rect 14028 45332 14084 45342
rect 13916 45330 14084 45332
rect 13916 45278 14030 45330
rect 14082 45278 14084 45330
rect 13916 45276 14084 45278
rect 14028 45266 14084 45276
rect 14252 45332 14308 45342
rect 14252 45238 14308 45276
rect 14364 45108 14420 45118
rect 14364 45014 14420 45052
rect 14476 44660 14532 45614
rect 14588 45556 14644 49534
rect 14588 45490 14644 45500
rect 14700 48244 14756 52108
rect 14924 52052 14980 54462
rect 15036 55298 15092 55310
rect 15036 55246 15038 55298
rect 15090 55246 15092 55298
rect 15036 53730 15092 55246
rect 15148 55300 15204 55338
rect 15148 55234 15204 55244
rect 15260 55298 15316 55310
rect 15260 55246 15262 55298
rect 15314 55246 15316 55298
rect 15148 55074 15204 55086
rect 15148 55022 15150 55074
rect 15202 55022 15204 55074
rect 15148 54740 15204 55022
rect 15148 54674 15204 54684
rect 15036 53678 15038 53730
rect 15090 53678 15092 53730
rect 15036 53666 15092 53678
rect 15260 53508 15316 55246
rect 15260 53442 15316 53452
rect 15372 54292 15428 54302
rect 15148 53284 15204 53294
rect 15036 53172 15092 53182
rect 15036 52388 15092 53116
rect 15148 52836 15204 53228
rect 15148 52770 15204 52780
rect 15260 52834 15316 52846
rect 15260 52782 15262 52834
rect 15314 52782 15316 52834
rect 15036 52322 15092 52332
rect 15036 52052 15092 52062
rect 14924 52050 15092 52052
rect 14924 51998 15038 52050
rect 15090 51998 15092 52050
rect 14924 51996 15092 51998
rect 14924 51828 14980 51838
rect 14924 51602 14980 51772
rect 14924 51550 14926 51602
rect 14978 51550 14980 51602
rect 14924 51156 14980 51550
rect 14924 51090 14980 51100
rect 15036 50036 15092 51996
rect 15260 51604 15316 52782
rect 15372 52050 15428 54236
rect 15372 51998 15374 52050
rect 15426 51998 15428 52050
rect 15372 51940 15428 51998
rect 15372 51874 15428 51884
rect 15260 51548 15428 51604
rect 15148 51378 15204 51390
rect 15148 51326 15150 51378
rect 15202 51326 15204 51378
rect 15148 50372 15204 51326
rect 15148 50306 15204 50316
rect 15260 50482 15316 50494
rect 15260 50430 15262 50482
rect 15314 50430 15316 50482
rect 14924 49698 14980 49710
rect 14924 49646 14926 49698
rect 14978 49646 14980 49698
rect 14924 49586 14980 49646
rect 14924 49534 14926 49586
rect 14978 49534 14980 49586
rect 14924 49522 14980 49534
rect 15036 49140 15092 49980
rect 14924 49084 15092 49140
rect 14924 48916 14980 49084
rect 15260 49028 15316 50430
rect 15372 50036 15428 51548
rect 15484 50428 15540 55918
rect 15708 55972 15764 55982
rect 15596 55188 15652 55198
rect 15596 54514 15652 55132
rect 15596 54462 15598 54514
rect 15650 54462 15652 54514
rect 15596 54450 15652 54462
rect 15596 53732 15652 53742
rect 15596 53638 15652 53676
rect 15596 52834 15652 52846
rect 15596 52782 15598 52834
rect 15650 52782 15652 52834
rect 15596 52388 15652 52782
rect 15596 52322 15652 52332
rect 15708 51828 15764 55916
rect 15932 55972 15988 55982
rect 15932 55970 16100 55972
rect 15932 55918 15934 55970
rect 15986 55918 16100 55970
rect 15932 55916 16100 55918
rect 15932 55906 15988 55916
rect 15820 55858 15876 55870
rect 15820 55806 15822 55858
rect 15874 55806 15876 55858
rect 15820 53732 15876 55806
rect 15932 54516 15988 54526
rect 15932 54422 15988 54460
rect 15820 53666 15876 53676
rect 16044 53730 16100 55916
rect 16380 55858 16436 56254
rect 17388 56532 17444 56542
rect 16380 55806 16382 55858
rect 16434 55806 16436 55858
rect 16380 55794 16436 55806
rect 16828 55970 16884 55982
rect 16828 55918 16830 55970
rect 16882 55918 16884 55970
rect 16828 55524 16884 55918
rect 16828 55458 16884 55468
rect 16940 55860 16996 55870
rect 16156 55300 16212 55310
rect 16156 54514 16212 55244
rect 16156 54462 16158 54514
rect 16210 54462 16212 54514
rect 16156 53956 16212 54462
rect 16156 53890 16212 53900
rect 16268 55186 16324 55198
rect 16268 55134 16270 55186
rect 16322 55134 16324 55186
rect 16044 53678 16046 53730
rect 16098 53678 16100 53730
rect 16044 52052 16100 53678
rect 16268 53732 16324 55134
rect 16604 55188 16660 55198
rect 16604 55094 16660 55132
rect 16380 55076 16436 55086
rect 16380 54402 16436 55020
rect 16492 54516 16548 54526
rect 16492 54422 16548 54460
rect 16604 54514 16660 54526
rect 16604 54462 16606 54514
rect 16658 54462 16660 54514
rect 16380 54350 16382 54402
rect 16434 54350 16436 54402
rect 16380 53956 16436 54350
rect 16604 54292 16660 54462
rect 16380 53890 16436 53900
rect 16492 54236 16660 54292
rect 16492 53732 16548 54236
rect 16940 53956 16996 55804
rect 17164 55186 17220 55198
rect 17164 55134 17166 55186
rect 17218 55134 17220 55186
rect 17164 54964 17220 55134
rect 17276 55188 17332 55198
rect 17276 55094 17332 55132
rect 17164 54404 17220 54908
rect 17164 54338 17220 54348
rect 17388 54292 17444 56476
rect 17500 56084 17556 56094
rect 17500 55990 17556 56028
rect 17948 55970 18004 55982
rect 17948 55918 17950 55970
rect 18002 55918 18004 55970
rect 17948 55860 18004 55918
rect 18172 55972 18228 59200
rect 21868 58100 21924 58110
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 21868 56420 21924 58044
rect 21868 56354 21924 56364
rect 22652 56196 22708 56206
rect 22652 56194 22820 56196
rect 22652 56142 22654 56194
rect 22706 56142 22820 56194
rect 22652 56140 22820 56142
rect 22652 56130 22708 56140
rect 18508 56084 18564 56094
rect 18508 55990 18564 56028
rect 21644 56084 21700 56094
rect 18172 55906 18228 55916
rect 19068 55972 19124 55982
rect 19068 55878 19124 55916
rect 20188 55970 20244 55982
rect 20188 55918 20190 55970
rect 20242 55918 20244 55970
rect 17948 55794 18004 55804
rect 20188 55858 20244 55918
rect 20188 55806 20190 55858
rect 20242 55806 20244 55858
rect 20188 55794 20244 55806
rect 20748 55970 20804 55982
rect 21308 55972 21364 55982
rect 20748 55918 20750 55970
rect 20802 55918 20804 55970
rect 17836 55636 17892 55646
rect 17500 55074 17556 55086
rect 17500 55022 17502 55074
rect 17554 55022 17556 55074
rect 17500 54516 17556 55022
rect 17724 54516 17780 54526
rect 17500 54514 17780 54516
rect 17500 54462 17726 54514
rect 17778 54462 17780 54514
rect 17500 54460 17780 54462
rect 17724 54450 17780 54460
rect 17836 54516 17892 55580
rect 19852 55636 19908 55646
rect 19516 55524 19572 55534
rect 19180 55298 19236 55310
rect 19180 55246 19182 55298
rect 19234 55246 19236 55298
rect 18172 55186 18228 55198
rect 18172 55134 18174 55186
rect 18226 55134 18228 55186
rect 18172 54852 18228 55134
rect 19180 55188 19236 55246
rect 18172 54786 18228 54796
rect 18284 55074 18340 55086
rect 18284 55022 18286 55074
rect 18338 55022 18340 55074
rect 18172 54516 18228 54526
rect 17836 54514 18228 54516
rect 17836 54462 18174 54514
rect 18226 54462 18228 54514
rect 17836 54460 18228 54462
rect 17388 54226 17444 54236
rect 17836 54068 17892 54460
rect 18172 54450 18228 54460
rect 17948 54292 18004 54302
rect 18172 54292 18228 54302
rect 17948 54198 18004 54236
rect 18060 54236 18172 54292
rect 16268 53676 16548 53732
rect 16828 53900 16996 53956
rect 17724 54012 17892 54068
rect 16268 53508 16324 53676
rect 16268 53442 16324 53452
rect 16604 53618 16660 53630
rect 16604 53566 16606 53618
rect 16658 53566 16660 53618
rect 16380 53396 16436 53406
rect 16156 52836 16212 52846
rect 16156 52742 16212 52780
rect 16380 52164 16436 53340
rect 16492 52836 16548 52846
rect 16604 52836 16660 53566
rect 16716 53506 16772 53518
rect 16716 53454 16718 53506
rect 16770 53454 16772 53506
rect 16716 53060 16772 53454
rect 16828 53172 16884 53900
rect 16940 53732 16996 53742
rect 17612 53732 17668 53742
rect 16940 53730 17668 53732
rect 16940 53678 16942 53730
rect 16994 53678 17614 53730
rect 17666 53678 17668 53730
rect 16940 53676 17668 53678
rect 16940 53666 16996 53676
rect 17612 53666 17668 53676
rect 16828 53106 16884 53116
rect 17052 53508 17108 53518
rect 17724 53508 17780 54012
rect 17836 53844 17892 53854
rect 17836 53730 17892 53788
rect 17836 53678 17838 53730
rect 17890 53678 17892 53730
rect 17836 53666 17892 53678
rect 18060 53730 18116 54236
rect 18172 54226 18228 54236
rect 18060 53678 18062 53730
rect 18114 53678 18116 53730
rect 16716 52994 16772 53004
rect 16940 52836 16996 52846
rect 16604 52834 16996 52836
rect 16604 52782 16942 52834
rect 16994 52782 16996 52834
rect 16604 52780 16996 52782
rect 16492 52742 16548 52780
rect 16380 52098 16436 52108
rect 16604 52612 16660 52622
rect 16268 52052 16324 52062
rect 16044 51996 16212 52052
rect 16156 51828 16212 51996
rect 16268 51958 16324 51996
rect 16492 52052 16548 52090
rect 16492 51986 16548 51996
rect 16380 51938 16436 51950
rect 16380 51886 16382 51938
rect 16434 51886 16436 51938
rect 16156 51772 16324 51828
rect 15708 51762 15764 51772
rect 16156 51380 16212 51390
rect 15708 51378 16212 51380
rect 15708 51326 16158 51378
rect 16210 51326 16212 51378
rect 15708 51324 16212 51326
rect 15708 50706 15764 51324
rect 16156 51314 16212 51324
rect 16268 50932 16324 51772
rect 16380 51716 16436 51886
rect 16380 51650 16436 51660
rect 16492 51828 16548 51838
rect 16380 51490 16436 51502
rect 16380 51438 16382 51490
rect 16434 51438 16436 51490
rect 16380 51380 16436 51438
rect 16492 51490 16548 51772
rect 16492 51438 16494 51490
rect 16546 51438 16548 51490
rect 16492 51426 16548 51438
rect 16380 51314 16436 51324
rect 16492 51266 16548 51278
rect 16492 51214 16494 51266
rect 16546 51214 16548 51266
rect 16492 51044 16548 51214
rect 16492 50978 16548 50988
rect 15708 50654 15710 50706
rect 15762 50654 15764 50706
rect 15708 50642 15764 50654
rect 16044 50706 16100 50718
rect 16044 50654 16046 50706
rect 16098 50654 16100 50706
rect 15484 50372 15764 50428
rect 15372 49970 15428 49980
rect 15484 50260 15540 50270
rect 15484 49812 15540 50204
rect 15484 49718 15540 49756
rect 15708 49810 15764 50372
rect 15708 49758 15710 49810
rect 15762 49758 15764 49810
rect 15708 49588 15764 49758
rect 15260 48972 15652 49028
rect 14924 48354 14980 48860
rect 15148 48804 15204 48814
rect 15148 48802 15428 48804
rect 15148 48750 15150 48802
rect 15202 48750 15428 48802
rect 15148 48748 15428 48750
rect 15148 48738 15204 48748
rect 14924 48302 14926 48354
rect 14978 48302 14980 48354
rect 14924 48290 14980 48302
rect 15148 48580 15204 48590
rect 14812 48244 14868 48254
rect 14700 48242 14868 48244
rect 14700 48190 14814 48242
rect 14866 48190 14868 48242
rect 14700 48188 14868 48190
rect 14476 44594 14532 44604
rect 14140 44436 14196 44446
rect 14140 44100 14196 44380
rect 14140 44006 14196 44044
rect 14252 44324 14308 44334
rect 14028 43540 14084 43550
rect 14028 43446 14084 43484
rect 14140 43428 14196 43438
rect 14140 43334 14196 43372
rect 14252 42980 14308 44268
rect 14588 44098 14644 44110
rect 14588 44046 14590 44098
rect 14642 44046 14644 44098
rect 14588 43764 14644 44046
rect 14364 43708 14644 43764
rect 14364 43316 14420 43708
rect 14588 43540 14644 43550
rect 14364 43250 14420 43260
rect 14476 43538 14644 43540
rect 14476 43486 14590 43538
rect 14642 43486 14644 43538
rect 14476 43484 14644 43486
rect 14140 42978 14308 42980
rect 14140 42926 14254 42978
rect 14306 42926 14308 42978
rect 14140 42924 14308 42926
rect 14028 42868 14084 42878
rect 13916 42644 13972 42654
rect 13804 42588 13916 42644
rect 13692 42550 13748 42588
rect 13916 42550 13972 42588
rect 13692 42420 13748 42430
rect 13580 41972 13636 41982
rect 13580 41188 13636 41916
rect 13580 40516 13636 41132
rect 13692 40626 13748 42364
rect 14028 41970 14084 42812
rect 14140 42196 14196 42924
rect 14252 42914 14308 42924
rect 14140 42130 14196 42140
rect 14252 42754 14308 42766
rect 14252 42702 14254 42754
rect 14306 42702 14308 42754
rect 14252 41972 14308 42702
rect 14364 42756 14420 42766
rect 14364 42082 14420 42700
rect 14476 42530 14532 43484
rect 14588 43474 14644 43484
rect 14476 42478 14478 42530
rect 14530 42478 14532 42530
rect 14476 42466 14532 42478
rect 14588 43316 14644 43326
rect 14588 42308 14644 43260
rect 14588 42242 14644 42252
rect 14364 42030 14366 42082
rect 14418 42030 14420 42082
rect 14364 42018 14420 42030
rect 14028 41918 14030 41970
rect 14082 41918 14084 41970
rect 13916 41748 13972 41758
rect 13916 41654 13972 41692
rect 14028 41412 14084 41918
rect 14028 41346 14084 41356
rect 14140 41916 14308 41972
rect 13692 40574 13694 40626
rect 13746 40574 13748 40626
rect 13692 40562 13748 40574
rect 13916 41298 13972 41310
rect 13916 41246 13918 41298
rect 13970 41246 13972 41298
rect 13580 40450 13636 40460
rect 13916 40404 13972 41246
rect 14028 41186 14084 41198
rect 14028 41134 14030 41186
rect 14082 41134 14084 41186
rect 14028 40964 14084 41134
rect 14028 40898 14084 40908
rect 14140 40740 14196 41916
rect 14252 41748 14308 41758
rect 14252 41654 14308 41692
rect 14364 41412 14420 41422
rect 14252 41188 14308 41198
rect 14252 41094 14308 41132
rect 13916 40338 13972 40348
rect 14028 40684 14196 40740
rect 13356 40226 13412 40236
rect 13580 40180 13636 40190
rect 13468 40178 13636 40180
rect 13468 40126 13582 40178
rect 13634 40126 13636 40178
rect 13468 40124 13636 40126
rect 13020 37426 13076 37436
rect 13356 40068 13412 40078
rect 13356 39058 13412 40012
rect 13468 39620 13524 40124
rect 13580 40114 13636 40124
rect 13916 40178 13972 40190
rect 13916 40126 13918 40178
rect 13970 40126 13972 40178
rect 13692 40068 13748 40078
rect 13692 39844 13748 40012
rect 13916 40068 13972 40126
rect 13916 40002 13972 40012
rect 13692 39788 13972 39844
rect 13468 39554 13524 39564
rect 13580 39732 13636 39742
rect 13356 39006 13358 39058
rect 13410 39006 13412 39058
rect 12908 36484 12964 36494
rect 12908 36390 12964 36428
rect 13020 36148 13076 36158
rect 12908 36036 12964 36046
rect 12796 35812 12852 35822
rect 12572 35810 12852 35812
rect 12572 35758 12798 35810
rect 12850 35758 12852 35810
rect 12572 35756 12852 35758
rect 12460 35698 12516 35710
rect 12460 35646 12462 35698
rect 12514 35646 12516 35698
rect 12460 35476 12516 35646
rect 12460 35410 12516 35420
rect 12572 35028 12628 35038
rect 12572 34934 12628 34972
rect 12796 34804 12852 35756
rect 12908 35252 12964 35980
rect 12908 34914 12964 35196
rect 12908 34862 12910 34914
rect 12962 34862 12964 34914
rect 12908 34850 12964 34862
rect 12796 34738 12852 34748
rect 12572 34692 12628 34702
rect 12572 34356 12628 34636
rect 12572 34224 12628 34300
rect 13020 34020 13076 36092
rect 13244 36036 13300 36046
rect 13020 33926 13076 33964
rect 13132 35812 13188 35822
rect 12124 33292 12292 33348
rect 12908 33348 12964 33358
rect 11900 32562 11956 32574
rect 11900 32510 11902 32562
rect 11954 32510 11956 32562
rect 11900 32452 11956 32510
rect 11900 32004 11956 32396
rect 11900 31938 11956 31948
rect 12124 32004 12180 33292
rect 12908 33254 12964 33292
rect 12236 33124 12292 33134
rect 12236 33030 12292 33068
rect 12796 33124 12852 33134
rect 12796 32562 12852 33068
rect 13132 32786 13188 35756
rect 13244 35810 13300 35980
rect 13244 35758 13246 35810
rect 13298 35758 13300 35810
rect 13244 35746 13300 35758
rect 13356 33572 13412 39006
rect 13468 38948 13524 38958
rect 13468 36148 13524 38892
rect 13580 38164 13636 39676
rect 13916 39618 13972 39788
rect 13916 39566 13918 39618
rect 13970 39566 13972 39618
rect 13916 39554 13972 39566
rect 13692 39506 13748 39518
rect 13692 39454 13694 39506
rect 13746 39454 13748 39506
rect 13692 39396 13748 39454
rect 13692 39330 13748 39340
rect 13580 38098 13636 38108
rect 13692 38834 13748 38846
rect 13692 38782 13694 38834
rect 13746 38782 13748 38834
rect 13692 37940 13748 38782
rect 14028 38052 14084 40684
rect 14364 40404 14420 41356
rect 14252 40348 14420 40404
rect 14252 39842 14308 40348
rect 14588 40292 14644 40302
rect 14252 39790 14254 39842
rect 14306 39790 14308 39842
rect 14252 39778 14308 39790
rect 14364 40290 14644 40292
rect 14364 40238 14590 40290
rect 14642 40238 14644 40290
rect 14364 40236 14644 40238
rect 14252 39620 14308 39630
rect 14252 39526 14308 39564
rect 14252 38948 14308 38958
rect 14252 38854 14308 38892
rect 14140 38724 14196 38734
rect 14364 38668 14420 40236
rect 14588 40226 14644 40236
rect 14476 39956 14532 39966
rect 14476 39394 14532 39900
rect 14476 39342 14478 39394
rect 14530 39342 14532 39394
rect 14476 39330 14532 39342
rect 14588 38948 14644 38958
rect 14588 38854 14644 38892
rect 14140 38612 14420 38668
rect 14700 38668 14756 48188
rect 14812 48178 14868 48188
rect 15036 47684 15092 47694
rect 14812 47236 14868 47246
rect 14924 47236 14980 47246
rect 14868 47234 14980 47236
rect 14868 47182 14926 47234
rect 14978 47182 14980 47234
rect 14868 47180 14980 47182
rect 14812 43540 14868 47180
rect 14924 47170 14980 47180
rect 14924 46564 14980 46574
rect 14924 46470 14980 46508
rect 15036 45780 15092 47628
rect 15148 47236 15204 48524
rect 15260 48468 15316 48478
rect 15260 48374 15316 48412
rect 15260 47796 15316 47806
rect 15260 47458 15316 47740
rect 15260 47406 15262 47458
rect 15314 47406 15316 47458
rect 15260 47394 15316 47406
rect 15148 47142 15204 47180
rect 15260 47124 15316 47134
rect 15260 46900 15316 47068
rect 15148 46844 15316 46900
rect 15148 46002 15204 46844
rect 15372 46788 15428 48748
rect 15148 45950 15150 46002
rect 15202 45950 15204 46002
rect 15148 45938 15204 45950
rect 15260 46732 15428 46788
rect 15484 48802 15540 48814
rect 15484 48750 15486 48802
rect 15538 48750 15540 48802
rect 15036 45714 15092 45724
rect 15148 45220 15204 45230
rect 15148 44100 15204 45164
rect 15260 44882 15316 46732
rect 15372 46564 15428 46574
rect 15372 45892 15428 46508
rect 15484 46340 15540 48750
rect 15484 46274 15540 46284
rect 15596 46676 15652 48972
rect 15708 47124 15764 49532
rect 15820 50036 15876 50046
rect 15820 48916 15876 49980
rect 16044 50034 16100 50654
rect 16156 50596 16212 50634
rect 16156 50530 16212 50540
rect 16044 49982 16046 50034
rect 16098 49982 16100 50034
rect 16044 49970 16100 49982
rect 16156 50372 16212 50382
rect 15932 49924 15988 49934
rect 15932 49830 15988 49868
rect 16156 49028 16212 50316
rect 16156 48934 16212 48972
rect 16268 49364 16324 50876
rect 16492 50036 16548 50046
rect 16380 49812 16436 49822
rect 16380 49718 16436 49756
rect 15820 48242 15876 48860
rect 16268 48914 16324 49308
rect 16268 48862 16270 48914
rect 16322 48862 16324 48914
rect 16268 48850 16324 48862
rect 16044 48804 16100 48814
rect 15820 48190 15822 48242
rect 15874 48190 15876 48242
rect 15820 48178 15876 48190
rect 15932 48354 15988 48366
rect 15932 48302 15934 48354
rect 15986 48302 15988 48354
rect 15708 47058 15764 47068
rect 15596 46116 15652 46620
rect 15596 46050 15652 46060
rect 15708 46788 15764 46798
rect 15708 45892 15764 46732
rect 15932 46788 15988 48302
rect 15932 46722 15988 46732
rect 15820 46564 15876 46574
rect 15820 46470 15876 46508
rect 16044 46228 16100 48748
rect 16492 48132 16548 49980
rect 16604 49588 16660 52556
rect 16940 52388 16996 52780
rect 16940 52322 16996 52332
rect 16828 52052 16884 52062
rect 16716 51940 16772 51950
rect 16716 51846 16772 51884
rect 16828 50372 16884 51996
rect 16940 51380 16996 51390
rect 16940 51286 16996 51324
rect 17052 50428 17108 53452
rect 17388 53452 17780 53508
rect 17164 52612 17220 52622
rect 17164 52052 17220 52556
rect 17388 52052 17444 53452
rect 18060 53396 18116 53678
rect 17612 53340 18116 53396
rect 18172 53730 18228 53742
rect 18172 53678 18174 53730
rect 18226 53678 18228 53730
rect 17500 53284 17556 53294
rect 17500 52724 17556 53228
rect 17612 53170 17668 53340
rect 17612 53118 17614 53170
rect 17666 53118 17668 53170
rect 17612 53106 17668 53118
rect 17500 52274 17556 52668
rect 17500 52222 17502 52274
rect 17554 52222 17556 52274
rect 17500 52210 17556 52222
rect 17724 52500 17780 52510
rect 17388 51996 17556 52052
rect 17164 51986 17220 51996
rect 16828 50306 16884 50316
rect 16940 50372 17108 50428
rect 17388 50484 17444 50522
rect 17388 50418 17444 50428
rect 16716 50036 16772 50046
rect 16716 49942 16772 49980
rect 16940 49922 16996 50372
rect 16940 49870 16942 49922
rect 16994 49870 16996 49922
rect 16940 49812 16996 49870
rect 16940 49746 16996 49756
rect 17388 49924 17444 49934
rect 17052 49588 17108 49598
rect 16604 49532 16772 49588
rect 16604 48356 16660 48366
rect 16604 48262 16660 48300
rect 16492 48076 16660 48132
rect 16044 46162 16100 46172
rect 16268 47570 16324 47582
rect 16268 47518 16270 47570
rect 16322 47518 16324 47570
rect 16156 45892 16212 45902
rect 15708 45836 15876 45892
rect 15372 45826 15428 45836
rect 15820 45780 15876 45836
rect 16156 45798 16212 45836
rect 15708 45666 15764 45678
rect 15708 45614 15710 45666
rect 15762 45614 15764 45666
rect 15260 44830 15262 44882
rect 15314 44830 15316 44882
rect 15260 44818 15316 44830
rect 15372 45556 15428 45566
rect 15260 44548 15316 44558
rect 15260 44454 15316 44492
rect 15148 44034 15204 44044
rect 15372 44322 15428 45500
rect 15708 45444 15764 45614
rect 15708 45378 15764 45388
rect 15596 45332 15652 45342
rect 15596 44996 15652 45276
rect 15596 44902 15652 44940
rect 15372 44270 15374 44322
rect 15426 44270 15428 44322
rect 15148 43652 15204 43662
rect 15148 43558 15204 43596
rect 14812 43474 14868 43484
rect 15036 43538 15092 43550
rect 15036 43486 15038 43538
rect 15090 43486 15092 43538
rect 15036 42868 15092 43486
rect 15260 43540 15316 43550
rect 15260 43446 15316 43484
rect 14812 42812 15092 42868
rect 14812 42644 14868 42812
rect 15372 42756 15428 44270
rect 15596 44322 15652 44334
rect 15596 44270 15598 44322
rect 15650 44270 15652 44322
rect 15596 43764 15652 44270
rect 15708 44212 15764 44222
rect 15708 44118 15764 44156
rect 15596 43316 15652 43708
rect 15820 43652 15876 45724
rect 15932 45666 15988 45678
rect 15932 45614 15934 45666
rect 15986 45614 15988 45666
rect 15932 45556 15988 45614
rect 15932 45490 15988 45500
rect 16044 45666 16100 45678
rect 16044 45614 16046 45666
rect 16098 45614 16100 45666
rect 16044 45332 16100 45614
rect 16044 45266 16100 45276
rect 16044 44994 16100 45006
rect 16044 44942 16046 44994
rect 16098 44942 16100 44994
rect 15820 43586 15876 43596
rect 15932 44882 15988 44894
rect 15932 44830 15934 44882
rect 15986 44830 15988 44882
rect 15820 43428 15876 43438
rect 15596 43250 15652 43260
rect 15708 43426 15876 43428
rect 15708 43374 15822 43426
rect 15874 43374 15876 43426
rect 15708 43372 15876 43374
rect 15708 43204 15764 43372
rect 15820 43362 15876 43372
rect 14812 40964 14868 42588
rect 15036 42700 15428 42756
rect 15484 42980 15540 42990
rect 14812 40292 14868 40908
rect 14812 40226 14868 40236
rect 14924 41076 14980 41086
rect 14924 38948 14980 41020
rect 14700 38612 14868 38668
rect 14028 37958 14084 37996
rect 13692 37874 13748 37884
rect 14364 37938 14420 38612
rect 14700 38500 14756 38510
rect 14364 37886 14366 37938
rect 14418 37886 14420 37938
rect 14252 37268 14308 37278
rect 14252 37174 14308 37212
rect 13468 35698 13524 36092
rect 13468 35646 13470 35698
rect 13522 35646 13524 35698
rect 13468 35634 13524 35646
rect 13804 36482 13860 36494
rect 13804 36430 13806 36482
rect 13858 36430 13860 36482
rect 13692 34802 13748 34814
rect 13692 34750 13694 34802
rect 13746 34750 13748 34802
rect 13468 34132 13524 34142
rect 13692 34132 13748 34750
rect 13804 34468 13860 36430
rect 14028 36372 14084 36382
rect 14028 36278 14084 36316
rect 14252 36370 14308 36382
rect 14252 36318 14254 36370
rect 14306 36318 14308 36370
rect 14028 35700 14084 35710
rect 14028 35606 14084 35644
rect 14028 34916 14084 34926
rect 14028 34802 14084 34860
rect 14028 34750 14030 34802
rect 14082 34750 14084 34802
rect 14028 34738 14084 34750
rect 13804 34402 13860 34412
rect 14028 34356 14084 34366
rect 13524 34076 13748 34132
rect 13804 34132 13860 34142
rect 13468 34038 13524 34076
rect 13804 34038 13860 34076
rect 14028 33684 14084 34300
rect 14252 34020 14308 36318
rect 14364 36372 14420 37886
rect 14476 38162 14532 38174
rect 14476 38110 14478 38162
rect 14530 38110 14532 38162
rect 14476 37378 14532 38110
rect 14700 37490 14756 38444
rect 14700 37438 14702 37490
rect 14754 37438 14756 37490
rect 14700 37426 14756 37438
rect 14476 37326 14478 37378
rect 14530 37326 14532 37378
rect 14476 37314 14532 37326
rect 14476 36372 14532 36382
rect 14364 36370 14532 36372
rect 14364 36318 14478 36370
rect 14530 36318 14532 36370
rect 14364 36316 14532 36318
rect 14476 36260 14532 36316
rect 14476 36204 14756 36260
rect 14364 36148 14420 36158
rect 14420 36092 14644 36148
rect 14364 36082 14420 36092
rect 14588 35922 14644 36092
rect 14588 35870 14590 35922
rect 14642 35870 14644 35922
rect 14588 35858 14644 35870
rect 14700 34580 14756 36204
rect 14812 35700 14868 38612
rect 14924 38050 14980 38892
rect 14924 37998 14926 38050
rect 14978 37998 14980 38050
rect 14924 37986 14980 37998
rect 15036 39730 15092 42700
rect 15372 42532 15428 42542
rect 15484 42532 15540 42924
rect 15372 42530 15540 42532
rect 15372 42478 15374 42530
rect 15426 42478 15540 42530
rect 15372 42476 15540 42478
rect 15372 42466 15428 42476
rect 15148 42420 15204 42430
rect 15148 42194 15204 42364
rect 15148 42142 15150 42194
rect 15202 42142 15204 42194
rect 15148 40516 15204 42142
rect 15148 40450 15204 40460
rect 15372 42308 15428 42318
rect 15372 40402 15428 42252
rect 15596 41858 15652 41870
rect 15596 41806 15598 41858
rect 15650 41806 15652 41858
rect 15596 41076 15652 41806
rect 15708 41860 15764 43148
rect 15820 42644 15876 42654
rect 15820 42550 15876 42588
rect 15932 42532 15988 44830
rect 16044 43988 16100 44942
rect 16100 43932 16212 43988
rect 16044 43922 16100 43932
rect 15932 42466 15988 42476
rect 16044 42530 16100 42542
rect 16044 42478 16046 42530
rect 16098 42478 16100 42530
rect 16044 41972 16100 42478
rect 16156 42532 16212 43932
rect 16268 42868 16324 47518
rect 16492 47458 16548 47470
rect 16492 47406 16494 47458
rect 16546 47406 16548 47458
rect 16380 46900 16436 46910
rect 16380 46806 16436 46844
rect 16492 46898 16548 47406
rect 16604 47236 16660 48076
rect 16604 47170 16660 47180
rect 16492 46846 16494 46898
rect 16546 46846 16548 46898
rect 16492 46834 16548 46846
rect 16716 46788 16772 49532
rect 17052 49586 17220 49588
rect 17052 49534 17054 49586
rect 17106 49534 17220 49586
rect 17052 49532 17220 49534
rect 17052 49522 17108 49532
rect 16940 49140 16996 49216
rect 16828 49084 16940 49140
rect 16828 48692 16884 49084
rect 16940 49074 16996 49084
rect 16940 48916 16996 48926
rect 16940 48914 17108 48916
rect 16940 48862 16942 48914
rect 16994 48862 17108 48914
rect 16940 48860 17108 48862
rect 16940 48850 16996 48860
rect 16828 48636 16996 48692
rect 16828 48356 16884 48366
rect 16828 48262 16884 48300
rect 16940 48130 16996 48636
rect 16940 48078 16942 48130
rect 16994 48078 16996 48130
rect 16940 48066 16996 48078
rect 17052 47458 17108 48860
rect 17164 47684 17220 49532
rect 17388 49026 17444 49868
rect 17388 48974 17390 49026
rect 17442 48974 17444 49026
rect 17388 48692 17444 48974
rect 17388 48626 17444 48636
rect 17164 47618 17220 47628
rect 17276 48244 17332 48254
rect 17052 47406 17054 47458
rect 17106 47406 17108 47458
rect 17052 47394 17108 47406
rect 17164 47460 17220 47470
rect 17164 47366 17220 47404
rect 17052 46900 17108 46910
rect 16828 46788 16884 46798
rect 16716 46732 16828 46788
rect 16604 46674 16660 46686
rect 16604 46622 16606 46674
rect 16658 46622 16660 46674
rect 16604 46340 16660 46622
rect 16604 46274 16660 46284
rect 16828 46452 16884 46732
rect 16716 45778 16772 45790
rect 16716 45726 16718 45778
rect 16770 45726 16772 45778
rect 16716 45220 16772 45726
rect 16716 45154 16772 45164
rect 16492 44994 16548 45006
rect 16492 44942 16494 44994
rect 16546 44942 16548 44994
rect 16492 44882 16548 44942
rect 16492 44830 16494 44882
rect 16546 44830 16548 44882
rect 16492 44212 16548 44830
rect 16716 44996 16772 45006
rect 16604 44212 16660 44222
rect 16492 44210 16660 44212
rect 16492 44158 16606 44210
rect 16658 44158 16660 44210
rect 16492 44156 16660 44158
rect 16604 44146 16660 44156
rect 16716 44210 16772 44940
rect 16716 44158 16718 44210
rect 16770 44158 16772 44210
rect 16380 44098 16436 44110
rect 16380 44046 16382 44098
rect 16434 44046 16436 44098
rect 16380 43538 16436 44046
rect 16716 43988 16772 44158
rect 16716 43922 16772 43932
rect 16716 43652 16772 43662
rect 16716 43558 16772 43596
rect 16380 43486 16382 43538
rect 16434 43486 16436 43538
rect 16380 43474 16436 43486
rect 16492 43538 16548 43550
rect 16492 43486 16494 43538
rect 16546 43486 16548 43538
rect 16380 42980 16436 42990
rect 16492 42980 16548 43486
rect 16380 42978 16548 42980
rect 16380 42926 16382 42978
rect 16434 42926 16548 42978
rect 16380 42924 16548 42926
rect 16380 42914 16436 42924
rect 16268 42802 16324 42812
rect 16156 42466 16212 42476
rect 16268 42530 16324 42542
rect 16268 42478 16270 42530
rect 16322 42478 16324 42530
rect 16268 42308 16324 42478
rect 16268 42242 16324 42252
rect 16492 42532 16548 42542
rect 16492 41972 16548 42476
rect 16604 42196 16660 42206
rect 16604 42102 16660 42140
rect 16100 41916 16212 41972
rect 16044 41878 16100 41916
rect 15708 41794 15764 41804
rect 15596 41010 15652 41020
rect 15372 40350 15374 40402
rect 15426 40350 15428 40402
rect 15372 40338 15428 40350
rect 15484 40962 15540 40974
rect 15484 40910 15486 40962
rect 15538 40910 15540 40962
rect 15148 40292 15204 40302
rect 15148 40198 15204 40236
rect 15036 39678 15038 39730
rect 15090 39678 15092 39730
rect 15036 36484 15092 39678
rect 15484 39284 15540 40910
rect 15932 40964 15988 40974
rect 15932 40962 16100 40964
rect 15932 40910 15934 40962
rect 15986 40910 16100 40962
rect 15932 40908 16100 40910
rect 15932 40898 15988 40908
rect 15820 40404 15876 40414
rect 15820 40310 15876 40348
rect 15932 39508 15988 39518
rect 15484 39218 15540 39228
rect 15596 39394 15652 39406
rect 15596 39342 15598 39394
rect 15650 39342 15652 39394
rect 15260 38722 15316 38734
rect 15260 38670 15262 38722
rect 15314 38670 15316 38722
rect 15036 36418 15092 36428
rect 15148 37828 15204 37838
rect 15148 37266 15204 37772
rect 15148 37214 15150 37266
rect 15202 37214 15204 37266
rect 15036 36148 15092 36158
rect 14812 35634 14868 35644
rect 14924 35698 14980 35710
rect 14924 35646 14926 35698
rect 14978 35646 14980 35698
rect 14924 35028 14980 35646
rect 14924 34914 14980 34972
rect 14924 34862 14926 34914
rect 14978 34862 14980 34914
rect 14924 34850 14980 34862
rect 14700 34514 14756 34524
rect 14924 34356 14980 34366
rect 15036 34356 15092 36092
rect 15148 34802 15204 37214
rect 15260 35364 15316 38670
rect 15372 38164 15428 38174
rect 15372 37266 15428 38108
rect 15596 38052 15652 39342
rect 15708 39060 15764 39070
rect 15708 38668 15764 39004
rect 15708 38612 15876 38668
rect 15596 37986 15652 37996
rect 15708 37828 15764 37838
rect 15372 37214 15374 37266
rect 15426 37214 15428 37266
rect 15372 37202 15428 37214
rect 15596 37826 15764 37828
rect 15596 37774 15710 37826
rect 15762 37774 15764 37826
rect 15596 37772 15764 37774
rect 15596 37492 15652 37772
rect 15708 37762 15764 37772
rect 15820 37716 15876 38612
rect 15820 37650 15876 37660
rect 15596 36482 15652 37436
rect 15596 36430 15598 36482
rect 15650 36430 15652 36482
rect 15596 36418 15652 36430
rect 15708 37042 15764 37054
rect 15708 36990 15710 37042
rect 15762 36990 15764 37042
rect 15484 36372 15540 36382
rect 15484 36278 15540 36316
rect 15708 36372 15764 36990
rect 15708 36306 15764 36316
rect 15596 35588 15652 35626
rect 15596 35522 15652 35532
rect 15260 35298 15316 35308
rect 15596 35364 15652 35374
rect 15148 34750 15150 34802
rect 15202 34750 15204 34802
rect 15148 34738 15204 34750
rect 14476 34354 15092 34356
rect 14476 34302 14926 34354
rect 14978 34302 15092 34354
rect 14476 34300 15092 34302
rect 15596 34356 15652 35308
rect 15708 35028 15764 35038
rect 15708 34934 15764 34972
rect 15820 34804 15876 34814
rect 15820 34710 15876 34748
rect 15708 34356 15764 34366
rect 15596 34300 15708 34356
rect 14252 33954 14308 33964
rect 14364 34132 14420 34142
rect 14140 33906 14196 33918
rect 14140 33854 14142 33906
rect 14194 33854 14196 33906
rect 14140 33796 14196 33854
rect 14140 33730 14196 33740
rect 14028 33618 14084 33628
rect 13356 33506 13412 33516
rect 14364 33458 14420 34076
rect 14364 33406 14366 33458
rect 14418 33406 14420 33458
rect 14364 33394 14420 33406
rect 13804 33348 13860 33358
rect 13132 32734 13134 32786
rect 13186 32734 13188 32786
rect 13132 32722 13188 32734
rect 13692 33234 13748 33246
rect 13692 33182 13694 33234
rect 13746 33182 13748 33234
rect 12796 32510 12798 32562
rect 12850 32510 12852 32562
rect 12572 32452 12628 32462
rect 12572 32358 12628 32396
rect 12124 31938 12180 31948
rect 11900 31780 11956 31790
rect 12460 31780 12516 31790
rect 11788 31778 12516 31780
rect 11788 31726 11902 31778
rect 11954 31726 12462 31778
rect 12514 31726 12516 31778
rect 11788 31724 12516 31726
rect 11900 31714 11956 31724
rect 12460 31714 12516 31724
rect 11676 31614 11678 31666
rect 11730 31614 11732 31666
rect 11676 31602 11732 31614
rect 11452 31490 11508 31500
rect 11452 31220 11508 31230
rect 11340 31218 11508 31220
rect 11340 31166 11454 31218
rect 11506 31166 11508 31218
rect 11340 31164 11508 31166
rect 11452 31154 11508 31164
rect 11116 30884 11172 30894
rect 11116 30790 11172 30828
rect 12012 30884 12068 30894
rect 12012 30790 12068 30828
rect 12796 30548 12852 32510
rect 13580 32564 13636 32574
rect 13692 32564 13748 33182
rect 13804 33234 13860 33292
rect 13804 33182 13806 33234
rect 13858 33182 13860 33234
rect 13804 33170 13860 33182
rect 14028 33124 14084 33134
rect 14028 33030 14084 33068
rect 14140 32788 14196 32798
rect 14140 32694 14196 32732
rect 13580 32562 13748 32564
rect 13580 32510 13582 32562
rect 13634 32510 13748 32562
rect 13580 32508 13748 32510
rect 14028 32562 14084 32574
rect 14028 32510 14030 32562
rect 14082 32510 14084 32562
rect 13580 31780 13636 32508
rect 13580 31714 13636 31724
rect 13020 31556 13076 31566
rect 13020 31332 13076 31500
rect 13020 31266 13076 31276
rect 13580 31554 13636 31566
rect 13580 31502 13582 31554
rect 13634 31502 13636 31554
rect 13356 31108 13412 31118
rect 13356 31106 13524 31108
rect 13356 31054 13358 31106
rect 13410 31054 13524 31106
rect 13356 31052 13524 31054
rect 13356 31042 13412 31052
rect 12796 30482 12852 30492
rect 11452 30212 11508 30222
rect 11452 30098 11508 30156
rect 11900 30212 11956 30222
rect 11900 30118 11956 30156
rect 11452 30046 11454 30098
rect 11506 30046 11508 30098
rect 11452 30034 11508 30046
rect 11564 30100 11620 30110
rect 10556 29922 10612 29932
rect 10668 29932 11060 29988
rect 11116 29988 11172 29998
rect 9996 24098 10052 24108
rect 10108 29820 10500 29876
rect 10108 22708 10164 29820
rect 10444 29428 10500 29438
rect 10444 29334 10500 29372
rect 10332 28084 10388 28094
rect 10332 27990 10388 28028
rect 10108 22642 10164 22652
rect 10668 10836 10724 29932
rect 11116 29894 11172 29932
rect 11452 29428 11508 29438
rect 11452 29334 11508 29372
rect 10892 29314 10948 29326
rect 10892 29262 10894 29314
rect 10946 29262 10948 29314
rect 10892 27076 10948 29262
rect 11340 27860 11396 27870
rect 11340 27766 11396 27804
rect 11340 27412 11396 27422
rect 11004 27076 11060 27086
rect 10892 27074 11060 27076
rect 10892 27022 11006 27074
rect 11058 27022 11060 27074
rect 10892 27020 11060 27022
rect 11004 27010 11060 27020
rect 11340 26850 11396 27356
rect 11564 26908 11620 30044
rect 12908 30100 12964 30110
rect 12908 30006 12964 30044
rect 12348 29988 12404 29998
rect 13468 29988 13524 31052
rect 13580 30996 13636 31502
rect 13580 30930 13636 30940
rect 14028 30996 14084 32510
rect 14252 32562 14308 32574
rect 14252 32510 14254 32562
rect 14306 32510 14308 32562
rect 14252 31892 14308 32510
rect 14476 32452 14532 34300
rect 14924 34290 14980 34300
rect 15708 34262 15764 34300
rect 14588 34130 14644 34142
rect 14588 34078 14590 34130
rect 14642 34078 14644 34130
rect 14588 34020 14644 34078
rect 14588 33954 14644 33964
rect 14252 31826 14308 31836
rect 14364 32396 14532 32452
rect 14812 33684 14868 33694
rect 14812 32674 14868 33628
rect 15932 33572 15988 39452
rect 16044 38612 16100 40908
rect 16156 39732 16212 41916
rect 16492 41186 16548 41916
rect 16492 41134 16494 41186
rect 16546 41134 16548 41186
rect 16492 41122 16548 41134
rect 16604 41748 16660 41758
rect 16828 41748 16884 46396
rect 16940 46676 16996 46686
rect 16940 46340 16996 46620
rect 16940 46274 16996 46284
rect 17052 46114 17108 46844
rect 17052 46062 17054 46114
rect 17106 46062 17108 46114
rect 17052 46050 17108 46062
rect 17052 45892 17108 45902
rect 17052 45798 17108 45836
rect 17164 45778 17220 45790
rect 17164 45726 17166 45778
rect 17218 45726 17220 45778
rect 16940 45108 16996 45118
rect 16940 43764 16996 45052
rect 17164 44882 17220 45726
rect 17164 44830 17166 44882
rect 17218 44830 17220 44882
rect 17164 44818 17220 44830
rect 16940 43698 16996 43708
rect 16940 43540 16996 43550
rect 16940 43446 16996 43484
rect 17052 43426 17108 43438
rect 17052 43374 17054 43426
rect 17106 43374 17108 43426
rect 17052 42978 17108 43374
rect 17052 42926 17054 42978
rect 17106 42926 17108 42978
rect 17052 42914 17108 42926
rect 16940 42868 16996 42878
rect 16940 42774 16996 42812
rect 17276 42308 17332 48188
rect 17500 47684 17556 51996
rect 17724 51602 17780 52444
rect 17724 51550 17726 51602
rect 17778 51550 17780 51602
rect 17612 51380 17668 51390
rect 17612 51286 17668 51324
rect 17724 51156 17780 51550
rect 17612 51100 17780 51156
rect 17612 49924 17668 51100
rect 17612 49858 17668 49868
rect 17724 50594 17780 50606
rect 17724 50542 17726 50594
rect 17778 50542 17780 50594
rect 17724 50372 17780 50542
rect 17836 50428 17892 53340
rect 17948 53172 18004 53182
rect 17948 52500 18004 53116
rect 18172 52612 18228 53678
rect 18284 53620 18340 55022
rect 18396 55076 18452 55086
rect 18396 54290 18452 55020
rect 19068 54738 19124 54750
rect 19068 54686 19070 54738
rect 19122 54686 19124 54738
rect 19068 54628 19124 54686
rect 19068 54562 19124 54572
rect 19180 54404 19236 55132
rect 19404 55076 19460 55086
rect 19404 54982 19460 55020
rect 19068 54348 19236 54404
rect 18396 54238 18398 54290
rect 18450 54238 18452 54290
rect 18396 54226 18452 54238
rect 18620 54292 18676 54302
rect 18620 54198 18676 54236
rect 18844 54290 18900 54302
rect 18844 54238 18846 54290
rect 18898 54238 18900 54290
rect 18844 54068 18900 54238
rect 18844 54002 18900 54012
rect 18284 53554 18340 53564
rect 18844 53620 18900 53630
rect 18844 53526 18900 53564
rect 18956 53506 19012 53518
rect 18956 53454 18958 53506
rect 19010 53454 19012 53506
rect 18396 53172 18452 53182
rect 18396 53078 18452 53116
rect 18956 53060 19012 53454
rect 18732 53004 19012 53060
rect 18172 52546 18228 52556
rect 18284 52722 18340 52734
rect 18284 52670 18286 52722
rect 18338 52670 18340 52722
rect 17948 52164 18004 52444
rect 18284 52386 18340 52670
rect 18508 52724 18564 52734
rect 18284 52334 18286 52386
rect 18338 52334 18340 52386
rect 18284 52322 18340 52334
rect 18396 52388 18452 52398
rect 18172 52164 18228 52174
rect 17948 52162 18228 52164
rect 17948 52110 18174 52162
rect 18226 52110 18228 52162
rect 17948 52108 18228 52110
rect 18172 52098 18228 52108
rect 18172 51940 18228 51950
rect 18172 51846 18228 51884
rect 18284 51828 18340 51838
rect 17948 51604 18004 51614
rect 17948 51510 18004 51548
rect 18172 51380 18228 51390
rect 18172 51286 18228 51324
rect 18284 51156 18340 51772
rect 18172 51100 18340 51156
rect 17836 50372 18004 50428
rect 17612 49698 17668 49710
rect 17612 49646 17614 49698
rect 17666 49646 17668 49698
rect 17612 47908 17668 49646
rect 17724 49028 17780 50316
rect 17724 48962 17780 48972
rect 17948 48580 18004 50372
rect 18172 49028 18228 51100
rect 18284 50484 18340 50522
rect 18284 50418 18340 50428
rect 18396 50428 18452 52332
rect 18508 52386 18564 52668
rect 18508 52334 18510 52386
rect 18562 52334 18564 52386
rect 18508 52322 18564 52334
rect 18396 50372 18564 50428
rect 18508 49812 18564 50372
rect 18396 49698 18452 49710
rect 18396 49646 18398 49698
rect 18450 49646 18452 49698
rect 18284 49028 18340 49038
rect 17724 48524 18004 48580
rect 18060 49026 18340 49028
rect 18060 48974 18286 49026
rect 18338 48974 18340 49026
rect 18060 48972 18340 48974
rect 17724 48244 17780 48524
rect 17724 48150 17780 48188
rect 17836 48356 17892 48366
rect 17612 47852 17780 47908
rect 17388 47628 17556 47684
rect 17612 47682 17668 47694
rect 17612 47630 17614 47682
rect 17666 47630 17668 47682
rect 17388 46900 17444 47628
rect 17612 47572 17668 47630
rect 17612 47506 17668 47516
rect 17500 47460 17556 47498
rect 17500 47394 17556 47404
rect 17388 46834 17444 46844
rect 17500 47236 17556 47246
rect 17500 46676 17556 47180
rect 17388 46620 17556 46676
rect 17612 46900 17668 46910
rect 17388 44546 17444 46620
rect 17500 46340 17556 46350
rect 17500 45666 17556 46284
rect 17500 45614 17502 45666
rect 17554 45614 17556 45666
rect 17500 45220 17556 45614
rect 17500 45154 17556 45164
rect 17388 44494 17390 44546
rect 17442 44494 17444 44546
rect 17388 44482 17444 44494
rect 17500 44436 17556 44446
rect 17500 44210 17556 44380
rect 17500 44158 17502 44210
rect 17554 44158 17556 44210
rect 17388 44100 17444 44110
rect 17388 44006 17444 44044
rect 17500 43876 17556 44158
rect 17500 43810 17556 43820
rect 17612 43316 17668 46844
rect 17724 44436 17780 47852
rect 17836 44996 17892 48300
rect 18060 46900 18116 48972
rect 18284 48962 18340 48972
rect 18396 48468 18452 49646
rect 18508 49364 18564 49756
rect 18620 50370 18676 50382
rect 18620 50318 18622 50370
rect 18674 50318 18676 50370
rect 18620 49700 18676 50318
rect 18620 49634 18676 49644
rect 18508 49298 18564 49308
rect 18620 49140 18676 49150
rect 18620 49046 18676 49084
rect 18508 49028 18564 49038
rect 18508 48580 18564 48972
rect 18620 48804 18676 48814
rect 18620 48710 18676 48748
rect 18508 48514 18564 48524
rect 18732 48468 18788 53004
rect 18956 52834 19012 52846
rect 18956 52782 18958 52834
rect 19010 52782 19012 52834
rect 18844 52500 18900 52510
rect 18844 50036 18900 52444
rect 18956 51604 19012 52782
rect 19068 52724 19124 54348
rect 19180 53508 19236 53518
rect 19180 53414 19236 53452
rect 19404 52836 19460 52846
rect 19292 52834 19460 52836
rect 19292 52782 19406 52834
rect 19458 52782 19460 52834
rect 19292 52780 19460 52782
rect 19180 52724 19236 52734
rect 19068 52722 19236 52724
rect 19068 52670 19182 52722
rect 19234 52670 19236 52722
rect 19068 52668 19236 52670
rect 19180 52274 19236 52668
rect 19180 52222 19182 52274
rect 19234 52222 19236 52274
rect 19180 52210 19236 52222
rect 18956 51538 19012 51548
rect 19180 52052 19236 52062
rect 18956 51378 19012 51390
rect 18956 51326 18958 51378
rect 19010 51326 19012 51378
rect 18956 51156 19012 51326
rect 18956 51090 19012 51100
rect 19180 50932 19236 51996
rect 19292 51828 19348 52780
rect 19404 52770 19460 52780
rect 19404 52388 19460 52398
rect 19516 52388 19572 55468
rect 19852 55410 19908 55580
rect 19852 55358 19854 55410
rect 19906 55358 19908 55410
rect 19852 55346 19908 55358
rect 20300 55522 20356 55534
rect 20300 55470 20302 55522
rect 20354 55470 20356 55522
rect 20300 55410 20356 55470
rect 20300 55358 20302 55410
rect 20354 55358 20356 55410
rect 20300 55346 20356 55358
rect 20748 55076 20804 55918
rect 21084 55970 21364 55972
rect 21084 55918 21310 55970
rect 21362 55918 21364 55970
rect 21084 55916 21364 55918
rect 20860 55860 20916 55870
rect 20860 55858 21028 55860
rect 20860 55806 20862 55858
rect 20914 55806 21028 55858
rect 20860 55804 21028 55806
rect 20860 55794 20916 55804
rect 20860 55076 20916 55086
rect 20748 55074 20916 55076
rect 20748 55022 20862 55074
rect 20914 55022 20916 55074
rect 20748 55020 20916 55022
rect 20860 54964 20916 55020
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20860 54898 20916 54908
rect 19836 54842 20100 54852
rect 20412 54740 20468 54750
rect 20412 54646 20468 54684
rect 20524 54740 20580 54750
rect 20524 54738 20916 54740
rect 20524 54686 20526 54738
rect 20578 54686 20916 54738
rect 20524 54684 20916 54686
rect 20524 54674 20580 54684
rect 20636 54516 20692 54526
rect 20412 54514 20692 54516
rect 20412 54462 20638 54514
rect 20690 54462 20692 54514
rect 20412 54460 20692 54462
rect 19740 54404 19796 54414
rect 19628 54402 19796 54404
rect 19628 54350 19742 54402
rect 19794 54350 19796 54402
rect 19628 54348 19796 54350
rect 19628 53172 19684 54348
rect 19740 54338 19796 54348
rect 20412 53956 20468 54460
rect 20636 54450 20692 54460
rect 20748 54516 20804 54526
rect 20748 54422 20804 54460
rect 20524 53956 20580 53966
rect 20412 53954 20580 53956
rect 20412 53902 20526 53954
rect 20578 53902 20580 53954
rect 20412 53900 20580 53902
rect 20524 53890 20580 53900
rect 19964 53732 20020 53742
rect 19964 53638 20020 53676
rect 20188 53732 20244 53742
rect 20188 53730 20468 53732
rect 20188 53678 20190 53730
rect 20242 53678 20468 53730
rect 20188 53676 20468 53678
rect 20188 53666 20244 53676
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19628 53116 19908 53172
rect 19460 52332 19572 52388
rect 19404 52256 19460 52332
rect 19292 51762 19348 51772
rect 19628 52162 19684 52174
rect 19628 52110 19630 52162
rect 19682 52110 19684 52162
rect 19292 51604 19348 51614
rect 19628 51604 19684 52110
rect 19852 52052 19908 53116
rect 20188 52836 20244 52846
rect 20188 52742 20244 52780
rect 20076 52500 20132 52510
rect 20076 52386 20132 52444
rect 20076 52334 20078 52386
rect 20130 52334 20132 52386
rect 20076 52322 20132 52334
rect 19852 51986 19908 51996
rect 20188 52164 20244 52174
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19292 51602 19684 51604
rect 19292 51550 19294 51602
rect 19346 51550 19684 51602
rect 19292 51548 19684 51550
rect 20188 51602 20244 52108
rect 20188 51550 20190 51602
rect 20242 51550 20244 51602
rect 19292 51538 19348 51548
rect 20188 51538 20244 51550
rect 19180 50594 19236 50876
rect 19404 51378 19460 51390
rect 19404 51326 19406 51378
rect 19458 51326 19460 51378
rect 19404 50708 19460 51326
rect 19404 50642 19460 50652
rect 19516 51378 19572 51390
rect 19516 51326 19518 51378
rect 19570 51326 19572 51378
rect 19180 50542 19182 50594
rect 19234 50542 19236 50594
rect 19180 50530 19236 50542
rect 19516 50372 19572 51326
rect 20412 51156 20468 53676
rect 20524 53172 20580 53182
rect 20524 52612 20580 53116
rect 20524 52546 20580 52556
rect 20636 52948 20692 52958
rect 20524 52276 20580 52286
rect 20524 52162 20580 52220
rect 20524 52110 20526 52162
rect 20578 52110 20580 52162
rect 20524 52098 20580 52110
rect 20636 52164 20692 52892
rect 20860 52388 20916 54684
rect 20636 52050 20692 52108
rect 20636 51998 20638 52050
rect 20690 51998 20692 52050
rect 20636 51986 20692 51998
rect 20748 52332 20916 52388
rect 20972 53172 21028 55804
rect 21084 55524 21140 55916
rect 21308 55906 21364 55916
rect 21084 55522 21252 55524
rect 21084 55470 21086 55522
rect 21138 55470 21252 55522
rect 21084 55468 21252 55470
rect 21084 55458 21140 55468
rect 21084 55300 21140 55310
rect 21084 54514 21140 55244
rect 21084 54462 21086 54514
rect 21138 54462 21140 54514
rect 21084 54450 21140 54462
rect 20748 51716 20804 52332
rect 20860 52164 20916 52174
rect 20860 52070 20916 52108
rect 20972 51828 21028 53116
rect 21196 52948 21252 55468
rect 21644 54514 21700 56028
rect 22540 56084 22596 56094
rect 22540 55990 22596 56028
rect 22092 55972 22148 55982
rect 22092 55970 22260 55972
rect 22092 55918 22094 55970
rect 22146 55918 22260 55970
rect 22092 55916 22260 55918
rect 22092 55906 22148 55916
rect 22092 55298 22148 55310
rect 22092 55246 22094 55298
rect 22146 55246 22148 55298
rect 22092 55076 22148 55246
rect 22204 55188 22260 55916
rect 22652 55860 22708 55870
rect 22652 55766 22708 55804
rect 22204 55122 22260 55132
rect 22092 54738 22148 55020
rect 22316 55076 22372 55086
rect 22316 54982 22372 55020
rect 22764 54964 22820 56140
rect 23548 55970 23604 59200
rect 25900 57204 25956 57214
rect 23548 55918 23550 55970
rect 23602 55918 23604 55970
rect 23548 55906 23604 55918
rect 24444 56084 24500 56094
rect 23548 55412 23604 55422
rect 22764 54898 22820 54908
rect 23100 55186 23156 55198
rect 23100 55134 23102 55186
rect 23154 55134 23156 55186
rect 22092 54686 22094 54738
rect 22146 54686 22148 54738
rect 22092 54674 22148 54686
rect 22204 54740 22260 54750
rect 21644 54462 21646 54514
rect 21698 54462 21700 54514
rect 21196 52816 21252 52892
rect 21308 54404 21364 54414
rect 21308 52724 21364 54348
rect 21644 54180 21700 54462
rect 21868 54514 21924 54526
rect 21868 54462 21870 54514
rect 21922 54462 21924 54514
rect 21644 54114 21700 54124
rect 21756 54402 21812 54414
rect 21756 54350 21758 54402
rect 21810 54350 21812 54402
rect 21644 53732 21700 53742
rect 21756 53732 21812 54350
rect 21868 54404 21924 54462
rect 21868 54338 21924 54348
rect 22092 54516 22148 54526
rect 21644 53730 21812 53732
rect 21644 53678 21646 53730
rect 21698 53678 21812 53730
rect 21644 53676 21812 53678
rect 21644 53666 21700 53676
rect 21868 53508 21924 53518
rect 22092 53508 22148 54460
rect 22204 53954 22260 54684
rect 22764 54404 22820 54414
rect 22204 53902 22206 53954
rect 22258 53902 22260 53954
rect 22204 53890 22260 53902
rect 22316 54402 22820 54404
rect 22316 54350 22766 54402
rect 22818 54350 22820 54402
rect 22316 54348 22820 54350
rect 21644 53506 21924 53508
rect 21644 53454 21870 53506
rect 21922 53454 21924 53506
rect 21644 53452 21924 53454
rect 20748 51650 20804 51660
rect 20860 51772 21028 51828
rect 21196 52668 21364 52724
rect 21420 53058 21476 53070
rect 21420 53006 21422 53058
rect 21474 53006 21476 53058
rect 21420 52836 21476 53006
rect 20524 51604 20580 51614
rect 20524 51510 20580 51548
rect 20860 51380 20916 51772
rect 20860 51314 20916 51324
rect 20972 51604 21028 51614
rect 20412 51100 20580 51156
rect 20188 50932 20244 50942
rect 20076 50708 20132 50718
rect 18844 49970 18900 49980
rect 19404 50370 19572 50372
rect 19404 50318 19518 50370
rect 19570 50318 19572 50370
rect 19404 50316 19572 50318
rect 18956 49924 19012 49934
rect 18844 49700 18900 49710
rect 18844 49606 18900 49644
rect 18284 48412 18452 48468
rect 18620 48412 18788 48468
rect 18844 49028 18900 49038
rect 18956 49028 19012 49868
rect 19404 49924 19460 50316
rect 19516 50306 19572 50316
rect 19628 50596 19684 50606
rect 19628 49924 19684 50540
rect 20076 50594 20132 50652
rect 20076 50542 20078 50594
rect 20130 50542 20132 50594
rect 20076 50530 20132 50542
rect 20188 50370 20244 50876
rect 20188 50318 20190 50370
rect 20242 50318 20244 50370
rect 20188 50306 20244 50318
rect 20412 50370 20468 50382
rect 20412 50318 20414 50370
rect 20466 50318 20468 50370
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19852 50036 19908 50046
rect 19852 49942 19908 49980
rect 19964 50036 20020 50046
rect 19964 50034 20244 50036
rect 19964 49982 19966 50034
rect 20018 49982 20244 50034
rect 19964 49980 20244 49982
rect 19964 49970 20020 49980
rect 19628 49868 19796 49924
rect 19404 49586 19460 49868
rect 19404 49534 19406 49586
rect 19458 49534 19460 49586
rect 19404 49522 19460 49534
rect 19628 49698 19684 49710
rect 19628 49646 19630 49698
rect 19682 49646 19684 49698
rect 19628 49588 19684 49646
rect 19740 49700 19796 49868
rect 20076 49812 20132 49822
rect 20076 49718 20132 49756
rect 19740 49644 19908 49700
rect 19628 49522 19684 49532
rect 18900 48972 19012 49028
rect 19068 49476 19124 49486
rect 19068 49026 19124 49420
rect 19068 48974 19070 49026
rect 19122 48974 19124 49026
rect 18172 48356 18228 48366
rect 18172 48262 18228 48300
rect 18060 46834 18116 46844
rect 18172 47684 18228 47694
rect 18060 46674 18116 46686
rect 18060 46622 18062 46674
rect 18114 46622 18116 46674
rect 17948 46116 18004 46126
rect 17948 46002 18004 46060
rect 17948 45950 17950 46002
rect 18002 45950 18004 46002
rect 17948 45668 18004 45950
rect 17948 45602 18004 45612
rect 17948 44996 18004 45006
rect 17836 44994 18004 44996
rect 17836 44942 17950 44994
rect 18002 44942 18004 44994
rect 17836 44940 18004 44942
rect 17724 44100 17780 44380
rect 17724 44034 17780 44044
rect 17724 43540 17780 43550
rect 17724 43446 17780 43484
rect 17500 43260 17668 43316
rect 17500 42980 17556 43260
rect 17948 42980 18004 44940
rect 18060 44996 18116 46622
rect 18060 44930 18116 44940
rect 18172 44436 18228 47628
rect 18284 46564 18340 48412
rect 18396 48244 18452 48254
rect 18396 48150 18452 48188
rect 18508 46900 18564 46910
rect 18620 46900 18676 48412
rect 18844 48242 18900 48972
rect 19068 48356 19124 48974
rect 19068 48290 19124 48300
rect 19180 49364 19236 49374
rect 18844 48190 18846 48242
rect 18898 48190 18900 48242
rect 18844 48178 18900 48190
rect 18508 46898 18676 46900
rect 18508 46846 18510 46898
rect 18562 46846 18676 46898
rect 18508 46844 18676 46846
rect 18732 48132 18788 48142
rect 18508 46834 18564 46844
rect 18396 46676 18452 46686
rect 18396 46582 18452 46620
rect 18620 46674 18676 46686
rect 18620 46622 18622 46674
rect 18674 46622 18676 46674
rect 18284 45556 18340 46508
rect 18620 46452 18676 46622
rect 18620 46386 18676 46396
rect 18284 45490 18340 45500
rect 18396 46114 18452 46126
rect 18396 46062 18398 46114
rect 18450 46062 18452 46114
rect 18396 46002 18452 46062
rect 18396 45950 18398 46002
rect 18450 45950 18452 46002
rect 18284 44436 18340 44446
rect 18172 44434 18340 44436
rect 18172 44382 18286 44434
rect 18338 44382 18340 44434
rect 18172 44380 18340 44382
rect 18284 44100 18340 44380
rect 18284 44034 18340 44044
rect 18396 43876 18452 45950
rect 18732 45892 18788 48076
rect 18956 47796 19012 47806
rect 18956 47570 19012 47740
rect 18956 47518 18958 47570
rect 19010 47518 19012 47570
rect 18956 47506 19012 47518
rect 19068 46900 19124 46910
rect 19068 46806 19124 46844
rect 19180 46116 19236 49308
rect 19628 49364 19684 49374
rect 19404 49140 19460 49150
rect 19292 48692 19348 48702
rect 19292 48242 19348 48636
rect 19292 48190 19294 48242
rect 19346 48190 19348 48242
rect 19292 48132 19348 48190
rect 19292 48066 19348 48076
rect 19180 46050 19236 46060
rect 19292 47684 19348 47694
rect 18284 43820 18452 43876
rect 18508 45836 18788 45892
rect 18508 44884 18564 45836
rect 18844 45780 18900 45790
rect 18284 43540 18340 43820
rect 18508 43652 18564 44828
rect 18508 43586 18564 43596
rect 18620 45778 18900 45780
rect 18620 45726 18846 45778
rect 18898 45726 18900 45778
rect 18620 45724 18900 45726
rect 18620 43876 18676 45724
rect 18844 45714 18900 45724
rect 18844 45556 18900 45566
rect 18844 45220 18900 45500
rect 18732 45218 18900 45220
rect 18732 45166 18846 45218
rect 18898 45166 18900 45218
rect 18732 45164 18900 45166
rect 18732 44322 18788 45164
rect 18844 45108 18900 45164
rect 18956 45220 19012 45230
rect 18956 45218 19124 45220
rect 18956 45166 18958 45218
rect 19010 45166 19124 45218
rect 18956 45164 19124 45166
rect 18956 45154 19012 45164
rect 18844 45042 18900 45052
rect 18844 44884 18900 44894
rect 18844 44434 18900 44828
rect 18956 44882 19012 44894
rect 18956 44830 18958 44882
rect 19010 44830 19012 44882
rect 18956 44548 19012 44830
rect 19068 44772 19124 45164
rect 19292 44772 19348 47628
rect 19404 45220 19460 49084
rect 19628 49028 19684 49308
rect 19852 49138 19908 49644
rect 20188 49364 20244 49980
rect 20412 49924 20468 50318
rect 20412 49858 20468 49868
rect 19852 49086 19854 49138
rect 19906 49086 19908 49138
rect 19852 49074 19908 49086
rect 19964 49308 20244 49364
rect 19964 49140 20020 49308
rect 20188 49140 20244 49150
rect 19964 49074 20020 49084
rect 20076 49084 20188 49140
rect 19740 49028 19796 49038
rect 19628 49026 19796 49028
rect 19628 48974 19742 49026
rect 19794 48974 19796 49026
rect 19628 48972 19796 48974
rect 19740 48962 19796 48972
rect 19964 48916 20020 48926
rect 20076 48916 20132 49084
rect 20188 49074 20244 49084
rect 19964 48914 20132 48916
rect 19964 48862 19966 48914
rect 20018 48862 20132 48914
rect 19964 48860 20132 48862
rect 19964 48850 20020 48860
rect 20188 48802 20244 48814
rect 20188 48750 20190 48802
rect 20242 48750 20244 48802
rect 19516 48692 19572 48702
rect 19516 46900 19572 48636
rect 19836 48636 20100 48646
rect 19628 48580 19684 48590
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19628 48356 19684 48524
rect 19852 48356 19908 48366
rect 19628 48354 19908 48356
rect 19628 48302 19854 48354
rect 19906 48302 19908 48354
rect 19628 48300 19908 48302
rect 19852 48290 19908 48300
rect 19964 48356 20020 48366
rect 19852 48020 19908 48030
rect 19852 47684 19908 47964
rect 19628 47460 19684 47470
rect 19628 47366 19684 47404
rect 19852 47458 19908 47628
rect 19852 47406 19854 47458
rect 19906 47406 19908 47458
rect 19852 47394 19908 47406
rect 19964 47458 20020 48300
rect 20076 48354 20132 48366
rect 20076 48302 20078 48354
rect 20130 48302 20132 48354
rect 20076 48132 20132 48302
rect 20076 48066 20132 48076
rect 20188 48130 20244 48750
rect 20188 48078 20190 48130
rect 20242 48078 20244 48130
rect 20188 47684 20244 48078
rect 20188 47618 20244 47628
rect 20300 48804 20356 48814
rect 20300 47682 20356 48748
rect 20524 48580 20580 51100
rect 20860 50372 20916 50382
rect 20524 48514 20580 48524
rect 20636 50370 20916 50372
rect 20636 50318 20862 50370
rect 20914 50318 20916 50370
rect 20636 50316 20916 50318
rect 20636 48356 20692 50316
rect 20860 50306 20916 50316
rect 20524 48300 20692 48356
rect 20748 49700 20804 49710
rect 20748 48916 20804 49644
rect 20748 48802 20804 48860
rect 20748 48750 20750 48802
rect 20802 48750 20804 48802
rect 20524 48020 20580 48300
rect 20524 47954 20580 47964
rect 20636 48130 20692 48142
rect 20636 48078 20638 48130
rect 20690 48078 20692 48130
rect 20300 47630 20302 47682
rect 20354 47630 20356 47682
rect 20300 47618 20356 47630
rect 20524 47684 20580 47694
rect 20524 47590 20580 47628
rect 19964 47406 19966 47458
rect 20018 47406 20020 47458
rect 19964 47348 20020 47406
rect 19964 47282 20020 47292
rect 19740 47236 19796 47274
rect 19740 47170 19796 47180
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19852 46900 19908 46910
rect 19516 46898 19908 46900
rect 19516 46846 19854 46898
rect 19906 46846 19908 46898
rect 19516 46844 19908 46846
rect 19852 46834 19908 46844
rect 19964 46900 20020 46910
rect 19628 46676 19684 46686
rect 19964 46676 20020 46844
rect 19628 46582 19684 46620
rect 19852 46620 20020 46676
rect 20076 46674 20132 46686
rect 20076 46622 20078 46674
rect 20130 46622 20132 46674
rect 19740 46564 19796 46574
rect 19740 46470 19796 46508
rect 19516 45778 19572 45790
rect 19516 45726 19518 45778
rect 19570 45726 19572 45778
rect 19516 45668 19572 45726
rect 19852 45780 19908 46620
rect 20076 46452 20132 46622
rect 20076 46386 20132 46396
rect 20412 46674 20468 46686
rect 20412 46622 20414 46674
rect 20466 46622 20468 46674
rect 20300 46116 20356 46126
rect 19852 45778 20132 45780
rect 19852 45726 19854 45778
rect 19906 45726 20132 45778
rect 19852 45724 20132 45726
rect 19852 45714 19908 45724
rect 20076 45668 20132 45724
rect 20076 45612 20244 45668
rect 19516 45602 19572 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20188 45332 20244 45612
rect 20076 45276 20244 45332
rect 19404 45154 19460 45164
rect 19740 45218 19796 45230
rect 19740 45166 19742 45218
rect 19794 45166 19796 45218
rect 19628 45106 19684 45118
rect 19628 45054 19630 45106
rect 19682 45054 19684 45106
rect 19628 44884 19684 45054
rect 19740 45108 19796 45166
rect 19740 45042 19796 45052
rect 19628 44818 19684 44828
rect 19292 44716 19572 44772
rect 19068 44706 19124 44716
rect 18956 44482 19012 44492
rect 18844 44382 18846 44434
rect 18898 44382 18900 44434
rect 18844 44370 18900 44382
rect 19068 44436 19124 44446
rect 18732 44270 18734 44322
rect 18786 44270 18788 44322
rect 18732 44258 18788 44270
rect 19068 44324 19124 44380
rect 19292 44324 19348 44334
rect 19068 44322 19348 44324
rect 19068 44270 19294 44322
rect 19346 44270 19348 44322
rect 19068 44268 19348 44270
rect 19292 44258 19348 44268
rect 18956 44100 19012 44110
rect 18844 44098 19012 44100
rect 18844 44046 18958 44098
rect 19010 44046 19012 44098
rect 18844 44044 19012 44046
rect 18844 43988 18900 44044
rect 18956 44034 19012 44044
rect 18844 43922 18900 43932
rect 18060 43428 18116 43438
rect 18060 43426 18228 43428
rect 18060 43374 18062 43426
rect 18114 43374 18228 43426
rect 18060 43372 18228 43374
rect 18060 43362 18116 43372
rect 17500 42914 17556 42924
rect 17612 42924 18004 42980
rect 18060 42980 18116 42990
rect 17388 42532 17444 42542
rect 17388 42438 17444 42476
rect 17276 42252 17444 42308
rect 16940 41972 16996 41982
rect 16940 41878 16996 41916
rect 16828 41692 16996 41748
rect 16604 41076 16660 41692
rect 16604 41074 16772 41076
rect 16604 41022 16606 41074
rect 16658 41022 16772 41074
rect 16604 41020 16772 41022
rect 16604 41010 16660 41020
rect 16604 40852 16660 40862
rect 16604 40626 16660 40796
rect 16604 40574 16606 40626
rect 16658 40574 16660 40626
rect 16156 38834 16212 39676
rect 16156 38782 16158 38834
rect 16210 38782 16212 38834
rect 16380 40516 16436 40526
rect 16380 38948 16436 40460
rect 16604 40516 16660 40574
rect 16604 40450 16660 40460
rect 16492 39396 16548 39406
rect 16492 39394 16660 39396
rect 16492 39342 16494 39394
rect 16546 39342 16660 39394
rect 16492 39340 16660 39342
rect 16492 39330 16548 39340
rect 16380 38816 16436 38892
rect 16492 39060 16548 39070
rect 16492 38946 16548 39004
rect 16492 38894 16494 38946
rect 16546 38894 16548 38946
rect 16156 38770 16212 38782
rect 16492 38668 16548 38894
rect 16044 38546 16100 38556
rect 16380 38612 16548 38668
rect 16044 37940 16100 37950
rect 16044 37846 16100 37884
rect 16268 36484 16324 36494
rect 16268 36390 16324 36428
rect 16156 36372 16212 36382
rect 16156 36278 16212 36316
rect 16268 36148 16324 36158
rect 16268 35812 16324 36092
rect 16044 35586 16100 35598
rect 16044 35534 16046 35586
rect 16098 35534 16100 35586
rect 16044 35476 16100 35534
rect 16044 35410 16100 35420
rect 15820 33516 15988 33572
rect 16044 34804 16100 34814
rect 16044 34132 16100 34748
rect 16268 34804 16324 35756
rect 16268 34738 16324 34748
rect 16156 34580 16212 34590
rect 16156 34354 16212 34524
rect 16156 34302 16158 34354
rect 16210 34302 16212 34354
rect 16156 34290 16212 34302
rect 14924 33348 14980 33358
rect 14924 33254 14980 33292
rect 15260 33122 15316 33134
rect 15260 33070 15262 33122
rect 15314 33070 15316 33122
rect 15260 33012 15316 33070
rect 15148 32788 15204 32798
rect 15148 32694 15204 32732
rect 14812 32622 14814 32674
rect 14866 32622 14868 32674
rect 14140 31668 14196 31678
rect 14364 31668 14420 32396
rect 14588 31892 14644 31902
rect 14812 31892 14868 32622
rect 15260 32452 15316 32956
rect 15260 32386 15316 32396
rect 15708 32452 15764 32462
rect 14588 31890 14868 31892
rect 14588 31838 14590 31890
rect 14642 31838 14868 31890
rect 14588 31836 14868 31838
rect 14924 31892 14980 31902
rect 14588 31826 14644 31836
rect 14924 31798 14980 31836
rect 15708 31890 15764 32396
rect 15708 31838 15710 31890
rect 15762 31838 15764 31890
rect 15708 31826 15764 31838
rect 14140 31574 14196 31612
rect 14252 31612 14420 31668
rect 14476 31780 14532 31790
rect 14140 31220 14196 31230
rect 14140 31126 14196 31164
rect 14028 30930 14084 30940
rect 13692 29988 13748 29998
rect 13468 29986 13748 29988
rect 13468 29934 13694 29986
rect 13746 29934 13748 29986
rect 13468 29932 13748 29934
rect 11676 29316 11732 29326
rect 11676 29222 11732 29260
rect 12348 29204 12404 29932
rect 12348 29138 12404 29148
rect 13356 29314 13412 29326
rect 13356 29262 13358 29314
rect 13410 29262 13412 29314
rect 13356 28980 13412 29262
rect 13356 28914 13412 28924
rect 13692 28532 13748 29932
rect 13692 28466 13748 28476
rect 14028 29540 14084 29550
rect 14028 28642 14084 29484
rect 14028 28590 14030 28642
rect 14082 28590 14084 28642
rect 13468 27858 13524 27870
rect 14028 27860 14084 28590
rect 14252 29426 14308 31612
rect 14476 31220 14532 31724
rect 14588 31220 14644 31230
rect 14476 31218 14644 31220
rect 14476 31166 14590 31218
rect 14642 31166 14644 31218
rect 14476 31164 14644 31166
rect 14588 31108 14644 31164
rect 15484 31220 15540 31230
rect 15484 31126 15540 31164
rect 14588 31042 14644 31052
rect 15260 31108 15316 31118
rect 15260 31014 15316 31052
rect 15036 30994 15092 31006
rect 15036 30942 15038 30994
rect 15090 30942 15092 30994
rect 15036 30884 15092 30942
rect 15036 30818 15092 30828
rect 15148 30882 15204 30894
rect 15148 30830 15150 30882
rect 15202 30830 15204 30882
rect 14700 30436 14756 30446
rect 14700 30342 14756 30380
rect 15148 30436 15204 30830
rect 15148 30370 15204 30380
rect 15260 30884 15316 30894
rect 14924 30212 14980 30222
rect 14252 29374 14254 29426
rect 14306 29374 14308 29426
rect 14252 28084 14308 29374
rect 14252 28018 14308 28028
rect 14364 29986 14420 29998
rect 14364 29934 14366 29986
rect 14418 29934 14420 29986
rect 13468 27806 13470 27858
rect 13522 27806 13524 27858
rect 13468 27412 13524 27806
rect 13468 27346 13524 27356
rect 13580 27858 14084 27860
rect 13580 27806 14030 27858
rect 14082 27806 14084 27858
rect 13580 27804 14084 27806
rect 13020 26964 13076 27002
rect 11564 26852 11732 26908
rect 11340 26798 11342 26850
rect 11394 26798 11396 26850
rect 11340 26786 11396 26798
rect 11676 24276 11732 26852
rect 11676 24210 11732 24220
rect 13020 14308 13076 26908
rect 13580 26292 13636 27804
rect 14028 27794 14084 27804
rect 13804 26964 13860 27002
rect 13804 26898 13860 26908
rect 14364 26908 14420 29934
rect 14700 29426 14756 29438
rect 14700 29374 14702 29426
rect 14754 29374 14756 29426
rect 14700 28980 14756 29374
rect 14812 29428 14868 29438
rect 14812 29334 14868 29372
rect 14924 29316 14980 30156
rect 14924 29250 14980 29260
rect 14700 28914 14756 28924
rect 14476 28644 14532 28654
rect 14476 28550 14532 28588
rect 14588 27970 14644 27982
rect 14588 27918 14590 27970
rect 14642 27918 14644 27970
rect 14588 27860 14644 27918
rect 14588 27794 14644 27804
rect 14924 27858 14980 27870
rect 14924 27806 14926 27858
rect 14978 27806 14980 27858
rect 14924 27412 14980 27806
rect 15148 27412 15204 27422
rect 14924 27356 15148 27412
rect 15148 27186 15204 27356
rect 15148 27134 15150 27186
rect 15202 27134 15204 27186
rect 15148 27122 15204 27134
rect 14364 26852 14644 26908
rect 14028 26292 14084 26302
rect 13580 26290 13972 26292
rect 13580 26238 13582 26290
rect 13634 26238 13972 26290
rect 13580 26236 13972 26238
rect 13580 26226 13636 26236
rect 13916 25172 13972 26236
rect 14028 26290 14420 26292
rect 14028 26238 14030 26290
rect 14082 26238 14420 26290
rect 14028 26236 14420 26238
rect 14028 26226 14084 26236
rect 14364 25394 14420 26236
rect 14588 25506 14644 26852
rect 14588 25454 14590 25506
rect 14642 25454 14644 25506
rect 14588 25442 14644 25454
rect 14364 25342 14366 25394
rect 14418 25342 14420 25394
rect 14364 25330 14420 25342
rect 15260 25396 15316 30828
rect 15708 30324 15764 30334
rect 15596 30212 15652 30222
rect 15596 30118 15652 30156
rect 15708 30210 15764 30268
rect 15708 30158 15710 30210
rect 15762 30158 15764 30210
rect 15708 30146 15764 30158
rect 15820 29764 15876 33516
rect 15932 33346 15988 33358
rect 15932 33294 15934 33346
rect 15986 33294 15988 33346
rect 15932 33012 15988 33294
rect 15932 32788 15988 32956
rect 15932 32722 15988 32732
rect 16044 31892 16100 34076
rect 16156 33236 16212 33246
rect 16156 33142 16212 33180
rect 16268 33012 16324 33022
rect 16268 32562 16324 32956
rect 16380 32788 16436 38612
rect 16604 38052 16660 39340
rect 16492 37940 16548 37950
rect 16492 37846 16548 37884
rect 16604 37828 16660 37996
rect 16604 37762 16660 37772
rect 16716 37492 16772 41020
rect 16940 40964 16996 41692
rect 16828 40908 16996 40964
rect 17164 41188 17220 41198
rect 17276 41188 17332 41198
rect 17220 41186 17332 41188
rect 17220 41134 17278 41186
rect 17330 41134 17332 41186
rect 17220 41132 17332 41134
rect 16828 39284 16884 40908
rect 16940 40740 16996 40750
rect 16940 40404 16996 40684
rect 17164 40740 17220 41132
rect 17276 41122 17332 41132
rect 17388 40964 17444 42252
rect 17164 40674 17220 40684
rect 17276 40908 17444 40964
rect 17500 41972 17556 41982
rect 16940 40310 16996 40348
rect 16940 39844 16996 39854
rect 16940 39750 16996 39788
rect 17052 39732 17108 39742
rect 17052 39618 17108 39676
rect 17052 39566 17054 39618
rect 17106 39566 17108 39618
rect 17052 39554 17108 39566
rect 16828 39228 17108 39284
rect 16940 38836 16996 38846
rect 16940 38742 16996 38780
rect 17052 38668 17108 39228
rect 16716 37426 16772 37436
rect 16828 38612 17108 38668
rect 16604 37268 16660 37278
rect 16492 37266 16660 37268
rect 16492 37214 16606 37266
rect 16658 37214 16660 37266
rect 16492 37212 16660 37214
rect 16492 35364 16548 37212
rect 16604 37202 16660 37212
rect 16604 36932 16660 36942
rect 16604 35922 16660 36876
rect 16604 35870 16606 35922
rect 16658 35870 16660 35922
rect 16604 35858 16660 35870
rect 16492 35298 16548 35308
rect 16716 35364 16772 35374
rect 16604 34804 16660 34814
rect 16492 34130 16548 34142
rect 16492 34078 16494 34130
rect 16546 34078 16548 34130
rect 16492 33124 16548 34078
rect 16604 33348 16660 34748
rect 16716 34802 16772 35308
rect 16716 34750 16718 34802
rect 16770 34750 16772 34802
rect 16716 34738 16772 34750
rect 16604 33282 16660 33292
rect 16716 33346 16772 33358
rect 16716 33294 16718 33346
rect 16770 33294 16772 33346
rect 16716 33124 16772 33294
rect 16492 33068 16772 33124
rect 16492 33012 16548 33068
rect 16492 32946 16548 32956
rect 16828 32900 16884 38612
rect 16940 37940 16996 37950
rect 16940 37846 16996 37884
rect 16940 37492 16996 37502
rect 16940 37398 16996 37436
rect 17164 36596 17220 36606
rect 17164 36482 17220 36540
rect 17164 36430 17166 36482
rect 17218 36430 17220 36482
rect 17164 36418 17220 36430
rect 17164 36260 17220 36270
rect 17052 35812 17108 35822
rect 16940 35700 16996 35710
rect 16940 35364 16996 35644
rect 16940 35298 16996 35308
rect 16940 34916 16996 34926
rect 17052 34916 17108 35756
rect 16940 34914 17108 34916
rect 16940 34862 16942 34914
rect 16994 34862 17108 34914
rect 16940 34860 17108 34862
rect 16940 34850 16996 34860
rect 16940 34580 16996 34590
rect 16940 34354 16996 34524
rect 16940 34302 16942 34354
rect 16994 34302 16996 34354
rect 16940 34290 16996 34302
rect 16940 33348 16996 33358
rect 16940 33254 16996 33292
rect 16828 32844 17108 32900
rect 16380 32732 16660 32788
rect 16604 32676 16660 32732
rect 16604 32620 16772 32676
rect 16268 32510 16270 32562
rect 16322 32510 16324 32562
rect 16268 32498 16324 32510
rect 16716 32564 16772 32620
rect 16940 32564 16996 32574
rect 16716 32562 16996 32564
rect 16716 32510 16942 32562
rect 16994 32510 16996 32562
rect 16716 32508 16996 32510
rect 16940 32498 16996 32508
rect 16604 32452 16660 32462
rect 16604 32358 16660 32396
rect 17052 32116 17108 32844
rect 16940 32060 17108 32116
rect 16156 31892 16212 31902
rect 16044 31890 16212 31892
rect 16044 31838 16158 31890
rect 16210 31838 16212 31890
rect 16044 31836 16212 31838
rect 16156 31826 16212 31836
rect 16940 31780 16996 32060
rect 17052 31892 17108 31902
rect 17164 31892 17220 36204
rect 17276 35924 17332 40908
rect 17388 40740 17444 40750
rect 17388 36148 17444 40684
rect 17500 40628 17556 41916
rect 17612 41748 17668 42924
rect 17948 42754 18004 42766
rect 17948 42702 17950 42754
rect 18002 42702 18004 42754
rect 17836 42642 17892 42654
rect 17836 42590 17838 42642
rect 17890 42590 17892 42642
rect 17724 42084 17780 42094
rect 17724 41990 17780 42028
rect 17836 41972 17892 42590
rect 17948 42644 18004 42702
rect 17948 42578 18004 42588
rect 18060 42084 18116 42924
rect 17948 41972 18004 41982
rect 17836 41970 18004 41972
rect 17836 41918 17950 41970
rect 18002 41918 18004 41970
rect 17836 41916 18004 41918
rect 17948 41906 18004 41916
rect 17612 41682 17668 41692
rect 17612 41412 17668 41422
rect 17612 41318 17668 41356
rect 17836 41076 17892 41086
rect 17612 40628 17668 40638
rect 17500 40626 17668 40628
rect 17500 40574 17614 40626
rect 17666 40574 17668 40626
rect 17500 40572 17668 40574
rect 17612 40562 17668 40572
rect 17836 40626 17892 41020
rect 17836 40574 17838 40626
rect 17890 40574 17892 40626
rect 17836 40562 17892 40574
rect 17948 40964 18004 40974
rect 17948 40514 18004 40908
rect 17948 40462 17950 40514
rect 18002 40462 18004 40514
rect 17500 39844 17556 39854
rect 17948 39844 18004 40462
rect 17500 39842 18004 39844
rect 17500 39790 17502 39842
rect 17554 39790 18004 39842
rect 17500 39788 18004 39790
rect 17500 39778 17556 39788
rect 17500 38052 17556 38062
rect 17500 37938 17556 37996
rect 17500 37886 17502 37938
rect 17554 37886 17556 37938
rect 17500 37492 17556 37886
rect 17612 37828 17668 39788
rect 17724 39618 17780 39630
rect 17724 39566 17726 39618
rect 17778 39566 17780 39618
rect 17724 39060 17780 39566
rect 17836 39396 17892 39406
rect 17836 39302 17892 39340
rect 17724 38994 17780 39004
rect 17724 38834 17780 38846
rect 17724 38782 17726 38834
rect 17778 38782 17780 38834
rect 17724 38724 17780 38782
rect 18060 38834 18116 42028
rect 18172 39732 18228 43372
rect 18284 42978 18340 43484
rect 18284 42926 18286 42978
rect 18338 42926 18340 42978
rect 18284 42914 18340 42926
rect 18396 42980 18452 42990
rect 18396 42886 18452 42924
rect 18620 42644 18676 43820
rect 18844 43652 18900 43662
rect 18844 43558 18900 43596
rect 19404 43540 19460 43550
rect 19292 43538 19460 43540
rect 19292 43486 19406 43538
rect 19458 43486 19460 43538
rect 19292 43484 19460 43486
rect 18172 39666 18228 39676
rect 18396 42532 18452 42542
rect 18060 38782 18062 38834
rect 18114 38782 18116 38834
rect 18060 38770 18116 38782
rect 18396 39618 18452 42476
rect 18508 40964 18564 40974
rect 18508 40870 18564 40908
rect 18396 39566 18398 39618
rect 18450 39566 18452 39618
rect 18396 38668 18452 39566
rect 18620 39508 18676 42588
rect 18732 43092 18788 43102
rect 18732 41076 18788 43036
rect 18956 42980 19012 42990
rect 18956 42886 19012 42924
rect 19180 42756 19236 42766
rect 19180 42662 19236 42700
rect 19292 42308 19348 43484
rect 19404 43474 19460 43484
rect 19404 43092 19460 43102
rect 19404 42866 19460 43036
rect 19404 42814 19406 42866
rect 19458 42814 19460 42866
rect 19404 42802 19460 42814
rect 19516 42868 19572 44716
rect 19852 44212 19908 44222
rect 19628 44210 19908 44212
rect 19628 44158 19854 44210
rect 19906 44158 19908 44210
rect 19628 44156 19908 44158
rect 19628 42980 19684 44156
rect 19852 44146 19908 44156
rect 20076 44210 20132 45276
rect 20188 44548 20244 44558
rect 20188 44454 20244 44492
rect 20076 44158 20078 44210
rect 20130 44158 20132 44210
rect 20076 44146 20132 44158
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19740 43764 19796 43774
rect 20300 43708 20356 46060
rect 20412 46114 20468 46622
rect 20412 46062 20414 46114
rect 20466 46062 20468 46114
rect 20412 46050 20468 46062
rect 20636 46676 20692 48078
rect 20524 45780 20580 45818
rect 20636 45780 20692 46620
rect 20580 45724 20692 45780
rect 20748 45778 20804 48750
rect 20860 49700 20916 49710
rect 20972 49700 21028 51548
rect 20860 49698 21028 49700
rect 20860 49646 20862 49698
rect 20914 49646 21028 49698
rect 20860 49644 21028 49646
rect 20860 48356 20916 49644
rect 21084 49252 21140 49262
rect 20860 48290 20916 48300
rect 20972 48580 21028 48590
rect 20748 45726 20750 45778
rect 20802 45726 20804 45778
rect 20524 45714 20580 45724
rect 20748 45556 20804 45726
rect 20748 45490 20804 45500
rect 20860 47796 20916 47806
rect 20636 45330 20692 45342
rect 20636 45278 20638 45330
rect 20690 45278 20692 45330
rect 20636 45108 20692 45278
rect 20636 45042 20692 45052
rect 20748 45108 20804 45118
rect 20860 45108 20916 47740
rect 20972 46564 21028 48524
rect 21084 47684 21140 49196
rect 21196 47796 21252 52668
rect 21420 51828 21476 52780
rect 21420 51762 21476 51772
rect 21308 51604 21364 51614
rect 21308 50484 21364 51548
rect 21308 50418 21364 50428
rect 21532 50820 21588 50830
rect 21532 49810 21588 50764
rect 21644 50596 21700 53452
rect 21868 53442 21924 53452
rect 21980 53506 22148 53508
rect 21980 53454 22094 53506
rect 22146 53454 22148 53506
rect 21980 53452 22148 53454
rect 21980 52946 22036 53452
rect 22092 53442 22148 53452
rect 21980 52894 21982 52946
rect 22034 52894 22036 52946
rect 21980 52882 22036 52894
rect 22204 52948 22260 52958
rect 22316 52948 22372 54348
rect 22764 54338 22820 54348
rect 23100 53844 23156 55134
rect 23436 55188 23492 55198
rect 23212 55076 23268 55086
rect 23212 54982 23268 55020
rect 23324 55074 23380 55086
rect 23324 55022 23326 55074
rect 23378 55022 23380 55074
rect 23324 54964 23380 55022
rect 23324 54898 23380 54908
rect 23436 54290 23492 55132
rect 23548 54738 23604 55356
rect 23884 55300 23940 55310
rect 23548 54686 23550 54738
rect 23602 54686 23604 54738
rect 23548 54674 23604 54686
rect 23660 54852 23716 54862
rect 23660 54738 23716 54796
rect 23660 54686 23662 54738
rect 23714 54686 23716 54738
rect 23660 54674 23716 54686
rect 23436 54238 23438 54290
rect 23490 54238 23492 54290
rect 23436 53956 23492 54238
rect 23436 53890 23492 53900
rect 23100 53778 23156 53788
rect 22652 53730 22708 53742
rect 22652 53678 22654 53730
rect 22706 53678 22708 53730
rect 22204 52946 22372 52948
rect 22204 52894 22206 52946
rect 22258 52894 22372 52946
rect 22204 52892 22372 52894
rect 22428 53620 22484 53630
rect 21756 51938 21812 51950
rect 21756 51886 21758 51938
rect 21810 51886 21812 51938
rect 21756 51828 21812 51886
rect 21756 51762 21812 51772
rect 22092 51940 22148 51950
rect 22092 51378 22148 51884
rect 22092 51326 22094 51378
rect 22146 51326 22148 51378
rect 22092 51314 22148 51326
rect 21868 51268 21924 51278
rect 21868 51174 21924 51212
rect 21644 50530 21700 50540
rect 21756 50932 21812 50942
rect 21532 49758 21534 49810
rect 21586 49758 21588 49810
rect 21420 49476 21476 49486
rect 21420 49250 21476 49420
rect 21420 49198 21422 49250
rect 21474 49198 21476 49250
rect 21420 49186 21476 49198
rect 21532 49140 21588 49758
rect 21532 49074 21588 49084
rect 21756 50034 21812 50876
rect 21756 49982 21758 50034
rect 21810 49982 21812 50034
rect 21644 48802 21700 48814
rect 21644 48750 21646 48802
rect 21698 48750 21700 48802
rect 21644 48468 21700 48750
rect 21644 48402 21700 48412
rect 21756 48356 21812 49982
rect 21980 50370 22036 50382
rect 21980 50318 21982 50370
rect 22034 50318 22036 50370
rect 21980 49812 22036 50318
rect 21980 49746 22036 49756
rect 22204 49476 22260 52892
rect 22428 52836 22484 53564
rect 22540 53172 22596 53182
rect 22652 53172 22708 53678
rect 23436 53620 23492 53630
rect 22764 53508 22820 53518
rect 22764 53414 22820 53452
rect 22988 53506 23044 53518
rect 22988 53454 22990 53506
rect 23042 53454 23044 53506
rect 22988 53396 23044 53454
rect 22988 53330 23044 53340
rect 22540 53170 22708 53172
rect 22540 53118 22542 53170
rect 22594 53118 22708 53170
rect 22540 53116 22708 53118
rect 22540 53106 22596 53116
rect 22316 52612 22372 52622
rect 22316 52050 22372 52556
rect 22428 52164 22484 52780
rect 23100 52836 23156 52846
rect 23100 52742 23156 52780
rect 23324 52836 23380 52846
rect 22540 52164 22596 52174
rect 22428 52162 22596 52164
rect 22428 52110 22542 52162
rect 22594 52110 22596 52162
rect 22428 52108 22596 52110
rect 22316 51998 22318 52050
rect 22370 51998 22372 52050
rect 22316 50820 22372 51998
rect 22540 51602 22596 52108
rect 22876 52052 22932 52062
rect 22876 51958 22932 51996
rect 22764 51938 22820 51950
rect 22764 51886 22766 51938
rect 22818 51886 22820 51938
rect 22764 51828 22820 51886
rect 22764 51762 22820 51772
rect 23324 51938 23380 52780
rect 23324 51886 23326 51938
rect 23378 51886 23380 51938
rect 22540 51550 22542 51602
rect 22594 51550 22596 51602
rect 22428 51380 22484 51390
rect 22428 51286 22484 51324
rect 22316 50754 22372 50764
rect 22540 50708 22596 51550
rect 22764 51378 22820 51390
rect 22764 51326 22766 51378
rect 22818 51326 22820 51378
rect 22652 51268 22708 51278
rect 22652 51174 22708 51212
rect 22764 50932 22820 51326
rect 22764 50866 22820 50876
rect 23212 51380 23268 51390
rect 22428 50652 22596 50708
rect 22316 50596 22372 50606
rect 22428 50596 22484 50652
rect 22316 50594 22484 50596
rect 22316 50542 22318 50594
rect 22370 50542 22484 50594
rect 22316 50540 22484 50542
rect 22316 50036 22372 50540
rect 22876 50484 22932 50494
rect 22876 50390 22932 50428
rect 23212 50370 23268 51324
rect 23324 51156 23380 51886
rect 23436 51828 23492 53564
rect 23548 53172 23604 53182
rect 23548 53078 23604 53116
rect 23548 52276 23604 52286
rect 23548 52182 23604 52220
rect 23660 52164 23716 52174
rect 23660 52050 23716 52108
rect 23660 51998 23662 52050
rect 23714 51998 23716 52050
rect 23660 51986 23716 51998
rect 23436 51490 23492 51772
rect 23436 51438 23438 51490
rect 23490 51438 23492 51490
rect 23436 51426 23492 51438
rect 23548 51938 23604 51950
rect 23548 51886 23550 51938
rect 23602 51886 23604 51938
rect 23548 51380 23604 51886
rect 23772 51940 23828 51950
rect 23772 51602 23828 51884
rect 23772 51550 23774 51602
rect 23826 51550 23828 51602
rect 23772 51538 23828 51550
rect 23884 51604 23940 55244
rect 24220 55300 24276 55310
rect 24220 55206 24276 55244
rect 23996 55074 24052 55086
rect 23996 55022 23998 55074
rect 24050 55022 24052 55074
rect 23996 54516 24052 55022
rect 24444 54852 24500 56028
rect 25676 56084 25732 56094
rect 25676 55990 25732 56028
rect 25340 55970 25396 55982
rect 25340 55918 25342 55970
rect 25394 55918 25396 55970
rect 24892 55860 24948 55870
rect 24892 55298 24948 55804
rect 24892 55246 24894 55298
rect 24946 55246 24948 55298
rect 24892 55234 24948 55246
rect 25228 55300 25284 55310
rect 25228 55206 25284 55244
rect 25340 55188 25396 55918
rect 25788 55972 25844 55982
rect 25788 55410 25844 55916
rect 25788 55358 25790 55410
rect 25842 55358 25844 55410
rect 25788 55346 25844 55358
rect 25900 55860 25956 57148
rect 26460 56308 26516 56318
rect 26124 56196 26180 56206
rect 26124 56102 26180 56140
rect 25900 55804 26404 55860
rect 25900 55188 25956 55804
rect 25340 55122 25396 55132
rect 25788 55132 25956 55188
rect 26012 55636 26068 55646
rect 23996 54450 24052 54460
rect 24332 54796 24500 54852
rect 25004 55074 25060 55086
rect 25676 55076 25732 55086
rect 25004 55022 25006 55074
rect 25058 55022 25060 55074
rect 24108 53732 24164 53742
rect 23996 53620 24052 53630
rect 23996 53526 24052 53564
rect 23996 53172 24052 53182
rect 23996 51604 24052 53116
rect 24108 52500 24164 53676
rect 24108 52434 24164 52444
rect 24108 52164 24164 52174
rect 24108 52070 24164 52108
rect 23996 51548 24164 51604
rect 23884 51538 23940 51548
rect 23660 51492 23716 51502
rect 23660 51398 23716 51436
rect 23548 51314 23604 51324
rect 23884 51380 23940 51390
rect 23324 51090 23380 51100
rect 23212 50318 23214 50370
rect 23266 50318 23268 50370
rect 23212 50260 23268 50318
rect 23212 50194 23268 50204
rect 23436 50932 23492 50942
rect 22316 49904 22372 49980
rect 23324 50036 23380 50046
rect 23324 49942 23380 49980
rect 23212 49924 23268 49934
rect 23212 49830 23268 49868
rect 22652 49812 22708 49822
rect 22652 49718 22708 49756
rect 23324 49586 23380 49598
rect 23324 49534 23326 49586
rect 23378 49534 23380 49586
rect 22204 49410 22260 49420
rect 22876 49476 22932 49486
rect 22204 49252 22260 49262
rect 22204 49158 22260 49196
rect 22652 48916 22708 48926
rect 22092 48802 22148 48814
rect 22092 48750 22094 48802
rect 22146 48750 22148 48802
rect 22092 48468 22148 48750
rect 22540 48804 22596 48814
rect 22540 48710 22596 48748
rect 22092 48402 22148 48412
rect 21756 48290 21812 48300
rect 21196 47730 21252 47740
rect 21308 48130 21364 48142
rect 21308 48078 21310 48130
rect 21362 48078 21364 48130
rect 21308 47908 21364 48078
rect 21084 46898 21140 47628
rect 21084 46846 21086 46898
rect 21138 46846 21140 46898
rect 21084 46834 21140 46846
rect 21308 46900 21364 47852
rect 21644 48132 21700 48142
rect 21644 47346 21700 48076
rect 21644 47294 21646 47346
rect 21698 47294 21700 47346
rect 21644 47282 21700 47294
rect 21868 48130 21924 48142
rect 22316 48132 22372 48142
rect 21868 48078 21870 48130
rect 21922 48078 21924 48130
rect 21868 47012 21924 48078
rect 21980 48130 22372 48132
rect 21980 48078 22318 48130
rect 22370 48078 22372 48130
rect 21980 48076 22372 48078
rect 21980 47460 22036 48076
rect 22316 48066 22372 48076
rect 22540 47684 22596 47694
rect 22540 47590 22596 47628
rect 21980 47458 22148 47460
rect 21980 47406 21982 47458
rect 22034 47406 22148 47458
rect 21980 47404 22148 47406
rect 21980 47394 22036 47404
rect 21868 46946 21924 46956
rect 21308 46834 21364 46844
rect 20972 46498 21028 46508
rect 21420 46562 21476 46574
rect 21420 46510 21422 46562
rect 21474 46510 21476 46562
rect 20748 45106 20916 45108
rect 20748 45054 20750 45106
rect 20802 45054 20916 45106
rect 20748 45052 20916 45054
rect 20748 45042 20804 45052
rect 20524 44884 20580 44894
rect 20524 44100 20580 44828
rect 20636 44100 20692 44110
rect 20524 44098 20692 44100
rect 20524 44046 20638 44098
rect 20690 44046 20692 44098
rect 20524 44044 20692 44046
rect 19740 43538 19796 43708
rect 19740 43486 19742 43538
rect 19794 43486 19796 43538
rect 19740 43474 19796 43486
rect 19964 43650 20020 43662
rect 19964 43598 19966 43650
rect 20018 43598 20020 43650
rect 19964 43540 20020 43598
rect 20188 43652 20356 43708
rect 20412 43876 20468 43886
rect 20188 43650 20244 43652
rect 20188 43598 20190 43650
rect 20242 43598 20244 43650
rect 20188 43586 20244 43598
rect 19964 43474 20020 43484
rect 20300 43540 20356 43550
rect 20076 43426 20132 43438
rect 20076 43374 20078 43426
rect 20130 43374 20132 43426
rect 19628 42914 19684 42924
rect 19852 43204 19908 43214
rect 19516 42532 19572 42812
rect 19740 42868 19796 42878
rect 19740 42774 19796 42812
rect 19852 42754 19908 43148
rect 19852 42702 19854 42754
rect 19906 42702 19908 42754
rect 19852 42690 19908 42702
rect 20076 42644 20132 43374
rect 20076 42578 20132 42588
rect 19628 42532 19684 42542
rect 19516 42530 19684 42532
rect 19516 42478 19630 42530
rect 19682 42478 19684 42530
rect 19516 42476 19684 42478
rect 19292 42242 19348 42252
rect 18844 41972 18900 41982
rect 18844 41878 18900 41916
rect 19068 41972 19124 41982
rect 18956 41858 19012 41870
rect 18956 41806 18958 41858
rect 19010 41806 19012 41858
rect 18956 41412 19012 41806
rect 19068 41746 19124 41916
rect 19068 41694 19070 41746
rect 19122 41694 19124 41746
rect 19068 41682 19124 41694
rect 18956 41346 19012 41356
rect 18844 41076 18900 41086
rect 18732 41074 18900 41076
rect 18732 41022 18846 41074
rect 18898 41022 18900 41074
rect 18732 41020 18900 41022
rect 18844 41010 18900 41020
rect 19292 41076 19348 41086
rect 19516 41076 19572 41086
rect 19292 41074 19516 41076
rect 19292 41022 19294 41074
rect 19346 41022 19516 41074
rect 19292 41020 19516 41022
rect 19292 41010 19348 41020
rect 19516 41010 19572 41020
rect 19628 40964 19684 42476
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19964 41858 20020 41870
rect 19964 41806 19966 41858
rect 20018 41806 20020 41858
rect 19852 41524 19908 41534
rect 19852 41410 19908 41468
rect 19852 41358 19854 41410
rect 19906 41358 19908 41410
rect 19852 41346 19908 41358
rect 19964 41412 20020 41806
rect 20300 41860 20356 43484
rect 20300 41766 20356 41804
rect 20412 43316 20468 43820
rect 19964 41346 20020 41356
rect 20076 41188 20132 41198
rect 20412 41188 20468 43260
rect 20524 43092 20580 44044
rect 20636 44034 20692 44044
rect 20636 43652 20692 43662
rect 20636 43558 20692 43596
rect 20524 43026 20580 43036
rect 20860 42868 20916 45052
rect 21308 45106 21364 45118
rect 21308 45054 21310 45106
rect 21362 45054 21364 45106
rect 21308 44548 21364 45054
rect 21308 44482 21364 44492
rect 21308 43988 21364 43998
rect 21084 43428 21140 43438
rect 21084 43334 21140 43372
rect 20860 42866 21140 42868
rect 20860 42814 20862 42866
rect 20914 42814 21140 42866
rect 20860 42812 21140 42814
rect 20860 42802 20916 42812
rect 20524 42530 20580 42542
rect 20524 42478 20526 42530
rect 20578 42478 20580 42530
rect 20524 41636 20580 42478
rect 20748 41858 20804 41870
rect 20748 41806 20750 41858
rect 20802 41806 20804 41858
rect 20748 41748 20804 41806
rect 20804 41692 20916 41748
rect 20748 41682 20804 41692
rect 20524 41570 20580 41580
rect 20748 41412 20804 41422
rect 20636 41300 20692 41310
rect 20636 41206 20692 41244
rect 20076 41186 20244 41188
rect 20076 41134 20078 41186
rect 20130 41134 20244 41186
rect 20076 41132 20244 41134
rect 20076 41122 20132 41132
rect 19740 40964 19796 40974
rect 19628 40908 19740 40964
rect 19740 40898 19796 40908
rect 19516 40852 19572 40862
rect 19068 40402 19124 40414
rect 19068 40350 19070 40402
rect 19122 40350 19124 40402
rect 18732 40292 18788 40302
rect 19068 40292 19124 40350
rect 19516 40292 19572 40796
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 20188 40628 20244 41132
rect 20412 41056 20468 41132
rect 20748 41186 20804 41356
rect 20748 41134 20750 41186
rect 20802 41134 20804 41186
rect 20748 41122 20804 41134
rect 20524 40962 20580 40974
rect 20524 40910 20526 40962
rect 20578 40910 20580 40962
rect 20412 40628 20468 40638
rect 20188 40626 20468 40628
rect 20188 40574 20414 40626
rect 20466 40574 20468 40626
rect 20188 40572 20468 40574
rect 20412 40562 20468 40572
rect 20076 40516 20132 40526
rect 20076 40422 20132 40460
rect 20412 40404 20468 40414
rect 20412 40310 20468 40348
rect 18732 40290 18900 40292
rect 18732 40238 18734 40290
rect 18786 40238 18900 40290
rect 18732 40236 18900 40238
rect 18732 40226 18788 40236
rect 18732 39508 18788 39518
rect 18620 39506 18788 39508
rect 18620 39454 18734 39506
rect 18786 39454 18788 39506
rect 18620 39452 18788 39454
rect 18732 39442 18788 39452
rect 17724 38658 17780 38668
rect 18284 38612 18452 38668
rect 18620 39172 18676 39182
rect 17836 37828 17892 37838
rect 17612 37826 17892 37828
rect 17612 37774 17838 37826
rect 17890 37774 17892 37826
rect 17612 37772 17892 37774
rect 17500 37426 17556 37436
rect 17836 37268 17892 37772
rect 17836 37202 17892 37212
rect 17724 37154 17780 37166
rect 17724 37102 17726 37154
rect 17778 37102 17780 37154
rect 17724 36820 17780 37102
rect 17724 36754 17780 36764
rect 17724 36596 17780 36606
rect 17724 36258 17780 36540
rect 18284 36484 18340 38612
rect 18620 38162 18676 39116
rect 18620 38110 18622 38162
rect 18674 38110 18676 38162
rect 18620 38098 18676 38110
rect 18732 38164 18788 38174
rect 18732 38070 18788 38108
rect 18508 37828 18564 37838
rect 18844 37828 18900 40236
rect 19068 40226 19124 40236
rect 19404 40290 19572 40292
rect 19404 40238 19518 40290
rect 19570 40238 19572 40290
rect 19404 40236 19572 40238
rect 19068 38276 19124 38286
rect 18508 37826 18900 37828
rect 18508 37774 18510 37826
rect 18562 37774 18900 37826
rect 18508 37772 18900 37774
rect 18956 37828 19012 37838
rect 18508 37762 18564 37772
rect 18396 37268 18452 37278
rect 18620 37268 18676 37278
rect 18396 37266 18564 37268
rect 18396 37214 18398 37266
rect 18450 37214 18564 37266
rect 18396 37212 18564 37214
rect 18396 37202 18452 37212
rect 18508 37044 18564 37212
rect 18620 37174 18676 37212
rect 18508 36988 18676 37044
rect 18284 36428 18452 36484
rect 18172 36260 18228 36270
rect 17724 36206 17726 36258
rect 17778 36206 17780 36258
rect 17724 36194 17780 36206
rect 17836 36258 18228 36260
rect 17836 36206 18174 36258
rect 18226 36206 18228 36258
rect 17836 36204 18228 36206
rect 17388 36082 17444 36092
rect 17276 35858 17332 35868
rect 17724 35812 17780 35822
rect 17724 35718 17780 35756
rect 17836 35588 17892 36204
rect 18172 36194 18228 36204
rect 18284 36260 18340 36270
rect 17276 35532 17892 35588
rect 17276 33570 17332 35532
rect 17276 33518 17278 33570
rect 17330 33518 17332 33570
rect 17276 33506 17332 33518
rect 17500 35364 17556 35374
rect 17500 34802 17556 35308
rect 17836 34914 17892 35532
rect 17836 34862 17838 34914
rect 17890 34862 17892 34914
rect 17836 34850 17892 34862
rect 18172 35700 18228 35710
rect 17500 34750 17502 34802
rect 17554 34750 17556 34802
rect 17388 33236 17444 33246
rect 17052 31890 17220 31892
rect 17052 31838 17054 31890
rect 17106 31838 17220 31890
rect 17052 31836 17220 31838
rect 17276 32676 17332 32686
rect 17052 31826 17108 31836
rect 16380 30996 16436 31006
rect 16044 30884 16100 30894
rect 16044 30790 16100 30828
rect 15820 29698 15876 29708
rect 16268 30210 16324 30222
rect 16268 30158 16270 30210
rect 16322 30158 16324 30210
rect 15372 29538 15428 29550
rect 15372 29486 15374 29538
rect 15426 29486 15428 29538
rect 15372 28644 15428 29486
rect 16268 29540 16324 30158
rect 16268 29474 16324 29484
rect 16380 30212 16436 30940
rect 16940 30436 16996 31724
rect 16940 30370 16996 30380
rect 15596 29428 15652 29438
rect 15596 29334 15652 29372
rect 16268 29316 16324 29326
rect 16380 29316 16436 30156
rect 16828 30324 16884 30334
rect 17276 30324 17332 32620
rect 17388 32116 17444 33180
rect 17388 32050 17444 32060
rect 17500 31220 17556 34750
rect 17948 34244 18004 34254
rect 17948 34150 18004 34188
rect 17612 33348 17668 33358
rect 17612 33236 17668 33292
rect 17836 33236 17892 33246
rect 17612 33234 17892 33236
rect 17612 33182 17838 33234
rect 17890 33182 17892 33234
rect 17612 33180 17892 33182
rect 17612 32786 17668 33180
rect 17836 33170 17892 33180
rect 18172 33234 18228 35644
rect 18284 35698 18340 36204
rect 18284 35646 18286 35698
rect 18338 35646 18340 35698
rect 18284 35634 18340 35646
rect 18396 35364 18452 36428
rect 18508 36372 18564 36382
rect 18508 36278 18564 36316
rect 18620 36036 18676 36988
rect 18396 35298 18452 35308
rect 18508 35980 18676 36036
rect 18284 34914 18340 34926
rect 18284 34862 18286 34914
rect 18338 34862 18340 34914
rect 18284 34356 18340 34862
rect 18396 34804 18452 34814
rect 18396 34710 18452 34748
rect 18508 34690 18564 35980
rect 18732 35252 18788 37772
rect 18844 37154 18900 37166
rect 18844 37102 18846 37154
rect 18898 37102 18900 37154
rect 18844 36036 18900 37102
rect 18844 35970 18900 35980
rect 18732 35186 18788 35196
rect 18844 35700 18900 35710
rect 18508 34638 18510 34690
rect 18562 34638 18564 34690
rect 18508 34626 18564 34638
rect 18284 34290 18340 34300
rect 18732 34580 18788 34590
rect 18620 34244 18676 34254
rect 18620 34150 18676 34188
rect 18732 34242 18788 34524
rect 18732 34190 18734 34242
rect 18786 34190 18788 34242
rect 18732 33458 18788 34190
rect 18844 34242 18900 35644
rect 18956 35698 19012 37772
rect 19068 37042 19124 38220
rect 19292 37940 19348 37950
rect 19292 37846 19348 37884
rect 19404 37268 19460 40236
rect 19516 40226 19572 40236
rect 20524 40180 20580 40910
rect 20524 40114 20580 40124
rect 20636 40402 20692 40414
rect 20636 40350 20638 40402
rect 20690 40350 20692 40402
rect 19404 37202 19460 37212
rect 19516 40068 19572 40078
rect 19068 36990 19070 37042
rect 19122 36990 19124 37042
rect 19068 36978 19124 36990
rect 19068 36260 19124 36270
rect 19068 35812 19124 36204
rect 19068 35746 19124 35756
rect 18956 35646 18958 35698
rect 19010 35646 19012 35698
rect 18956 35634 19012 35646
rect 19292 35698 19348 35710
rect 19292 35646 19294 35698
rect 19346 35646 19348 35698
rect 19180 35588 19236 35598
rect 19180 34914 19236 35532
rect 19180 34862 19182 34914
rect 19234 34862 19236 34914
rect 19180 34850 19236 34862
rect 19292 34580 19348 35646
rect 19404 35700 19460 35710
rect 19404 35606 19460 35644
rect 19292 34514 19348 34524
rect 19292 34356 19348 34366
rect 19516 34356 19572 40012
rect 20636 39956 20692 40350
rect 20860 40404 20916 41692
rect 20860 40338 20916 40348
rect 20972 41746 21028 41758
rect 20972 41694 20974 41746
rect 21026 41694 21028 41746
rect 20188 39900 20692 39956
rect 20972 40292 21028 41694
rect 21084 41524 21140 42812
rect 21308 42084 21364 43932
rect 21420 43764 21476 46510
rect 21868 46114 21924 46126
rect 21868 46062 21870 46114
rect 21922 46062 21924 46114
rect 21868 46002 21924 46062
rect 21868 45950 21870 46002
rect 21922 45950 21924 46002
rect 21868 45938 21924 45950
rect 21532 45332 21588 45342
rect 21532 45238 21588 45276
rect 21868 45220 21924 45230
rect 21868 45126 21924 45164
rect 21756 45106 21812 45118
rect 21756 45054 21758 45106
rect 21810 45054 21812 45106
rect 21420 43698 21476 43708
rect 21644 44994 21700 45006
rect 21644 44942 21646 44994
rect 21698 44942 21700 44994
rect 21532 43540 21588 43550
rect 21532 43446 21588 43484
rect 21644 43316 21700 44942
rect 21756 44324 21812 45054
rect 22092 44436 22148 47404
rect 22540 46900 22596 46910
rect 22540 46806 22596 46844
rect 22204 46564 22260 46574
rect 22204 46562 22484 46564
rect 22204 46510 22206 46562
rect 22258 46510 22484 46562
rect 22204 46508 22484 46510
rect 22204 46114 22260 46508
rect 22204 46062 22206 46114
rect 22258 46062 22260 46114
rect 22204 46050 22260 46062
rect 22428 45778 22484 46508
rect 22428 45726 22430 45778
rect 22482 45726 22484 45778
rect 22428 45220 22484 45726
rect 22092 44380 22260 44436
rect 21868 44324 21924 44334
rect 21756 44268 21868 44324
rect 21868 44230 21924 44268
rect 21980 44210 22036 44222
rect 21980 44158 21982 44210
rect 22034 44158 22036 44210
rect 21980 43764 22036 44158
rect 22092 44210 22148 44222
rect 22092 44158 22094 44210
rect 22146 44158 22148 44210
rect 22092 44100 22148 44158
rect 22092 44034 22148 44044
rect 21980 43698 22036 43708
rect 22092 43652 22148 43662
rect 22092 43558 22148 43596
rect 21644 43250 21700 43260
rect 21532 43204 21588 43214
rect 21420 42084 21476 42094
rect 21308 42028 21420 42084
rect 21196 41860 21252 41870
rect 21196 41766 21252 41804
rect 21084 41458 21140 41468
rect 21308 41524 21364 41534
rect 20972 39956 21028 40236
rect 19852 39844 19908 39854
rect 19852 39750 19908 39788
rect 20188 39842 20244 39900
rect 20972 39890 21028 39900
rect 20188 39790 20190 39842
rect 20242 39790 20244 39842
rect 20188 39778 20244 39790
rect 19628 39508 19684 39546
rect 19628 39442 19684 39452
rect 20972 39394 21028 39406
rect 20972 39342 20974 39394
rect 21026 39342 21028 39394
rect 19628 39284 19684 39294
rect 19628 38834 19684 39228
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 20972 38948 21028 39342
rect 19628 38782 19630 38834
rect 19682 38782 19684 38834
rect 19628 38770 19684 38782
rect 20748 38836 20804 38846
rect 20748 38742 20804 38780
rect 20636 38724 20692 38734
rect 20300 38164 20356 38174
rect 20300 38050 20356 38108
rect 20636 38162 20692 38668
rect 20636 38110 20638 38162
rect 20690 38110 20692 38162
rect 20636 38098 20692 38110
rect 20300 37998 20302 38050
rect 20354 37998 20356 38050
rect 20300 37986 20356 37998
rect 19628 37940 19684 37950
rect 19628 37846 19684 37884
rect 20636 37940 20692 37950
rect 19628 37716 19684 37726
rect 19628 37154 19684 37660
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20636 37380 20692 37884
rect 20860 37940 20916 37950
rect 20860 37846 20916 37884
rect 20076 37268 20132 37278
rect 20076 37174 20132 37212
rect 19628 37102 19630 37154
rect 19682 37102 19684 37154
rect 19628 37090 19684 37102
rect 19852 36820 19908 36830
rect 19852 36482 19908 36764
rect 19852 36430 19854 36482
rect 19906 36430 19908 36482
rect 19628 36372 19684 36382
rect 19628 36278 19684 36316
rect 19852 36260 19908 36430
rect 19852 36194 19908 36204
rect 20524 36370 20580 36382
rect 20524 36318 20526 36370
rect 20578 36318 20580 36370
rect 20524 36260 20580 36318
rect 20524 36194 20580 36204
rect 20636 36258 20692 37324
rect 20972 36596 21028 38892
rect 21308 38668 21364 41468
rect 21420 40626 21476 42028
rect 21420 40574 21422 40626
rect 21474 40574 21476 40626
rect 21420 40404 21476 40574
rect 21420 40338 21476 40348
rect 20972 36530 21028 36540
rect 21196 38612 21364 38668
rect 21420 39956 21476 39966
rect 21420 39732 21476 39900
rect 21420 38724 21476 39676
rect 21420 38658 21476 38668
rect 20636 36206 20638 36258
rect 20690 36206 20692 36258
rect 19292 34354 19572 34356
rect 19292 34302 19294 34354
rect 19346 34302 19572 34354
rect 19292 34300 19572 34302
rect 19628 36148 19684 36158
rect 19292 34290 19348 34300
rect 18844 34190 18846 34242
rect 18898 34190 18900 34242
rect 18844 34178 18900 34190
rect 18732 33406 18734 33458
rect 18786 33406 18788 33458
rect 18732 33394 18788 33406
rect 18172 33182 18174 33234
rect 18226 33182 18228 33234
rect 18172 33170 18228 33182
rect 19292 33124 19348 33134
rect 19628 33124 19684 36092
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 20636 35810 20692 36206
rect 20860 36260 20916 36270
rect 20860 36166 20916 36204
rect 20636 35758 20638 35810
rect 20690 35758 20692 35810
rect 20636 35700 20692 35758
rect 20860 35700 20916 35710
rect 20076 35644 20692 35700
rect 20748 35698 20916 35700
rect 20748 35646 20862 35698
rect 20914 35646 20916 35698
rect 20748 35644 20916 35646
rect 19964 35476 20020 35486
rect 19964 35382 20020 35420
rect 20076 34804 20132 35644
rect 20076 34738 20132 34748
rect 20524 35252 20580 35262
rect 20524 34802 20580 35196
rect 20524 34750 20526 34802
rect 20578 34750 20580 34802
rect 20524 34738 20580 34750
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19740 34132 19796 34142
rect 19740 34038 19796 34076
rect 20188 34132 20244 34142
rect 19292 33122 19684 33124
rect 19292 33070 19294 33122
rect 19346 33070 19684 33122
rect 19292 33068 19684 33070
rect 20188 34018 20244 34076
rect 20748 34130 20804 35644
rect 20860 35634 20916 35644
rect 21084 35252 21140 35262
rect 20860 34916 20916 34926
rect 21084 34916 21140 35196
rect 20860 34914 21140 34916
rect 20860 34862 20862 34914
rect 20914 34862 21140 34914
rect 20860 34860 21140 34862
rect 20860 34850 20916 34860
rect 21084 34354 21140 34860
rect 21084 34302 21086 34354
rect 21138 34302 21140 34354
rect 21084 34290 21140 34302
rect 20748 34078 20750 34130
rect 20802 34078 20804 34130
rect 20188 33966 20190 34018
rect 20242 33966 20244 34018
rect 19292 32900 19348 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19292 32834 19348 32844
rect 17612 32734 17614 32786
rect 17666 32734 17668 32786
rect 17612 32452 17668 32734
rect 18172 32788 18228 32798
rect 18172 32694 18228 32732
rect 18956 32788 19012 32798
rect 18956 32562 19012 32732
rect 18956 32510 18958 32562
rect 19010 32510 19012 32562
rect 18956 32498 19012 32510
rect 19516 32564 19572 32574
rect 19516 32470 19572 32508
rect 17612 32386 17668 32396
rect 19628 32450 19684 32462
rect 19628 32398 19630 32450
rect 19682 32398 19684 32450
rect 19516 32004 19572 32014
rect 19628 32004 19684 32398
rect 20188 32340 20244 33966
rect 20412 34020 20468 34030
rect 20412 33458 20468 33964
rect 20748 34020 20804 34078
rect 20748 33954 20804 33964
rect 20412 33406 20414 33458
rect 20466 33406 20468 33458
rect 20412 33394 20468 33406
rect 20188 32274 20244 32284
rect 20860 33122 20916 33134
rect 20860 33070 20862 33122
rect 20914 33070 20916 33122
rect 20860 32340 20916 33070
rect 20860 32274 20916 32284
rect 19516 32002 19684 32004
rect 19516 31950 19518 32002
rect 19570 31950 19684 32002
rect 19516 31948 19684 31950
rect 19516 31938 19572 31948
rect 20300 31892 20356 31902
rect 19852 31780 19908 31790
rect 19852 31686 19908 31724
rect 19628 31556 19684 31566
rect 18844 31554 19684 31556
rect 18844 31502 19630 31554
rect 19682 31502 19684 31554
rect 18844 31500 19684 31502
rect 17612 31220 17668 31230
rect 17500 31218 18004 31220
rect 17500 31166 17614 31218
rect 17666 31166 18004 31218
rect 17500 31164 18004 31166
rect 17612 31154 17668 31164
rect 16828 29652 16884 30268
rect 17052 30268 17332 30324
rect 17724 30436 17780 30446
rect 16940 30212 16996 30222
rect 16940 30118 16996 30156
rect 16940 29652 16996 29662
rect 16828 29650 16996 29652
rect 16828 29598 16942 29650
rect 16994 29598 16996 29650
rect 16828 29596 16996 29598
rect 16940 29586 16996 29596
rect 17052 29428 17108 30268
rect 16268 29314 16436 29316
rect 16268 29262 16270 29314
rect 16322 29262 16436 29314
rect 16268 29260 16436 29262
rect 16828 29372 17108 29428
rect 17164 30098 17220 30110
rect 17164 30046 17166 30098
rect 17218 30046 17220 30098
rect 16268 29250 16324 29260
rect 15372 28578 15428 28588
rect 16044 28980 16100 28990
rect 15484 28084 15540 28094
rect 15484 27990 15540 28028
rect 15820 27746 15876 27758
rect 15820 27694 15822 27746
rect 15874 27694 15876 27746
rect 15820 27412 15876 27694
rect 15820 27346 15876 27356
rect 16044 25620 16100 28924
rect 16604 28642 16660 28654
rect 16604 28590 16606 28642
rect 16658 28590 16660 28642
rect 16268 27972 16324 27982
rect 16268 27748 16324 27916
rect 16604 27748 16660 28590
rect 16268 27746 16660 27748
rect 16268 27694 16270 27746
rect 16322 27694 16660 27746
rect 16268 27692 16660 27694
rect 16268 26964 16324 27692
rect 16268 26514 16324 26908
rect 16828 26908 16884 29372
rect 17164 29092 17220 30046
rect 17724 30098 17780 30380
rect 17724 30046 17726 30098
rect 17778 30046 17780 30098
rect 17724 30034 17780 30046
rect 17948 30210 18004 31164
rect 18396 30994 18452 31006
rect 18396 30942 18398 30994
rect 18450 30942 18452 30994
rect 17948 30158 17950 30210
rect 18002 30158 18004 30210
rect 17948 29876 18004 30158
rect 17948 29810 18004 29820
rect 18284 30436 18340 30446
rect 18284 29650 18340 30380
rect 18284 29598 18286 29650
rect 18338 29598 18340 29650
rect 18284 29586 18340 29598
rect 18396 29988 18452 30942
rect 18844 30994 18900 31500
rect 19628 31490 19684 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 18844 30942 18846 30994
rect 18898 30942 18900 30994
rect 18844 30930 18900 30942
rect 19180 30436 19236 30446
rect 19180 30342 19236 30380
rect 19740 30322 19796 30334
rect 19740 30270 19742 30322
rect 19794 30270 19796 30322
rect 18396 29428 18452 29932
rect 18956 30210 19012 30222
rect 18956 30158 18958 30210
rect 19010 30158 19012 30210
rect 18956 29652 19012 30158
rect 19628 30210 19684 30222
rect 19628 30158 19630 30210
rect 19682 30158 19684 30210
rect 18956 29586 19012 29596
rect 19404 30098 19460 30110
rect 19404 30046 19406 30098
rect 19458 30046 19460 30098
rect 18620 29428 18676 29438
rect 18396 29426 18676 29428
rect 18396 29374 18622 29426
rect 18674 29374 18676 29426
rect 18396 29372 18676 29374
rect 17164 29026 17220 29036
rect 17612 29314 17668 29326
rect 17612 29262 17614 29314
rect 17666 29262 17668 29314
rect 17612 29092 17668 29262
rect 17668 29036 17780 29092
rect 17612 29026 17668 29036
rect 17052 28532 17108 28542
rect 16940 28196 16996 28206
rect 16940 28082 16996 28140
rect 16940 28030 16942 28082
rect 16994 28030 16996 28082
rect 16940 28018 16996 28030
rect 16828 26852 16996 26908
rect 16268 26462 16270 26514
rect 16322 26462 16324 26514
rect 16268 26450 16324 26462
rect 15596 25618 16100 25620
rect 15596 25566 16046 25618
rect 16098 25566 16100 25618
rect 15596 25564 16100 25566
rect 15596 25506 15652 25564
rect 16044 25554 16100 25564
rect 15596 25454 15598 25506
rect 15650 25454 15652 25506
rect 15596 25442 15652 25454
rect 15260 25394 15428 25396
rect 15260 25342 15262 25394
rect 15314 25342 15428 25394
rect 15260 25340 15428 25342
rect 15260 25330 15316 25340
rect 13916 25116 14420 25172
rect 14364 24946 14420 25116
rect 14364 24894 14366 24946
rect 14418 24894 14420 24946
rect 14364 24882 14420 24894
rect 14700 24836 14756 24846
rect 14700 24742 14756 24780
rect 15260 24836 15316 24846
rect 15260 24742 15316 24780
rect 14364 24388 14420 24398
rect 14364 17666 14420 24332
rect 15372 23492 15428 25340
rect 15372 23426 15428 23436
rect 16604 20580 16660 20590
rect 16492 18450 16548 18462
rect 16492 18398 16494 18450
rect 16546 18398 16548 18450
rect 16492 17892 16548 18398
rect 16604 18452 16660 20524
rect 16940 18562 16996 26852
rect 17052 26066 17108 28476
rect 17612 28532 17668 28542
rect 17612 28418 17668 28476
rect 17612 28366 17614 28418
rect 17666 28366 17668 28418
rect 17612 28308 17668 28366
rect 17612 28242 17668 28252
rect 17724 27858 17780 29036
rect 18060 28418 18116 28430
rect 18060 28366 18062 28418
rect 18114 28366 18116 28418
rect 17724 27806 17726 27858
rect 17778 27806 17780 27858
rect 17724 27188 17780 27806
rect 17948 28196 18004 28206
rect 17948 27858 18004 28140
rect 17948 27806 17950 27858
rect 18002 27806 18004 27858
rect 17948 27794 18004 27806
rect 17724 27122 17780 27132
rect 17948 27636 18004 27646
rect 17164 26964 17220 27002
rect 17164 26898 17220 26908
rect 17052 26014 17054 26066
rect 17106 26014 17108 26066
rect 17052 22708 17108 26014
rect 17500 25506 17556 25518
rect 17500 25454 17502 25506
rect 17554 25454 17556 25506
rect 17500 25284 17556 25454
rect 17948 25506 18004 27580
rect 18060 26964 18116 28366
rect 18284 27860 18340 27870
rect 18284 27766 18340 27804
rect 18396 26908 18452 29372
rect 18620 29362 18676 29372
rect 19292 29428 19348 29438
rect 19404 29428 19460 30046
rect 19628 29540 19684 30158
rect 19740 30212 19796 30270
rect 20188 30212 20244 30222
rect 19740 30210 20244 30212
rect 19740 30158 20190 30210
rect 20242 30158 20244 30210
rect 19740 30156 20244 30158
rect 20188 30146 20244 30156
rect 20300 30100 20356 31836
rect 21084 30994 21140 31006
rect 21084 30942 21086 30994
rect 21138 30942 21140 30994
rect 20524 30884 20580 30894
rect 20524 30324 20580 30828
rect 20524 30210 20580 30268
rect 20524 30158 20526 30210
rect 20578 30158 20580 30210
rect 20524 30146 20580 30158
rect 20412 30100 20468 30110
rect 20300 30098 20468 30100
rect 20300 30046 20414 30098
rect 20466 30046 20468 30098
rect 20300 30044 20468 30046
rect 20412 30034 20468 30044
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 21084 29764 21140 30942
rect 21084 29698 21140 29708
rect 19628 29474 19684 29484
rect 19964 29652 20020 29662
rect 19292 29426 19460 29428
rect 19292 29374 19294 29426
rect 19346 29374 19460 29426
rect 19292 29372 19460 29374
rect 19292 29362 19348 29372
rect 19964 28754 20020 29596
rect 19964 28702 19966 28754
rect 20018 28702 20020 28754
rect 19964 28690 20020 28702
rect 20412 29540 20468 29550
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19180 27970 19236 27982
rect 19180 27918 19182 27970
rect 19234 27918 19236 27970
rect 18844 27860 18900 27870
rect 18844 27766 18900 27804
rect 19180 27636 19236 27918
rect 19180 27570 19236 27580
rect 18508 27188 18564 27198
rect 18508 27094 18564 27132
rect 18060 26898 18116 26908
rect 18284 26852 18452 26908
rect 20300 26964 20356 26974
rect 17948 25454 17950 25506
rect 18002 25454 18004 25506
rect 17948 25442 18004 25454
rect 18060 26402 18116 26414
rect 18060 26350 18062 26402
rect 18114 26350 18116 26402
rect 18060 25284 18116 26350
rect 18172 26068 18228 26078
rect 18172 25732 18228 26012
rect 18172 25666 18228 25676
rect 17500 25228 18116 25284
rect 18284 24612 18340 26852
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19180 26404 19236 26414
rect 18396 26292 18452 26302
rect 18396 26198 18452 26236
rect 18956 26292 19012 26302
rect 18956 26198 19012 26236
rect 18844 24836 18900 24846
rect 18844 24742 18900 24780
rect 17500 23940 17556 23950
rect 17500 23846 17556 23884
rect 17836 23938 17892 23950
rect 17836 23886 17838 23938
rect 17890 23886 17892 23938
rect 17052 22652 17332 22708
rect 16940 18510 16942 18562
rect 16994 18510 16996 18562
rect 16940 18498 16996 18510
rect 16604 18386 16660 18396
rect 16716 18338 16772 18350
rect 16716 18286 16718 18338
rect 16770 18286 16772 18338
rect 16604 17892 16660 17902
rect 16492 17890 16660 17892
rect 16492 17838 16606 17890
rect 16658 17838 16660 17890
rect 16492 17836 16660 17838
rect 15148 17780 15204 17790
rect 15148 17686 15204 17724
rect 16268 17780 16324 17818
rect 16268 17714 16324 17724
rect 14364 17614 14366 17666
rect 14418 17614 14420 17666
rect 14364 17602 14420 17614
rect 15260 17668 15316 17678
rect 15932 17668 15988 17678
rect 15260 17666 15428 17668
rect 15260 17614 15262 17666
rect 15314 17614 15428 17666
rect 15260 17612 15428 17614
rect 15260 17602 15316 17612
rect 15372 16994 15428 17612
rect 15372 16942 15374 16994
rect 15426 16942 15428 16994
rect 14812 16324 14868 16334
rect 14812 16230 14868 16268
rect 14700 15988 14756 15998
rect 14700 15894 14756 15932
rect 14812 15876 14868 15886
rect 14812 15782 14868 15820
rect 14476 15426 14532 15438
rect 14476 15374 14478 15426
rect 14530 15374 14532 15426
rect 14252 14756 14308 14766
rect 14252 14642 14308 14700
rect 14252 14590 14254 14642
rect 14306 14590 14308 14642
rect 14252 14578 14308 14590
rect 14476 14532 14532 15374
rect 13804 14420 13860 14430
rect 13804 14326 13860 14364
rect 13020 14242 13076 14252
rect 13916 13972 13972 13982
rect 13916 13878 13972 13916
rect 14476 13972 14532 14476
rect 14700 15314 14756 15326
rect 14700 15262 14702 15314
rect 14754 15262 14756 15314
rect 14700 14530 14756 15262
rect 14924 14756 14980 14766
rect 14924 14662 14980 14700
rect 14700 14478 14702 14530
rect 14754 14478 14756 14530
rect 14700 14420 14756 14478
rect 14700 14354 14756 14364
rect 14476 13746 14532 13916
rect 14924 14308 14980 14318
rect 14476 13694 14478 13746
rect 14530 13694 14532 13746
rect 14476 13682 14532 13694
rect 14700 13748 14756 13758
rect 14700 13654 14756 13692
rect 14924 13746 14980 14252
rect 15260 14306 15316 14318
rect 15260 14254 15262 14306
rect 15314 14254 15316 14306
rect 14924 13694 14926 13746
rect 14978 13694 14980 13746
rect 14924 13682 14980 13694
rect 15036 13748 15092 13758
rect 14364 13522 14420 13534
rect 14364 13470 14366 13522
rect 14418 13470 14420 13522
rect 14364 13188 14420 13470
rect 14364 13122 14420 13132
rect 15036 13074 15092 13692
rect 15260 13748 15316 14254
rect 15372 13972 15428 16942
rect 15932 16882 15988 17612
rect 15932 16830 15934 16882
rect 15986 16830 15988 16882
rect 15932 16818 15988 16830
rect 16044 17554 16100 17566
rect 16044 17502 16046 17554
rect 16098 17502 16100 17554
rect 15820 16324 15876 16334
rect 15372 13906 15428 13916
rect 15708 13970 15764 13982
rect 15708 13918 15710 13970
rect 15762 13918 15764 13970
rect 15484 13860 15540 13870
rect 15316 13692 15428 13748
rect 15260 13682 15316 13692
rect 15260 13188 15316 13198
rect 15036 13022 15038 13074
rect 15090 13022 15092 13074
rect 15036 13010 15092 13022
rect 15148 13132 15260 13188
rect 15148 12402 15204 13132
rect 15260 13094 15316 13132
rect 15148 12350 15150 12402
rect 15202 12350 15204 12402
rect 15148 12338 15204 12350
rect 15372 12402 15428 13692
rect 15484 13746 15540 13804
rect 15484 13694 15486 13746
rect 15538 13694 15540 13746
rect 15484 13188 15540 13694
rect 15484 13132 15652 13188
rect 15372 12350 15374 12402
rect 15426 12350 15428 12402
rect 15372 12338 15428 12350
rect 15484 12962 15540 12974
rect 15484 12910 15486 12962
rect 15538 12910 15540 12962
rect 15484 12404 15540 12910
rect 15484 12338 15540 12348
rect 15260 12180 15316 12190
rect 15596 12180 15652 13132
rect 15708 12404 15764 13918
rect 15820 13858 15876 16268
rect 16044 16324 16100 17502
rect 16268 17554 16324 17566
rect 16268 17502 16270 17554
rect 16322 17502 16324 17554
rect 16268 17444 16324 17502
rect 16268 17378 16324 17388
rect 16380 16884 16436 16894
rect 16492 16884 16548 17836
rect 16604 17826 16660 17836
rect 16716 17892 16772 18286
rect 16716 17826 16772 17836
rect 16828 17668 16884 17678
rect 16828 17574 16884 17612
rect 16940 17444 16996 17454
rect 16380 16882 16548 16884
rect 16380 16830 16382 16882
rect 16434 16830 16548 16882
rect 16380 16828 16548 16830
rect 16380 16818 16436 16828
rect 16044 16258 16100 16268
rect 16492 16210 16548 16828
rect 16492 16158 16494 16210
rect 16546 16158 16548 16210
rect 16492 16146 16548 16158
rect 16716 17106 16772 17118
rect 16716 17054 16718 17106
rect 16770 17054 16772 17106
rect 16044 16100 16100 16110
rect 16044 15538 16100 16044
rect 16380 16098 16436 16110
rect 16380 16046 16382 16098
rect 16434 16046 16436 16098
rect 16380 15988 16436 16046
rect 16380 15764 16436 15932
rect 16380 15698 16436 15708
rect 16044 15486 16046 15538
rect 16098 15486 16100 15538
rect 16044 15474 16100 15486
rect 16156 15540 16212 15550
rect 15932 15426 15988 15438
rect 15932 15374 15934 15426
rect 15986 15374 15988 15426
rect 15932 15316 15988 15374
rect 16156 15316 16212 15484
rect 15932 15260 16212 15316
rect 16156 14756 16212 15260
rect 16156 14624 16212 14700
rect 15932 14420 15988 14430
rect 15932 14326 15988 14364
rect 16044 14308 16100 14318
rect 16044 14214 16100 14252
rect 16604 14308 16660 14318
rect 16604 14214 16660 14252
rect 16716 14084 16772 17054
rect 16940 16994 16996 17388
rect 16940 16942 16942 16994
rect 16994 16942 16996 16994
rect 16940 16930 16996 16942
rect 17164 16100 17220 16110
rect 17164 16006 17220 16044
rect 17052 15876 17108 15886
rect 17052 15782 17108 15820
rect 16828 15540 16884 15550
rect 16828 15446 16884 15484
rect 17052 14420 17108 14430
rect 17052 14326 17108 14364
rect 16604 14028 16772 14084
rect 16492 13972 16548 13982
rect 16492 13878 16548 13916
rect 15820 13806 15822 13858
rect 15874 13806 15876 13858
rect 15820 13794 15876 13806
rect 16044 13748 16100 13758
rect 16044 13746 16436 13748
rect 16044 13694 16046 13746
rect 16098 13694 16436 13746
rect 16044 13692 16436 13694
rect 16044 13682 16100 13692
rect 15932 13524 15988 13534
rect 15932 13186 15988 13468
rect 15932 13134 15934 13186
rect 15986 13134 15988 13186
rect 15932 13122 15988 13134
rect 16380 13186 16436 13692
rect 16380 13134 16382 13186
rect 16434 13134 16436 13186
rect 16380 13122 16436 13134
rect 16492 13300 16548 13310
rect 16492 13074 16548 13244
rect 16492 13022 16494 13074
rect 16546 13022 16548 13074
rect 16492 13010 16548 13022
rect 15708 12348 15876 12404
rect 15260 12178 15652 12180
rect 15260 12126 15262 12178
rect 15314 12126 15652 12178
rect 15260 12124 15652 12126
rect 15708 12180 15764 12190
rect 15260 12114 15316 12124
rect 15708 12086 15764 12124
rect 14252 12068 14308 12078
rect 14252 11506 14308 12012
rect 14252 11454 14254 11506
rect 14306 11454 14308 11506
rect 14252 11442 14308 11454
rect 14924 11394 14980 11406
rect 14924 11342 14926 11394
rect 14978 11342 14980 11394
rect 10668 10770 10724 10780
rect 14812 10836 14868 10846
rect 14812 10742 14868 10780
rect 14700 10388 14756 10398
rect 14588 10386 14756 10388
rect 14588 10334 14702 10386
rect 14754 10334 14756 10386
rect 14588 10332 14756 10334
rect 14588 9938 14644 10332
rect 14700 10322 14756 10332
rect 14924 10052 14980 11342
rect 15148 11396 15204 11406
rect 15148 11302 15204 11340
rect 15708 11396 15764 11406
rect 15708 11302 15764 11340
rect 15820 10836 15876 12348
rect 15932 11452 16548 11508
rect 15932 11282 15988 11452
rect 15932 11230 15934 11282
rect 15986 11230 15988 11282
rect 15932 11218 15988 11230
rect 16044 11282 16100 11294
rect 16044 11230 16046 11282
rect 16098 11230 16100 11282
rect 15820 10724 15876 10780
rect 15932 10724 15988 10734
rect 15820 10722 15988 10724
rect 15820 10670 15934 10722
rect 15986 10670 15988 10722
rect 15820 10668 15988 10670
rect 15932 10658 15988 10668
rect 15596 10610 15652 10622
rect 15596 10558 15598 10610
rect 15650 10558 15652 10610
rect 15036 10500 15092 10510
rect 15036 10406 15092 10444
rect 14924 9986 14980 9996
rect 14588 9886 14590 9938
rect 14642 9886 14644 9938
rect 14588 9874 14644 9886
rect 15596 9938 15652 10558
rect 15596 9886 15598 9938
rect 15650 9886 15652 9938
rect 14700 9828 14756 9838
rect 14700 9734 14756 9772
rect 15596 9828 15652 9886
rect 16044 10498 16100 11230
rect 16492 10836 16548 11452
rect 16604 11060 16660 14028
rect 16716 13860 16772 13870
rect 16716 13766 16772 13804
rect 16828 13746 16884 13758
rect 16828 13694 16830 13746
rect 16882 13694 16884 13746
rect 16828 13524 16884 13694
rect 16828 13458 16884 13468
rect 17276 11284 17332 22652
rect 17836 22260 17892 23886
rect 18284 23940 18340 24556
rect 18284 23874 18340 23884
rect 17948 23492 18004 23502
rect 17948 23378 18004 23436
rect 17948 23326 17950 23378
rect 18002 23326 18004 23378
rect 17948 23314 18004 23326
rect 19180 23156 19236 26348
rect 19628 26290 19684 26302
rect 19628 26238 19630 26290
rect 19682 26238 19684 26290
rect 19628 26180 19684 26238
rect 19852 26292 19908 26302
rect 19852 26198 19908 26236
rect 19628 26114 19684 26124
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19836 23548 20100 23558
rect 19404 23492 19460 23502
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20300 23492 20356 26908
rect 20412 26292 20468 29484
rect 20412 26198 20468 26236
rect 20524 26964 20580 26974
rect 20412 25284 20468 25294
rect 20412 25190 20468 25228
rect 20412 23716 20468 23726
rect 20524 23716 20580 26908
rect 20860 26180 20916 26190
rect 20860 26086 20916 26124
rect 20972 25732 21028 25742
rect 20972 25638 21028 25676
rect 21196 24724 21252 38612
rect 21532 37490 21588 43148
rect 22204 42756 22260 44380
rect 22092 42700 22260 42756
rect 22316 43540 22372 43550
rect 21644 42530 21700 42542
rect 21644 42478 21646 42530
rect 21698 42478 21700 42530
rect 21644 42196 21700 42478
rect 21644 42084 21700 42140
rect 21644 42028 21924 42084
rect 21868 41972 21924 42028
rect 22092 41972 22148 42700
rect 22316 42644 22372 43484
rect 22428 43204 22484 45164
rect 22652 44996 22708 48860
rect 22764 47458 22820 47470
rect 22764 47406 22766 47458
rect 22818 47406 22820 47458
rect 22764 47012 22820 47406
rect 22764 46946 22820 46956
rect 22764 45666 22820 45678
rect 22764 45614 22766 45666
rect 22818 45614 22820 45666
rect 22764 45444 22820 45614
rect 22764 45378 22820 45388
rect 22764 45220 22820 45230
rect 22764 45126 22820 45164
rect 22652 44940 22820 44996
rect 22540 44100 22596 44110
rect 22540 44098 22708 44100
rect 22540 44046 22542 44098
rect 22594 44046 22708 44098
rect 22540 44044 22708 44046
rect 22540 44034 22596 44044
rect 22540 43538 22596 43550
rect 22540 43486 22542 43538
rect 22594 43486 22596 43538
rect 22540 43428 22596 43486
rect 22540 43362 22596 43372
rect 22428 43138 22484 43148
rect 22652 42980 22708 44044
rect 22652 42914 22708 42924
rect 22652 42756 22708 42766
rect 22428 42644 22484 42654
rect 22316 42642 22484 42644
rect 22316 42590 22430 42642
rect 22482 42590 22484 42642
rect 22316 42588 22484 42590
rect 22204 42532 22260 42542
rect 22204 42438 22260 42476
rect 22428 42196 22484 42588
rect 22540 42642 22596 42654
rect 22540 42590 22542 42642
rect 22594 42590 22596 42642
rect 22540 42532 22596 42590
rect 22652 42642 22708 42700
rect 22652 42590 22654 42642
rect 22706 42590 22708 42642
rect 22652 42578 22708 42590
rect 22540 42466 22596 42476
rect 22428 42130 22484 42140
rect 22652 42084 22708 42094
rect 22540 41972 22596 41982
rect 21868 41916 22036 41972
rect 21756 41858 21812 41870
rect 21756 41806 21758 41858
rect 21810 41806 21812 41858
rect 21756 41746 21812 41806
rect 21756 41694 21758 41746
rect 21810 41694 21812 41746
rect 21756 41682 21812 41694
rect 21868 41524 21924 41534
rect 21868 41410 21924 41468
rect 21868 41358 21870 41410
rect 21922 41358 21924 41410
rect 21868 41346 21924 41358
rect 21644 41076 21700 41086
rect 21644 40982 21700 41020
rect 21980 40964 22036 41916
rect 21980 40898 22036 40908
rect 22092 41970 22596 41972
rect 22092 41918 22094 41970
rect 22146 41918 22542 41970
rect 22594 41918 22596 41970
rect 22092 41916 22596 41918
rect 21980 40628 22036 40638
rect 22092 40628 22148 41916
rect 22540 41906 22596 41916
rect 22204 41412 22260 41422
rect 22204 41318 22260 41356
rect 22540 41076 22596 41086
rect 21644 40626 22148 40628
rect 21644 40574 21982 40626
rect 22034 40574 22148 40626
rect 21644 40572 22148 40574
rect 22204 40964 22260 40974
rect 21644 39730 21700 40572
rect 21980 40562 22036 40572
rect 21868 40404 21924 40414
rect 22092 40404 22148 40442
rect 21924 40348 22036 40404
rect 21868 40338 21924 40348
rect 21644 39678 21646 39730
rect 21698 39678 21700 39730
rect 21644 39508 21700 39678
rect 21644 39442 21700 39452
rect 21756 39844 21812 39854
rect 21644 38836 21700 38846
rect 21644 38610 21700 38780
rect 21644 38558 21646 38610
rect 21698 38558 21700 38610
rect 21644 38546 21700 38558
rect 21644 37940 21700 37950
rect 21644 37846 21700 37884
rect 21532 37438 21534 37490
rect 21586 37438 21588 37490
rect 21532 37426 21588 37438
rect 21420 37380 21476 37390
rect 21420 37286 21476 37324
rect 21644 37380 21700 37390
rect 21644 37286 21700 37324
rect 21644 36370 21700 36382
rect 21644 36318 21646 36370
rect 21698 36318 21700 36370
rect 21644 36260 21700 36318
rect 21756 36370 21812 39788
rect 21868 39620 21924 39630
rect 21868 39526 21924 39564
rect 21980 38164 22036 40348
rect 22092 40338 22148 40348
rect 22204 40402 22260 40908
rect 22204 40350 22206 40402
rect 22258 40350 22260 40402
rect 22204 40338 22260 40350
rect 22428 40514 22484 40526
rect 22428 40462 22430 40514
rect 22482 40462 22484 40514
rect 22092 40180 22148 40190
rect 22092 39842 22148 40124
rect 22092 39790 22094 39842
rect 22146 39790 22148 39842
rect 22092 39778 22148 39790
rect 22428 39844 22484 40462
rect 22540 40180 22596 41020
rect 22652 40404 22708 42028
rect 22652 40338 22708 40348
rect 22540 40124 22708 40180
rect 22428 39778 22484 39788
rect 22204 39732 22260 39742
rect 22204 38388 22260 39676
rect 22540 39620 22596 39630
rect 22540 39526 22596 39564
rect 22316 39508 22372 39518
rect 22316 38668 22372 39452
rect 22652 38724 22708 40124
rect 22316 38612 22484 38668
rect 22652 38630 22708 38668
rect 22204 38332 22372 38388
rect 22092 38164 22148 38174
rect 21980 38162 22148 38164
rect 21980 38110 22094 38162
rect 22146 38110 22148 38162
rect 21980 38108 22148 38110
rect 22092 38098 22148 38108
rect 22204 38164 22260 38174
rect 22204 37490 22260 38108
rect 22204 37438 22206 37490
rect 22258 37438 22260 37490
rect 22204 37426 22260 37438
rect 21980 37268 22036 37278
rect 21756 36318 21758 36370
rect 21810 36318 21812 36370
rect 21756 36306 21812 36318
rect 21868 36708 21924 36718
rect 21644 36194 21700 36204
rect 21868 36148 21924 36652
rect 21980 36482 22036 37212
rect 21980 36430 21982 36482
rect 22034 36430 22036 36482
rect 21980 36418 22036 36430
rect 21868 36082 21924 36092
rect 21644 35924 21700 35934
rect 21644 35830 21700 35868
rect 21532 35812 21588 35822
rect 21532 35718 21588 35756
rect 21868 35698 21924 35710
rect 21868 35646 21870 35698
rect 21922 35646 21924 35698
rect 21868 35252 21924 35646
rect 21868 35186 21924 35196
rect 22092 35364 22148 35374
rect 21532 34690 21588 34702
rect 21532 34638 21534 34690
rect 21586 34638 21588 34690
rect 21532 34020 21588 34638
rect 21644 34468 21700 34478
rect 21644 34354 21700 34412
rect 21644 34302 21646 34354
rect 21698 34302 21700 34354
rect 21644 34290 21700 34302
rect 21868 34132 21924 34142
rect 21868 34038 21924 34076
rect 21532 33954 21588 33964
rect 22092 33458 22148 35308
rect 22092 33406 22094 33458
rect 22146 33406 22148 33458
rect 22092 33394 22148 33406
rect 21644 33236 21700 33246
rect 21644 33142 21700 33180
rect 22092 32788 22148 32798
rect 22092 32694 22148 32732
rect 21980 31892 22036 31902
rect 21980 31798 22036 31836
rect 22316 31220 22372 38332
rect 22428 36260 22484 38612
rect 22540 38388 22596 38398
rect 22540 37940 22596 38332
rect 22652 37940 22708 37950
rect 22540 37938 22708 37940
rect 22540 37886 22654 37938
rect 22706 37886 22708 37938
rect 22540 37884 22708 37886
rect 22540 37716 22596 37726
rect 22540 37490 22596 37660
rect 22540 37438 22542 37490
rect 22594 37438 22596 37490
rect 22540 37426 22596 37438
rect 22652 37044 22708 37884
rect 22652 36820 22708 36988
rect 22540 36764 22708 36820
rect 22540 36482 22596 36764
rect 22540 36430 22542 36482
rect 22594 36430 22596 36482
rect 22540 36418 22596 36430
rect 22652 36260 22708 36270
rect 22428 36204 22652 36260
rect 22428 35922 22484 36204
rect 22652 36128 22708 36204
rect 22428 35870 22430 35922
rect 22482 35870 22484 35922
rect 22428 35858 22484 35870
rect 22652 35698 22708 35710
rect 22652 35646 22654 35698
rect 22706 35646 22708 35698
rect 22652 35252 22708 35646
rect 22428 34132 22484 34142
rect 22652 34132 22708 35196
rect 22764 35140 22820 44940
rect 22876 41412 22932 49420
rect 23212 49476 23268 49486
rect 23212 49250 23268 49420
rect 23212 49198 23214 49250
rect 23266 49198 23268 49250
rect 23212 49186 23268 49198
rect 23324 49252 23380 49534
rect 23436 49252 23492 50876
rect 23772 50482 23828 50494
rect 23772 50430 23774 50482
rect 23826 50430 23828 50482
rect 23772 49924 23828 50430
rect 23772 49858 23828 49868
rect 23884 50484 23940 51324
rect 23996 51378 24052 51390
rect 23996 51326 23998 51378
rect 24050 51326 24052 51378
rect 23996 50932 24052 51326
rect 24108 51380 24164 51548
rect 24108 51314 24164 51324
rect 23996 50866 24052 50876
rect 23324 49196 23716 49252
rect 23324 49026 23380 49038
rect 23548 49028 23604 49038
rect 23324 48974 23326 49026
rect 23378 48974 23380 49026
rect 23100 48916 23156 48926
rect 22988 48468 23044 48478
rect 22988 48242 23044 48412
rect 22988 48190 22990 48242
rect 23042 48190 23044 48242
rect 22988 48178 23044 48190
rect 23100 47458 23156 48860
rect 23212 48804 23268 48814
rect 23212 48710 23268 48748
rect 23212 48244 23268 48254
rect 23324 48244 23380 48974
rect 23436 49026 23604 49028
rect 23436 48974 23550 49026
rect 23602 48974 23604 49026
rect 23436 48972 23604 48974
rect 23436 48916 23492 48972
rect 23548 48962 23604 48972
rect 23436 48850 23492 48860
rect 23548 48692 23604 48702
rect 23268 48188 23380 48244
rect 23436 48356 23492 48366
rect 23212 48150 23268 48188
rect 23324 47684 23380 47694
rect 23324 47570 23380 47628
rect 23324 47518 23326 47570
rect 23378 47518 23380 47570
rect 23324 47506 23380 47518
rect 23100 47406 23102 47458
rect 23154 47406 23156 47458
rect 23100 47394 23156 47406
rect 23436 47460 23492 48300
rect 23548 48242 23604 48636
rect 23660 48580 23716 49196
rect 23884 48692 23940 50428
rect 24108 50372 24164 50382
rect 24108 50370 24276 50372
rect 24108 50318 24110 50370
rect 24162 50318 24276 50370
rect 24108 50316 24276 50318
rect 24108 50306 24164 50316
rect 24220 49922 24276 50316
rect 24332 50148 24388 54796
rect 24444 54628 24500 54638
rect 24444 54534 24500 54572
rect 24556 54626 24612 54638
rect 24556 54574 24558 54626
rect 24610 54574 24612 54626
rect 24556 54516 24612 54574
rect 24556 54450 24612 54460
rect 24780 54516 24836 54526
rect 25004 54516 25060 55022
rect 24780 54514 24948 54516
rect 24780 54462 24782 54514
rect 24834 54462 24948 54514
rect 24780 54460 24948 54462
rect 24780 54450 24836 54460
rect 24556 53508 24612 53518
rect 24556 53414 24612 53452
rect 24444 52834 24500 52846
rect 24444 52782 24446 52834
rect 24498 52782 24500 52834
rect 24444 52500 24500 52782
rect 24780 52836 24836 52846
rect 24780 52742 24836 52780
rect 24444 52444 24836 52500
rect 24556 52164 24612 52174
rect 24556 51828 24612 52108
rect 24668 52052 24724 52062
rect 24780 52052 24836 52444
rect 24892 52388 24948 54460
rect 25004 54450 25060 54460
rect 25564 55074 25732 55076
rect 25564 55022 25678 55074
rect 25730 55022 25732 55074
rect 25564 55020 25732 55022
rect 25452 54068 25508 54078
rect 25452 53844 25508 54012
rect 25452 53712 25508 53788
rect 25004 53620 25060 53630
rect 25004 53526 25060 53564
rect 25340 53060 25396 53070
rect 25228 52388 25284 52398
rect 24892 52332 25060 52388
rect 25004 52164 25060 52332
rect 25228 52294 25284 52332
rect 25004 52098 25060 52108
rect 24892 52052 24948 52062
rect 24780 51996 24892 52052
rect 24668 51958 24724 51996
rect 24892 51958 24948 51996
rect 25116 51938 25172 51950
rect 25116 51886 25118 51938
rect 25170 51886 25172 51938
rect 25116 51828 25172 51886
rect 24556 51772 25172 51828
rect 25340 51828 25396 53004
rect 25564 52724 25620 55020
rect 25676 55010 25732 55020
rect 25788 54738 25844 55132
rect 25788 54686 25790 54738
rect 25842 54686 25844 54738
rect 25788 54674 25844 54686
rect 24556 51602 24612 51772
rect 25340 51762 25396 51772
rect 25452 52668 25620 52724
rect 25676 53732 25732 53742
rect 24556 51550 24558 51602
rect 24610 51550 24612 51602
rect 24556 51538 24612 51550
rect 24780 51492 24836 51502
rect 24780 51398 24836 51436
rect 24892 51378 24948 51390
rect 24892 51326 24894 51378
rect 24946 51326 24948 51378
rect 24892 51268 24948 51326
rect 24668 51212 24948 51268
rect 24444 50708 24500 50718
rect 24668 50708 24724 51212
rect 24444 50706 24724 50708
rect 24444 50654 24446 50706
rect 24498 50654 24724 50706
rect 24444 50652 24724 50654
rect 24444 50642 24500 50652
rect 24332 50092 24500 50148
rect 24220 49870 24222 49922
rect 24274 49870 24276 49922
rect 24220 49858 24276 49870
rect 24332 49924 24388 49934
rect 24108 49140 24164 49150
rect 24108 49046 24164 49084
rect 23884 48636 24052 48692
rect 23660 48524 23940 48580
rect 23660 48356 23716 48366
rect 23660 48262 23716 48300
rect 23548 48190 23550 48242
rect 23602 48190 23604 48242
rect 23548 48178 23604 48190
rect 23884 48242 23940 48524
rect 23884 48190 23886 48242
rect 23938 48190 23940 48242
rect 23772 48130 23828 48142
rect 23772 48078 23774 48130
rect 23826 48078 23828 48130
rect 22988 47348 23044 47358
rect 23436 47328 23492 47404
rect 23548 47908 23604 47918
rect 22988 46900 23044 47292
rect 23212 47234 23268 47246
rect 23212 47182 23214 47234
rect 23266 47182 23268 47234
rect 23100 46900 23156 46910
rect 22988 46898 23156 46900
rect 22988 46846 23102 46898
rect 23154 46846 23156 46898
rect 22988 46844 23156 46846
rect 23100 46834 23156 46844
rect 23212 46900 23268 47182
rect 23212 46834 23268 46844
rect 23436 46674 23492 46686
rect 23436 46622 23438 46674
rect 23490 46622 23492 46674
rect 23100 45892 23156 45902
rect 23100 45332 23156 45836
rect 23436 45892 23492 46622
rect 23436 45760 23492 45836
rect 22988 45330 23156 45332
rect 22988 45278 23102 45330
rect 23154 45278 23156 45330
rect 22988 45276 23156 45278
rect 22988 43708 23044 45276
rect 23100 45266 23156 45276
rect 23212 44324 23268 44334
rect 23212 44230 23268 44268
rect 23324 44324 23380 44334
rect 23436 44324 23492 44334
rect 23324 44322 23436 44324
rect 23324 44270 23326 44322
rect 23378 44270 23436 44322
rect 23324 44268 23436 44270
rect 23100 44210 23156 44222
rect 23100 44158 23102 44210
rect 23154 44158 23156 44210
rect 23100 44100 23156 44158
rect 23100 44034 23156 44044
rect 23324 43876 23380 44268
rect 23436 44258 23492 44268
rect 23324 43810 23380 43820
rect 22988 43652 23156 43708
rect 22988 43538 23044 43550
rect 22988 43486 22990 43538
rect 23042 43486 23044 43538
rect 22988 42866 23044 43486
rect 22988 42814 22990 42866
rect 23042 42814 23044 42866
rect 22988 42802 23044 42814
rect 23100 42756 23156 43652
rect 23100 42532 23156 42700
rect 23100 42466 23156 42476
rect 23436 43650 23492 43662
rect 23436 43598 23438 43650
rect 23490 43598 23492 43650
rect 23324 42196 23380 42206
rect 23324 42102 23380 42140
rect 23100 41970 23156 41982
rect 23100 41918 23102 41970
rect 23154 41918 23156 41970
rect 23100 41748 23156 41918
rect 23100 41682 23156 41692
rect 23212 41858 23268 41870
rect 23212 41806 23214 41858
rect 23266 41806 23268 41858
rect 23212 41636 23268 41806
rect 23212 41570 23268 41580
rect 23324 41860 23380 41870
rect 22876 41346 22932 41356
rect 22988 41186 23044 41198
rect 22988 41134 22990 41186
rect 23042 41134 23044 41186
rect 22988 39620 23044 41134
rect 23100 40964 23156 40974
rect 23100 40962 23268 40964
rect 23100 40910 23102 40962
rect 23154 40910 23268 40962
rect 23100 40908 23268 40910
rect 23100 40898 23156 40908
rect 23100 40402 23156 40414
rect 23100 40350 23102 40402
rect 23154 40350 23156 40402
rect 23100 39842 23156 40350
rect 23100 39790 23102 39842
rect 23154 39790 23156 39842
rect 23100 39778 23156 39790
rect 22988 39488 23044 39564
rect 23100 39396 23156 39406
rect 23212 39396 23268 40908
rect 23324 40516 23380 41804
rect 23436 40740 23492 43598
rect 23548 43652 23604 47852
rect 23660 47796 23716 47806
rect 23660 45444 23716 47740
rect 23772 47348 23828 48078
rect 23884 47460 23940 48190
rect 23996 47796 24052 48636
rect 24332 48244 24388 49868
rect 24108 48188 24388 48244
rect 24108 47908 24164 48188
rect 24444 48020 24500 50092
rect 24556 49812 24612 49822
rect 24556 49718 24612 49756
rect 24556 49364 24612 49374
rect 24556 49138 24612 49308
rect 24556 49086 24558 49138
rect 24610 49086 24612 49138
rect 24556 49074 24612 49086
rect 24668 49140 24724 50652
rect 24668 49074 24724 49084
rect 24780 51044 24836 51054
rect 24668 48804 24724 48814
rect 24556 48132 24612 48142
rect 24668 48132 24724 48748
rect 24780 48692 24836 50988
rect 25340 50708 25396 50718
rect 24892 50484 24948 50522
rect 24892 50418 24948 50428
rect 24892 49924 24948 49934
rect 24892 49830 24948 49868
rect 25116 49252 25172 49262
rect 25116 49140 25172 49196
rect 25340 49250 25396 50652
rect 25452 49364 25508 52668
rect 25564 52052 25620 52062
rect 25564 51958 25620 51996
rect 25676 51604 25732 53676
rect 26012 53620 26068 55580
rect 26236 55188 26292 55198
rect 26236 55094 26292 55132
rect 26348 54738 26404 55804
rect 26348 54686 26350 54738
rect 26402 54686 26404 54738
rect 26348 54674 26404 54686
rect 25788 53564 26068 53620
rect 25788 52276 25844 53564
rect 26124 53508 26180 53518
rect 26012 53506 26180 53508
rect 26012 53454 26126 53506
rect 26178 53454 26180 53506
rect 26012 53452 26180 53454
rect 26012 53060 26068 53452
rect 26124 53442 26180 53452
rect 25900 53058 26068 53060
rect 25900 53006 26014 53058
rect 26066 53006 26068 53058
rect 25900 53004 26068 53006
rect 25900 52500 25956 53004
rect 26012 52994 26068 53004
rect 26124 53060 26180 53070
rect 26124 52966 26180 53004
rect 26460 52836 26516 56252
rect 27468 56308 27524 56318
rect 27468 56214 27524 56252
rect 28924 56308 28980 59200
rect 33852 58212 33908 58222
rect 33628 56756 33684 56766
rect 32956 56644 33012 56654
rect 31276 56420 31332 56430
rect 28924 56242 28980 56252
rect 30268 56308 30324 56318
rect 26572 56196 26628 56206
rect 26572 55524 26628 56140
rect 30268 56194 30324 56252
rect 31276 56306 31332 56364
rect 31276 56254 31278 56306
rect 31330 56254 31332 56306
rect 31276 56242 31332 56254
rect 30268 56142 30270 56194
rect 30322 56142 30324 56194
rect 30268 56130 30324 56142
rect 26572 55458 26628 55468
rect 27916 56082 27972 56094
rect 27916 56030 27918 56082
rect 27970 56030 27972 56082
rect 26684 55074 26740 55086
rect 26684 55022 26686 55074
rect 26738 55022 26740 55074
rect 26572 54626 26628 54638
rect 26572 54574 26574 54626
rect 26626 54574 26628 54626
rect 26572 53844 26628 54574
rect 26684 54628 26740 55022
rect 27132 55074 27188 55086
rect 27132 55022 27134 55074
rect 27186 55022 27188 55074
rect 27132 54852 27188 55022
rect 27916 54964 27972 56030
rect 28252 56082 28308 56094
rect 28252 56030 28254 56082
rect 28306 56030 28308 56082
rect 27916 54898 27972 54908
rect 28028 55298 28084 55310
rect 28028 55246 28030 55298
rect 28082 55246 28084 55298
rect 27132 54786 27188 54796
rect 27244 54740 27300 54750
rect 26684 54562 26740 54572
rect 26908 54628 26964 54638
rect 26908 54534 26964 54572
rect 26796 54516 26852 54526
rect 26796 54422 26852 54460
rect 26684 54404 26740 54414
rect 26684 54310 26740 54348
rect 26572 53778 26628 53788
rect 27020 53844 27076 53854
rect 26460 52770 26516 52780
rect 26572 53620 26628 53630
rect 26012 52722 26068 52734
rect 26012 52670 26014 52722
rect 26066 52670 26068 52722
rect 26012 52500 26068 52670
rect 26460 52500 26516 52510
rect 26012 52444 26404 52500
rect 25900 52434 25956 52444
rect 25788 52220 25956 52276
rect 25676 51538 25732 51548
rect 25564 51492 25620 51502
rect 25564 49924 25620 51436
rect 25788 50594 25844 50606
rect 25788 50542 25790 50594
rect 25842 50542 25844 50594
rect 25788 50372 25844 50542
rect 25788 50306 25844 50316
rect 25900 50260 25956 52220
rect 26348 52162 26404 52444
rect 26348 52110 26350 52162
rect 26402 52110 26404 52162
rect 26348 52098 26404 52110
rect 26124 52052 26180 52090
rect 26124 51986 26180 51996
rect 26460 51940 26516 52444
rect 26572 52164 26628 53564
rect 27020 53618 27076 53788
rect 27020 53566 27022 53618
rect 27074 53566 27076 53618
rect 27020 53554 27076 53566
rect 26796 53172 26852 53182
rect 26796 53078 26852 53116
rect 26684 52948 26740 52958
rect 26684 52388 26740 52892
rect 26908 52948 26964 52958
rect 26908 52946 27076 52948
rect 26908 52894 26910 52946
rect 26962 52894 27076 52946
rect 26908 52892 27076 52894
rect 26908 52882 26964 52892
rect 26684 52322 26740 52332
rect 26796 52836 26852 52846
rect 26572 52098 26628 52108
rect 26348 51884 26516 51940
rect 25900 50036 25956 50204
rect 26124 51828 26180 51838
rect 26124 50148 26180 51772
rect 26236 51604 26292 51614
rect 26236 51490 26292 51548
rect 26236 51438 26238 51490
rect 26290 51438 26292 51490
rect 26236 51426 26292 51438
rect 26012 50036 26068 50046
rect 25900 50034 26068 50036
rect 25900 49982 26014 50034
rect 26066 49982 26068 50034
rect 25900 49980 26068 49982
rect 26012 49970 26068 49980
rect 25564 49868 25844 49924
rect 25564 49698 25620 49710
rect 25564 49646 25566 49698
rect 25618 49646 25620 49698
rect 25564 49588 25620 49646
rect 25564 49522 25620 49532
rect 25452 49308 25732 49364
rect 25340 49198 25342 49250
rect 25394 49198 25396 49250
rect 25340 49186 25396 49198
rect 25116 49138 25284 49140
rect 25116 49086 25118 49138
rect 25170 49086 25284 49138
rect 25116 49084 25284 49086
rect 25116 49074 25172 49084
rect 24780 48626 24836 48636
rect 25228 48468 25284 49084
rect 25340 49028 25396 49038
rect 25340 48916 25396 48972
rect 25340 48860 25508 48916
rect 25452 48802 25508 48860
rect 25452 48750 25454 48802
rect 25506 48750 25508 48802
rect 25452 48738 25508 48750
rect 25564 48468 25620 48478
rect 25228 48466 25620 48468
rect 25228 48414 25566 48466
rect 25618 48414 25620 48466
rect 25228 48412 25620 48414
rect 25564 48402 25620 48412
rect 24556 48130 24724 48132
rect 24556 48078 24558 48130
rect 24610 48078 24724 48130
rect 24556 48076 24724 48078
rect 24780 48354 24836 48366
rect 24780 48302 24782 48354
rect 24834 48302 24836 48354
rect 24556 48066 24612 48076
rect 24108 47842 24164 47852
rect 24220 47964 24500 48020
rect 23996 47730 24052 47740
rect 24108 47460 24164 47470
rect 23884 47458 24164 47460
rect 23884 47406 24110 47458
rect 24162 47406 24164 47458
rect 23884 47404 24164 47406
rect 24108 47394 24164 47404
rect 23772 47282 23828 47292
rect 23884 46564 23940 46574
rect 23884 46562 24052 46564
rect 23884 46510 23886 46562
rect 23938 46510 24052 46562
rect 23884 46508 24052 46510
rect 23884 46498 23940 46508
rect 23660 45330 23716 45388
rect 23660 45278 23662 45330
rect 23714 45278 23716 45330
rect 23660 45266 23716 45278
rect 23884 45892 23940 45902
rect 23660 44210 23716 44222
rect 23660 44158 23662 44210
rect 23714 44158 23716 44210
rect 23660 43652 23716 44158
rect 23884 43764 23940 45836
rect 23996 45778 24052 46508
rect 23996 45726 23998 45778
rect 24050 45726 24052 45778
rect 23996 43988 24052 45726
rect 24108 45444 24164 45454
rect 24108 44996 24164 45388
rect 24220 45220 24276 47964
rect 24780 47908 24836 48302
rect 24892 48132 24948 48142
rect 24892 48038 24948 48076
rect 24444 47852 24836 47908
rect 25228 48020 25284 48030
rect 24444 47682 24500 47852
rect 24444 47630 24446 47682
rect 24498 47630 24500 47682
rect 24444 47618 24500 47630
rect 24444 47460 24500 47470
rect 24444 47366 24500 47404
rect 24892 47460 24948 47470
rect 24332 46676 24388 46686
rect 24332 46582 24388 46620
rect 24780 46562 24836 46574
rect 24780 46510 24782 46562
rect 24834 46510 24836 46562
rect 24780 46452 24836 46510
rect 24780 46386 24836 46396
rect 24220 45164 24388 45220
rect 24220 44996 24276 45006
rect 24108 44994 24276 44996
rect 24108 44942 24222 44994
rect 24274 44942 24276 44994
rect 24108 44940 24276 44942
rect 24220 44930 24276 44940
rect 24108 44324 24164 44334
rect 24108 44230 24164 44268
rect 23996 43922 24052 43932
rect 24220 44212 24276 44222
rect 23884 43708 24164 43764
rect 23660 43596 24052 43652
rect 23548 43540 23604 43596
rect 23548 43484 23828 43540
rect 23660 42756 23716 42766
rect 23548 42644 23604 42654
rect 23548 40852 23604 42588
rect 23660 42642 23716 42700
rect 23660 42590 23662 42642
rect 23714 42590 23716 42642
rect 23660 41860 23716 42590
rect 23772 42084 23828 43484
rect 23772 41970 23828 42028
rect 23772 41918 23774 41970
rect 23826 41918 23828 41970
rect 23772 41906 23828 41918
rect 23996 43538 24052 43596
rect 23996 43486 23998 43538
rect 24050 43486 24052 43538
rect 23996 42642 24052 43486
rect 23996 42590 23998 42642
rect 24050 42590 24052 42642
rect 23660 41794 23716 41804
rect 23772 41188 23828 41198
rect 23772 41094 23828 41132
rect 23548 40786 23604 40796
rect 23436 40674 23492 40684
rect 23436 40516 23492 40526
rect 23324 40514 23492 40516
rect 23324 40462 23438 40514
rect 23490 40462 23492 40514
rect 23324 40460 23492 40462
rect 23436 40450 23492 40460
rect 23548 40404 23604 40414
rect 23548 40310 23604 40348
rect 23660 40402 23716 40414
rect 23660 40350 23662 40402
rect 23714 40350 23716 40402
rect 23660 40292 23716 40350
rect 23660 40226 23716 40236
rect 23884 40178 23940 40190
rect 23884 40126 23886 40178
rect 23938 40126 23940 40178
rect 23156 39340 23268 39396
rect 23660 39844 23716 39854
rect 23660 39396 23716 39788
rect 23772 39396 23828 39406
rect 23660 39394 23828 39396
rect 23660 39342 23774 39394
rect 23826 39342 23828 39394
rect 23660 39340 23828 39342
rect 23100 39302 23156 39340
rect 23212 38948 23268 38958
rect 23212 38854 23268 38892
rect 23212 38724 23268 38734
rect 23212 38162 23268 38668
rect 23660 38668 23716 39340
rect 23772 39330 23828 39340
rect 23772 38836 23828 38846
rect 23884 38836 23940 40126
rect 23772 38834 23940 38836
rect 23772 38782 23774 38834
rect 23826 38782 23940 38834
rect 23772 38780 23940 38782
rect 23772 38770 23828 38780
rect 23660 38612 23940 38668
rect 23660 38388 23716 38398
rect 23660 38274 23716 38332
rect 23660 38222 23662 38274
rect 23714 38222 23716 38274
rect 23212 38110 23214 38162
rect 23266 38110 23268 38162
rect 23212 38098 23268 38110
rect 23436 38164 23492 38174
rect 23492 38108 23604 38164
rect 23436 38070 23492 38108
rect 23324 37828 23380 37838
rect 22876 37436 23268 37492
rect 22876 36482 22932 37436
rect 23212 37378 23268 37436
rect 23212 37326 23214 37378
rect 23266 37326 23268 37378
rect 23212 37314 23268 37326
rect 23324 37380 23380 37772
rect 23548 37492 23604 38108
rect 23660 38052 23716 38222
rect 23660 37986 23716 37996
rect 23772 37492 23828 37502
rect 23548 37436 23716 37492
rect 22876 36430 22878 36482
rect 22930 36430 22932 36482
rect 22876 36418 22932 36430
rect 23212 37044 23268 37054
rect 23212 35922 23268 36988
rect 23324 36370 23380 37324
rect 23324 36318 23326 36370
rect 23378 36318 23380 36370
rect 23324 36306 23380 36318
rect 23548 37266 23604 37278
rect 23548 37214 23550 37266
rect 23602 37214 23604 37266
rect 23212 35870 23214 35922
rect 23266 35870 23268 35922
rect 22764 35084 22932 35140
rect 22764 34916 22820 34926
rect 22764 34354 22820 34860
rect 22764 34302 22766 34354
rect 22818 34302 22820 34354
rect 22764 34290 22820 34302
rect 22764 34132 22820 34142
rect 22652 34130 22820 34132
rect 22652 34078 22766 34130
rect 22818 34078 22820 34130
rect 22652 34076 22820 34078
rect 22428 34038 22484 34076
rect 22764 34066 22820 34076
rect 22540 34020 22596 34030
rect 22428 31890 22484 31902
rect 22428 31838 22430 31890
rect 22482 31838 22484 31890
rect 22428 31780 22484 31838
rect 22428 31714 22484 31724
rect 22540 31892 22596 33964
rect 22540 31666 22596 31836
rect 22540 31614 22542 31666
rect 22594 31614 22596 31666
rect 22540 31602 22596 31614
rect 22652 33234 22708 33246
rect 22652 33182 22654 33234
rect 22706 33182 22708 33234
rect 22652 32564 22708 33182
rect 22764 33236 22820 33246
rect 22876 33236 22932 35084
rect 23212 34468 23268 35870
rect 23548 35476 23604 37214
rect 23660 36932 23716 37436
rect 23772 37154 23828 37436
rect 23772 37102 23774 37154
rect 23826 37102 23828 37154
rect 23772 37090 23828 37102
rect 23884 37044 23940 38612
rect 23996 37716 24052 42590
rect 24108 42420 24164 43708
rect 24220 43650 24276 44156
rect 24220 43598 24222 43650
rect 24274 43598 24276 43650
rect 24220 43586 24276 43598
rect 24108 42364 24276 42420
rect 24108 41524 24164 41534
rect 24108 41298 24164 41468
rect 24108 41246 24110 41298
rect 24162 41246 24164 41298
rect 24108 41234 24164 41246
rect 24220 41074 24276 42364
rect 24220 41022 24222 41074
rect 24274 41022 24276 41074
rect 24108 40852 24164 40862
rect 24108 40626 24164 40796
rect 24108 40574 24110 40626
rect 24162 40574 24164 40626
rect 24108 39508 24164 40574
rect 24220 40178 24276 41022
rect 24220 40126 24222 40178
rect 24274 40126 24276 40178
rect 24220 39730 24276 40126
rect 24220 39678 24222 39730
rect 24274 39678 24276 39730
rect 24220 39666 24276 39678
rect 24332 39620 24388 45164
rect 24444 45108 24500 45118
rect 24444 45014 24500 45052
rect 24780 44884 24836 44894
rect 24780 44790 24836 44828
rect 24556 44772 24612 44782
rect 24556 44100 24612 44716
rect 24556 44006 24612 44044
rect 24444 42532 24500 42542
rect 24444 42438 24500 42476
rect 24668 41972 24724 41982
rect 24668 41878 24724 41916
rect 24556 41858 24612 41870
rect 24556 41806 24558 41858
rect 24610 41806 24612 41858
rect 24556 41636 24612 41806
rect 24556 41570 24612 41580
rect 24892 41300 24948 47404
rect 25116 47234 25172 47246
rect 25116 47182 25118 47234
rect 25170 47182 25172 47234
rect 25004 47124 25060 47134
rect 25004 43652 25060 47068
rect 25116 47012 25172 47182
rect 25116 46004 25172 46956
rect 25116 45938 25172 45948
rect 25228 44212 25284 47964
rect 25452 47572 25508 47582
rect 25452 47478 25508 47516
rect 25452 46900 25508 46910
rect 25452 45890 25508 46844
rect 25676 46788 25732 49308
rect 25452 45838 25454 45890
rect 25506 45838 25508 45890
rect 25452 45826 25508 45838
rect 25564 46732 25732 46788
rect 25452 45668 25508 45678
rect 25340 44660 25396 44670
rect 25340 44434 25396 44604
rect 25340 44382 25342 44434
rect 25394 44382 25396 44434
rect 25340 44370 25396 44382
rect 25228 44156 25396 44212
rect 25004 43596 25172 43652
rect 25004 43428 25060 43438
rect 25004 42084 25060 43372
rect 25004 41636 25060 42028
rect 25004 41570 25060 41580
rect 24556 41244 24948 41300
rect 24556 40626 24612 41244
rect 24556 40574 24558 40626
rect 24610 40574 24612 40626
rect 24556 39956 24612 40574
rect 24556 39890 24612 39900
rect 25004 39732 25060 39742
rect 25116 39732 25172 43596
rect 25228 42530 25284 42542
rect 25228 42478 25230 42530
rect 25282 42478 25284 42530
rect 25228 42084 25284 42478
rect 25228 42018 25284 42028
rect 25228 41300 25284 41310
rect 25228 41206 25284 41244
rect 24556 39730 25172 39732
rect 24556 39678 25006 39730
rect 25058 39678 25172 39730
rect 24556 39676 25172 39678
rect 25228 41076 25284 41086
rect 24332 39564 24500 39620
rect 24108 39452 24388 39508
rect 24220 38836 24276 38846
rect 24332 38836 24388 39452
rect 24220 38834 24388 38836
rect 24220 38782 24222 38834
rect 24274 38782 24388 38834
rect 24220 38780 24388 38782
rect 24220 38770 24276 38780
rect 24220 38274 24276 38286
rect 24444 38276 24500 39564
rect 24220 38222 24222 38274
rect 24274 38222 24276 38274
rect 24108 38164 24164 38174
rect 24220 38164 24276 38222
rect 24108 38162 24276 38164
rect 24108 38110 24110 38162
rect 24162 38110 24276 38162
rect 24108 38108 24276 38110
rect 24332 38220 24500 38276
rect 24556 38834 24612 39676
rect 25004 39666 25060 39676
rect 24556 38782 24558 38834
rect 24610 38782 24612 38834
rect 24556 38274 24612 38782
rect 24780 39508 24836 39518
rect 24668 38724 24724 38762
rect 24668 38658 24724 38668
rect 24556 38222 24558 38274
rect 24610 38222 24612 38274
rect 24108 38098 24164 38108
rect 23996 37650 24052 37660
rect 24220 37604 24276 37614
rect 24220 37266 24276 37548
rect 24220 37214 24222 37266
rect 24274 37214 24276 37266
rect 24220 37202 24276 37214
rect 23884 36988 24276 37044
rect 23660 36876 23828 36932
rect 23660 36372 23716 36382
rect 23660 36278 23716 36316
rect 23772 35922 23828 36876
rect 24220 36370 24276 36988
rect 24220 36318 24222 36370
rect 24274 36318 24276 36370
rect 24220 36306 24276 36318
rect 23772 35870 23774 35922
rect 23826 35870 23828 35922
rect 23772 35858 23828 35870
rect 23548 35410 23604 35420
rect 23996 35698 24052 35710
rect 23996 35646 23998 35698
rect 24050 35646 24052 35698
rect 23212 34402 23268 34412
rect 23436 35364 23492 35374
rect 23100 34244 23156 34254
rect 23100 34150 23156 34188
rect 23436 33346 23492 35308
rect 23996 35252 24052 35646
rect 23884 34804 23940 34814
rect 23884 34710 23940 34748
rect 23884 34242 23940 34254
rect 23884 34190 23886 34242
rect 23938 34190 23940 34242
rect 23884 34132 23940 34190
rect 23996 34244 24052 35196
rect 23996 34178 24052 34188
rect 24220 34354 24276 34366
rect 24220 34302 24222 34354
rect 24274 34302 24276 34354
rect 23884 33908 23940 34076
rect 24220 34020 24276 34302
rect 24220 33954 24276 33964
rect 23884 33852 24052 33908
rect 23884 33570 23940 33582
rect 23884 33518 23886 33570
rect 23938 33518 23940 33570
rect 23436 33294 23438 33346
rect 23490 33294 23492 33346
rect 23436 33282 23492 33294
rect 23772 33348 23828 33358
rect 23884 33348 23940 33518
rect 23772 33346 23940 33348
rect 23772 33294 23774 33346
rect 23826 33294 23940 33346
rect 23772 33292 23940 33294
rect 23772 33282 23828 33292
rect 22820 33180 22932 33236
rect 22764 33104 22820 33180
rect 22988 33124 23044 33134
rect 23548 33124 23604 33134
rect 22988 33122 23156 33124
rect 22988 33070 22990 33122
rect 23042 33070 23156 33122
rect 22988 33068 23156 33070
rect 22988 33058 23044 33068
rect 22988 32900 23044 32910
rect 22652 31444 22708 32508
rect 22876 32788 22932 32798
rect 22876 32562 22932 32732
rect 22876 32510 22878 32562
rect 22930 32510 22932 32562
rect 22876 32498 22932 32510
rect 22764 31668 22820 31678
rect 22764 31666 22932 31668
rect 22764 31614 22766 31666
rect 22818 31614 22932 31666
rect 22764 31612 22932 31614
rect 22764 31602 22820 31612
rect 22876 31556 22932 31612
rect 22652 31388 22820 31444
rect 22316 31154 22372 31164
rect 22540 31332 22596 31342
rect 21980 30772 22036 30782
rect 21868 30716 21980 30772
rect 21532 29988 21588 29998
rect 21420 29986 21588 29988
rect 21420 29934 21534 29986
rect 21586 29934 21588 29986
rect 21420 29932 21588 29934
rect 21420 29540 21476 29932
rect 21532 29922 21588 29932
rect 21420 29474 21476 29484
rect 21532 29764 21588 29774
rect 21532 29650 21588 29708
rect 21532 29598 21534 29650
rect 21586 29598 21588 29650
rect 21196 24658 21252 24668
rect 21308 27858 21364 27870
rect 21308 27806 21310 27858
rect 21362 27806 21364 27858
rect 21308 26290 21364 27806
rect 21308 26238 21310 26290
rect 21362 26238 21364 26290
rect 20412 23714 20580 23716
rect 20412 23662 20414 23714
rect 20466 23662 20580 23714
rect 20412 23660 20580 23662
rect 20636 24612 20692 24622
rect 20412 23650 20468 23660
rect 19180 23154 19348 23156
rect 19180 23102 19182 23154
rect 19234 23102 19348 23154
rect 19180 23100 19348 23102
rect 19180 23090 19236 23100
rect 18508 23044 18564 23054
rect 18508 23042 18900 23044
rect 18508 22990 18510 23042
rect 18562 22990 18900 23042
rect 18508 22988 18900 22990
rect 18508 22978 18564 22988
rect 18844 22372 18900 22988
rect 19292 22596 19348 23100
rect 19404 23154 19460 23436
rect 20300 23378 20356 23436
rect 20300 23326 20302 23378
rect 20354 23326 20356 23378
rect 20300 23314 20356 23326
rect 19404 23102 19406 23154
rect 19458 23102 19460 23154
rect 19404 23090 19460 23102
rect 20636 23156 20692 24556
rect 20972 24388 21028 24398
rect 20972 23714 21028 24332
rect 21308 24052 21364 26238
rect 21532 26852 21588 29598
rect 21868 28420 21924 30716
rect 21980 30640 22036 30716
rect 21980 30324 22036 30334
rect 21980 30230 22036 30268
rect 22428 29988 22484 30026
rect 22428 29922 22484 29932
rect 22316 29876 22372 29886
rect 22316 29650 22372 29820
rect 22316 29598 22318 29650
rect 22370 29598 22372 29650
rect 22316 29204 22372 29598
rect 22316 29138 22372 29148
rect 22428 29764 22484 29774
rect 22428 28756 22484 29708
rect 22428 28624 22484 28700
rect 21868 28354 21924 28364
rect 21644 27858 21700 27870
rect 21644 27806 21646 27858
rect 21698 27806 21700 27858
rect 21644 27636 21700 27806
rect 21644 27570 21700 27580
rect 21980 26964 22036 27002
rect 21980 26898 22036 26908
rect 21644 26852 21700 26862
rect 21532 26850 21700 26852
rect 21532 26798 21646 26850
rect 21698 26798 21700 26850
rect 21532 26796 21700 26798
rect 21532 25284 21588 26796
rect 21644 26786 21700 26796
rect 21868 26290 21924 26302
rect 21868 26238 21870 26290
rect 21922 26238 21924 26290
rect 21532 25190 21588 25228
rect 21756 26180 21812 26190
rect 21420 24948 21476 24958
rect 21420 24854 21476 24892
rect 21756 24948 21812 26124
rect 21868 25732 21924 26238
rect 21868 25666 21924 25676
rect 21868 24948 21924 24958
rect 21756 24946 21924 24948
rect 21756 24894 21870 24946
rect 21922 24894 21924 24946
rect 21756 24892 21924 24894
rect 21308 23986 21364 23996
rect 20972 23662 20974 23714
rect 21026 23662 21028 23714
rect 20748 23156 20804 23166
rect 20636 23154 20804 23156
rect 20636 23102 20750 23154
rect 20802 23102 20804 23154
rect 20636 23100 20804 23102
rect 20748 23090 20804 23100
rect 19292 22540 19796 22596
rect 19740 22482 19796 22540
rect 19740 22430 19742 22482
rect 19794 22430 19796 22482
rect 19740 22418 19796 22430
rect 18956 22372 19012 22382
rect 18844 22370 19012 22372
rect 18844 22318 18958 22370
rect 19010 22318 19012 22370
rect 18844 22316 19012 22318
rect 18956 22306 19012 22316
rect 17836 22194 17892 22204
rect 18732 22260 18788 22270
rect 18732 22166 18788 22204
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20860 19124 20916 19134
rect 18956 19012 19012 19022
rect 18172 18452 18228 18462
rect 18172 18358 18228 18396
rect 18956 18450 19012 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 18956 18398 18958 18450
rect 19010 18398 19012 18450
rect 18956 18386 19012 18398
rect 19628 18450 19684 18462
rect 19628 18398 19630 18450
rect 19682 18398 19684 18450
rect 17500 17892 17556 17902
rect 17500 17798 17556 17836
rect 17836 17668 17892 17678
rect 17836 17554 17892 17612
rect 17836 17502 17838 17554
rect 17890 17502 17892 17554
rect 17612 17444 17668 17454
rect 17612 17350 17668 17388
rect 17836 17108 17892 17502
rect 17836 17042 17892 17052
rect 18396 17554 18452 17566
rect 18396 17502 18398 17554
rect 18450 17502 18452 17554
rect 18396 16884 18452 17502
rect 18620 17556 18676 17566
rect 18620 17462 18676 17500
rect 18508 17444 18564 17454
rect 18508 17350 18564 17388
rect 17612 15540 17668 15550
rect 17612 14642 17668 15484
rect 18396 15538 18452 16828
rect 19628 16884 19684 18398
rect 20188 18450 20244 18462
rect 20188 18398 20190 18450
rect 20242 18398 20244 18450
rect 19852 17780 19908 17790
rect 19852 17686 19908 17724
rect 20188 17556 20244 18398
rect 20860 17890 20916 19068
rect 20860 17838 20862 17890
rect 20914 17838 20916 17890
rect 20860 17826 20916 17838
rect 20524 17780 20580 17790
rect 20524 17686 20580 17724
rect 20300 17668 20356 17678
rect 20300 17574 20356 17612
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 16818 19684 16828
rect 19964 16884 20020 16894
rect 19964 16790 20020 16828
rect 20188 16884 20244 17500
rect 20188 16818 20244 16828
rect 19180 16212 19236 16222
rect 18956 15986 19012 15998
rect 18956 15934 18958 15986
rect 19010 15934 19012 15986
rect 18956 15876 19012 15934
rect 18956 15810 19012 15820
rect 18396 15486 18398 15538
rect 18450 15486 18452 15538
rect 18396 15474 18452 15486
rect 18844 15764 18900 15774
rect 17612 14590 17614 14642
rect 17666 14590 17668 14642
rect 17612 14578 17668 14590
rect 18844 14642 18900 15708
rect 19180 15314 19236 16156
rect 19964 16212 20020 16222
rect 19964 16118 20020 16156
rect 19180 15262 19182 15314
rect 19234 15262 19236 15314
rect 18844 14590 18846 14642
rect 18898 14590 18900 14642
rect 18844 14578 18900 14590
rect 18956 14756 19012 14766
rect 18956 14530 19012 14700
rect 18956 14478 18958 14530
rect 19010 14478 19012 14530
rect 18956 14466 19012 14478
rect 17948 14308 18004 14318
rect 17948 13748 18004 14252
rect 18732 14306 18788 14318
rect 18732 14254 18734 14306
rect 18786 14254 18788 14306
rect 18732 13970 18788 14254
rect 18732 13918 18734 13970
rect 18786 13918 18788 13970
rect 18732 13906 18788 13918
rect 19180 13972 19236 15262
rect 19516 15874 19572 15886
rect 19516 15822 19518 15874
rect 19570 15822 19572 15874
rect 19404 14532 19460 14542
rect 19516 14532 19572 15822
rect 20412 15874 20468 15886
rect 20412 15822 20414 15874
rect 20466 15822 20468 15874
rect 20412 15764 20468 15822
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 20412 15202 20468 15708
rect 20412 15150 20414 15202
rect 20466 15150 20468 15202
rect 20412 15148 20468 15150
rect 19404 14530 19572 14532
rect 19404 14478 19406 14530
rect 19458 14478 19572 14530
rect 19404 14476 19572 14478
rect 20188 15092 20468 15148
rect 20524 15426 20580 15438
rect 20524 15374 20526 15426
rect 20578 15374 20580 15426
rect 20524 15092 20580 15374
rect 19404 14466 19460 14476
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19740 13972 19796 13982
rect 19180 13970 19796 13972
rect 19180 13918 19742 13970
rect 19794 13918 19796 13970
rect 19180 13916 19796 13918
rect 17948 13682 18004 13692
rect 19068 13748 19124 13758
rect 19180 13748 19236 13916
rect 19740 13906 19796 13916
rect 20188 13970 20244 15092
rect 20524 14756 20580 15036
rect 20524 14690 20580 14700
rect 20300 14644 20356 14654
rect 20300 14550 20356 14588
rect 20636 14532 20692 14542
rect 20636 14438 20692 14476
rect 20188 13918 20190 13970
rect 20242 13918 20244 13970
rect 19068 13746 19236 13748
rect 19068 13694 19070 13746
rect 19122 13694 19236 13746
rect 19068 13692 19236 13694
rect 19068 13682 19124 13692
rect 19292 13634 19348 13646
rect 19292 13582 19294 13634
rect 19346 13582 19348 13634
rect 19292 13524 19348 13582
rect 19516 13524 19572 13534
rect 19292 13522 19572 13524
rect 19292 13470 19518 13522
rect 19570 13470 19572 13522
rect 19292 13468 19572 13470
rect 19516 13458 19572 13468
rect 20188 13522 20244 13918
rect 20860 14418 20916 14430
rect 20860 14366 20862 14418
rect 20914 14366 20916 14418
rect 20860 13636 20916 14366
rect 20860 13542 20916 13580
rect 20188 13470 20190 13522
rect 20242 13470 20244 13522
rect 20188 13458 20244 13470
rect 19852 13076 19908 13086
rect 18956 12850 19012 12862
rect 18956 12798 18958 12850
rect 19010 12798 19012 12850
rect 18508 12740 18564 12750
rect 18508 12646 18564 12684
rect 18620 12180 18676 12190
rect 18284 12178 18676 12180
rect 18284 12126 18622 12178
rect 18674 12126 18676 12178
rect 18284 12124 18676 12126
rect 18284 11506 18340 12124
rect 18620 12114 18676 12124
rect 18956 12068 19012 12798
rect 19852 12850 19908 13020
rect 20860 13076 20916 13086
rect 19852 12798 19854 12850
rect 19906 12798 19908 12850
rect 19852 12786 19908 12798
rect 19964 12852 20020 12862
rect 19964 12758 20020 12796
rect 20524 12852 20580 12862
rect 18956 12002 19012 12012
rect 19068 12740 19124 12750
rect 19068 11956 19124 12684
rect 19068 11890 19124 11900
rect 19292 12738 19348 12750
rect 19292 12686 19294 12738
rect 19346 12686 19348 12738
rect 18284 11454 18286 11506
rect 18338 11454 18340 11506
rect 18284 11442 18340 11454
rect 17276 11218 17332 11228
rect 19292 11396 19348 12686
rect 19628 12738 19684 12750
rect 19628 12686 19630 12738
rect 19682 12686 19684 12738
rect 19516 12178 19572 12190
rect 19516 12126 19518 12178
rect 19570 12126 19572 12178
rect 19404 12068 19460 12078
rect 19404 11974 19460 12012
rect 19516 11956 19572 12126
rect 19516 11890 19572 11900
rect 19628 11620 19684 12686
rect 20524 12738 20580 12796
rect 20524 12686 20526 12738
rect 20578 12686 20580 12738
rect 20524 12628 20580 12686
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20524 12562 20580 12572
rect 19836 12506 20100 12516
rect 20860 12178 20916 13020
rect 20860 12126 20862 12178
rect 20914 12126 20916 12178
rect 20860 12114 20916 12126
rect 20300 12068 20356 12078
rect 20300 11974 20356 12012
rect 20524 11956 20580 11966
rect 18172 11172 18228 11182
rect 19180 11172 19236 11182
rect 18060 11170 18228 11172
rect 18060 11118 18174 11170
rect 18226 11118 18228 11170
rect 18060 11116 18228 11118
rect 16604 11004 16772 11060
rect 16604 10836 16660 10846
rect 16492 10834 16660 10836
rect 16492 10782 16606 10834
rect 16658 10782 16660 10834
rect 16492 10780 16660 10782
rect 16604 10770 16660 10780
rect 16268 10724 16324 10734
rect 16044 10446 16046 10498
rect 16098 10446 16100 10498
rect 16044 9940 16100 10446
rect 16156 10610 16212 10622
rect 16156 10558 16158 10610
rect 16210 10558 16212 10610
rect 16156 10500 16212 10558
rect 16156 10434 16212 10444
rect 16044 9874 16100 9884
rect 15596 9762 15652 9772
rect 16268 9826 16324 10668
rect 16492 10612 16548 10622
rect 16492 9938 16548 10556
rect 16716 10500 16772 11004
rect 17948 10834 18004 10846
rect 17948 10782 17950 10834
rect 18002 10782 18004 10834
rect 16828 10724 16884 10734
rect 16828 10630 16884 10668
rect 16940 10612 16996 10622
rect 16940 10518 16996 10556
rect 17724 10612 17780 10622
rect 17724 10518 17780 10556
rect 16716 10434 16772 10444
rect 17612 10500 17668 10510
rect 17500 10052 17556 10062
rect 17500 9958 17556 9996
rect 16492 9886 16494 9938
rect 16546 9886 16548 9938
rect 16492 9874 16548 9886
rect 16268 9774 16270 9826
rect 16322 9774 16324 9826
rect 16268 9762 16324 9774
rect 13804 9714 13860 9726
rect 13804 9662 13806 9714
rect 13858 9662 13860 9714
rect 9212 4498 9268 4508
rect 12684 9154 12740 9166
rect 12684 9102 12686 9154
rect 12738 9102 12740 9154
rect 6972 3614 6974 3666
rect 7026 3614 7028 3666
rect 6972 3602 7028 3614
rect 12236 3556 12292 3566
rect 12684 3556 12740 9102
rect 13020 9156 13076 9166
rect 13020 9062 13076 9100
rect 13804 9156 13860 9662
rect 13804 9090 13860 9100
rect 16492 9716 16548 9726
rect 16492 8482 16548 9660
rect 17612 9714 17668 10444
rect 17836 10052 17892 10062
rect 17836 9958 17892 9996
rect 17612 9662 17614 9714
rect 17666 9662 17668 9714
rect 17612 9650 17668 9662
rect 16492 8430 16494 8482
rect 16546 8430 16548 8482
rect 16492 8418 16548 8430
rect 17164 8370 17220 8382
rect 17164 8318 17166 8370
rect 17218 8318 17220 8370
rect 17164 7364 17220 8318
rect 17276 8260 17332 8270
rect 17276 8166 17332 8204
rect 17948 8148 18004 10782
rect 18060 10724 18116 11116
rect 18172 11106 18228 11116
rect 19068 11170 19236 11172
rect 19068 11118 19182 11170
rect 19234 11118 19236 11170
rect 19068 11116 19236 11118
rect 18060 10630 18116 10668
rect 18284 10610 18340 10622
rect 18284 10558 18286 10610
rect 18338 10558 18340 10610
rect 18284 10500 18340 10558
rect 18284 10434 18340 10444
rect 18620 10052 18676 10062
rect 18284 9940 18340 9950
rect 18060 8148 18116 8158
rect 17948 8146 18116 8148
rect 17948 8094 18062 8146
rect 18114 8094 18116 8146
rect 17948 8092 18116 8094
rect 17724 7588 17780 7598
rect 17948 7588 18004 8092
rect 18060 8082 18116 8092
rect 18284 8146 18340 9884
rect 18508 8260 18564 8270
rect 18508 8166 18564 8204
rect 18620 8258 18676 9996
rect 19068 10052 19124 11116
rect 19180 11106 19236 11116
rect 19180 10724 19236 10734
rect 19292 10724 19348 11340
rect 19180 10722 19348 10724
rect 19180 10670 19182 10722
rect 19234 10670 19348 10722
rect 19180 10668 19348 10670
rect 19516 11564 19908 11620
rect 19516 10722 19572 11564
rect 19740 11396 19796 11406
rect 19740 11302 19796 11340
rect 19852 11394 19908 11564
rect 20524 11506 20580 11900
rect 20524 11454 20526 11506
rect 20578 11454 20580 11506
rect 20524 11442 20580 11454
rect 19852 11342 19854 11394
rect 19906 11342 19908 11394
rect 19852 11330 19908 11342
rect 19516 10670 19518 10722
rect 19570 10670 19572 10722
rect 19180 10658 19236 10668
rect 19516 10658 19572 10670
rect 19628 11282 19684 11294
rect 19628 11230 19630 11282
rect 19682 11230 19684 11282
rect 19628 10610 19684 11230
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19628 10558 19630 10610
rect 19682 10558 19684 10610
rect 19292 10500 19348 10510
rect 19628 10500 19684 10558
rect 19292 10406 19348 10444
rect 19516 10444 19684 10500
rect 19068 9986 19124 9996
rect 19516 8818 19572 10444
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19516 8766 19518 8818
rect 19570 8766 19572 8818
rect 19516 8754 19572 8766
rect 19628 9042 19684 9054
rect 19628 8990 19630 9042
rect 19682 8990 19684 9042
rect 19628 8428 19684 8990
rect 20300 9044 20356 9054
rect 19628 8372 19796 8428
rect 19628 8370 19684 8372
rect 19628 8318 19630 8370
rect 19682 8318 19684 8370
rect 19628 8306 19684 8318
rect 19740 8306 19796 8316
rect 18620 8206 18622 8258
rect 18674 8206 18676 8258
rect 18284 8094 18286 8146
rect 18338 8094 18340 8146
rect 18284 7812 18340 8094
rect 17724 7586 18004 7588
rect 17724 7534 17726 7586
rect 17778 7534 18004 7586
rect 17724 7532 18004 7534
rect 18060 7756 18340 7812
rect 18060 7586 18116 7756
rect 18060 7534 18062 7586
rect 18114 7534 18116 7586
rect 17724 7522 17780 7532
rect 18060 7522 18116 7534
rect 18284 7588 18340 7598
rect 18620 7588 18676 8206
rect 19180 8260 19236 8270
rect 18284 7586 18676 7588
rect 18284 7534 18286 7586
rect 18338 7534 18676 7586
rect 18284 7532 18676 7534
rect 18844 8034 18900 8046
rect 18844 7982 18846 8034
rect 18898 7982 18900 8034
rect 18284 7522 18340 7532
rect 17836 7364 17892 7374
rect 17164 7362 17892 7364
rect 17164 7310 17838 7362
rect 17890 7310 17892 7362
rect 17164 7308 17892 7310
rect 17836 7298 17892 7308
rect 18844 5124 18900 7982
rect 19180 6914 19236 8204
rect 20076 8036 20132 8046
rect 20076 8034 20244 8036
rect 20076 7982 20078 8034
rect 20130 7982 20244 8034
rect 20076 7980 20244 7982
rect 20076 7970 20132 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 20188 7700 20244 7980
rect 20076 7644 20244 7700
rect 20076 7586 20132 7644
rect 20076 7534 20078 7586
rect 20130 7534 20132 7586
rect 20076 7522 20132 7534
rect 20300 7586 20356 8988
rect 20636 8930 20692 8942
rect 20636 8878 20638 8930
rect 20690 8878 20692 8930
rect 20412 8372 20468 8382
rect 20412 8278 20468 8316
rect 20636 8260 20692 8878
rect 20300 7534 20302 7586
rect 20354 7534 20356 7586
rect 20300 7522 20356 7534
rect 20412 7698 20468 7710
rect 20412 7646 20414 7698
rect 20466 7646 20468 7698
rect 19180 6862 19182 6914
rect 19234 6862 19236 6914
rect 19180 6850 19236 6862
rect 19404 7028 19460 7038
rect 19292 6692 19348 6702
rect 19292 6598 19348 6636
rect 18844 5058 18900 5068
rect 19292 3668 19348 3678
rect 19404 3668 19460 6972
rect 19628 6690 19684 6702
rect 19628 6638 19630 6690
rect 19682 6638 19684 6690
rect 19628 6132 19684 6638
rect 20412 6692 20468 7646
rect 20636 6916 20692 8204
rect 20748 7476 20804 7486
rect 20748 7382 20804 7420
rect 20972 7028 21028 23662
rect 21756 23938 21812 24892
rect 21868 24882 21924 24892
rect 22540 24948 22596 31276
rect 22652 31220 22708 31230
rect 22652 31126 22708 31164
rect 22764 31218 22820 31388
rect 22764 31166 22766 31218
rect 22818 31166 22820 31218
rect 22764 31154 22820 31166
rect 22876 30996 22932 31500
rect 22764 30940 22932 30996
rect 22764 30324 22820 30940
rect 22876 30770 22932 30782
rect 22876 30718 22878 30770
rect 22930 30718 22932 30770
rect 22876 30434 22932 30718
rect 22876 30382 22878 30434
rect 22930 30382 22932 30434
rect 22876 30370 22932 30382
rect 22764 30258 22820 30268
rect 22652 29988 22708 29998
rect 22652 29650 22708 29932
rect 22876 29988 22932 29998
rect 22876 29894 22932 29932
rect 22652 29598 22654 29650
rect 22706 29598 22708 29650
rect 22652 29586 22708 29598
rect 22988 26908 23044 32844
rect 23100 32450 23156 33068
rect 23548 33030 23604 33068
rect 23996 32788 24052 33852
rect 24108 33124 24164 33134
rect 24108 33030 24164 33068
rect 24108 32788 24164 32798
rect 23996 32786 24164 32788
rect 23996 32734 24110 32786
rect 24162 32734 24164 32786
rect 23996 32732 24164 32734
rect 24108 32722 24164 32732
rect 23548 32452 23604 32462
rect 23100 32398 23102 32450
rect 23154 32398 23156 32450
rect 23100 32386 23156 32398
rect 23324 32450 23604 32452
rect 23324 32398 23550 32450
rect 23602 32398 23604 32450
rect 23324 32396 23604 32398
rect 23324 32002 23380 32396
rect 23548 32386 23604 32396
rect 23324 31950 23326 32002
rect 23378 31950 23380 32002
rect 23324 31938 23380 31950
rect 23660 31780 23716 31790
rect 23660 31686 23716 31724
rect 24332 31668 24388 38220
rect 24556 38210 24612 38222
rect 24444 38052 24500 38062
rect 24444 37958 24500 37996
rect 24780 37380 24836 39452
rect 24892 37828 24948 37838
rect 24892 37734 24948 37772
rect 24780 37324 24948 37380
rect 24780 37154 24836 37166
rect 24780 37102 24782 37154
rect 24834 37102 24836 37154
rect 24556 36372 24612 36382
rect 24780 36372 24836 37102
rect 24612 36316 24836 36372
rect 24556 36240 24612 36316
rect 24668 35586 24724 36316
rect 24668 35534 24670 35586
rect 24722 35534 24724 35586
rect 24668 35476 24724 35534
rect 24668 35410 24724 35420
rect 24780 35474 24836 35486
rect 24780 35422 24782 35474
rect 24834 35422 24836 35474
rect 24780 35252 24836 35422
rect 24780 35186 24836 35196
rect 24668 34916 24724 34926
rect 24668 34822 24724 34860
rect 24556 34804 24612 34814
rect 24444 34468 24500 34478
rect 24444 34242 24500 34412
rect 24444 34190 24446 34242
rect 24498 34190 24500 34242
rect 24444 34178 24500 34190
rect 24556 34244 24612 34748
rect 24780 34802 24836 34814
rect 24780 34750 24782 34802
rect 24834 34750 24836 34802
rect 24220 31612 24388 31668
rect 24556 33122 24612 34188
rect 24668 34356 24724 34366
rect 24668 34130 24724 34300
rect 24668 34078 24670 34130
rect 24722 34078 24724 34130
rect 24668 34066 24724 34078
rect 24668 33572 24724 33582
rect 24780 33572 24836 34750
rect 24668 33570 24836 33572
rect 24668 33518 24670 33570
rect 24722 33518 24836 33570
rect 24668 33516 24836 33518
rect 24668 33506 24724 33516
rect 24556 33070 24558 33122
rect 24610 33070 24612 33122
rect 23436 31556 23492 31566
rect 23324 31554 23492 31556
rect 23324 31502 23438 31554
rect 23490 31502 23492 31554
rect 23324 31500 23492 31502
rect 23212 30770 23268 30782
rect 23212 30718 23214 30770
rect 23266 30718 23268 30770
rect 23212 30434 23268 30718
rect 23212 30382 23214 30434
rect 23266 30382 23268 30434
rect 23212 29428 23268 30382
rect 23324 30436 23380 31500
rect 23436 31490 23492 31500
rect 24108 31556 24164 31566
rect 24108 31462 24164 31500
rect 23772 31220 23828 31230
rect 23772 31126 23828 31164
rect 23436 30882 23492 30894
rect 23436 30830 23438 30882
rect 23490 30830 23492 30882
rect 23436 30770 23492 30830
rect 23436 30718 23438 30770
rect 23490 30718 23492 30770
rect 23436 30706 23492 30718
rect 23324 30380 23492 30436
rect 23324 30210 23380 30222
rect 23324 30158 23326 30210
rect 23378 30158 23380 30210
rect 23324 29988 23380 30158
rect 23436 30212 23492 30380
rect 23884 30212 23940 30222
rect 23436 30210 23940 30212
rect 23436 30158 23886 30210
rect 23938 30158 23940 30210
rect 23436 30156 23940 30158
rect 23884 30146 23940 30156
rect 23324 29922 23380 29932
rect 24220 29876 24276 31612
rect 24220 29810 24276 29820
rect 24332 30882 24388 30894
rect 24332 30830 24334 30882
rect 24386 30830 24388 30882
rect 23548 29538 23604 29550
rect 23548 29486 23550 29538
rect 23602 29486 23604 29538
rect 23324 29428 23380 29438
rect 23212 29426 23380 29428
rect 23212 29374 23326 29426
rect 23378 29374 23380 29426
rect 23212 29372 23380 29374
rect 23324 29204 23380 29372
rect 23324 29138 23380 29148
rect 23548 28980 23604 29486
rect 23996 29314 24052 29326
rect 23996 29262 23998 29314
rect 24050 29262 24052 29314
rect 23996 29204 24052 29262
rect 23996 29138 24052 29148
rect 23548 28914 23604 28924
rect 23996 28756 24052 28766
rect 23996 28082 24052 28700
rect 24332 28756 24388 30830
rect 24556 30772 24612 33070
rect 24892 33124 24948 37324
rect 25004 36258 25060 36270
rect 25004 36206 25006 36258
rect 25058 36206 25060 36258
rect 25004 35476 25060 36206
rect 25004 35410 25060 35420
rect 25228 35026 25284 41020
rect 25340 39060 25396 44156
rect 25452 42196 25508 45612
rect 25452 42130 25508 42140
rect 25452 41972 25508 41982
rect 25452 41410 25508 41916
rect 25452 41358 25454 41410
rect 25506 41358 25508 41410
rect 25452 41346 25508 41358
rect 25340 38994 25396 39004
rect 25452 40740 25508 40750
rect 25452 39730 25508 40684
rect 25452 39678 25454 39730
rect 25506 39678 25508 39730
rect 25452 37492 25508 39678
rect 25564 39284 25620 46732
rect 25676 46562 25732 46574
rect 25676 46510 25678 46562
rect 25730 46510 25732 46562
rect 25676 46004 25732 46510
rect 25676 45938 25732 45948
rect 25788 45332 25844 49868
rect 25900 49250 25956 49262
rect 25900 49198 25902 49250
rect 25954 49198 25956 49250
rect 25900 49138 25956 49198
rect 25900 49086 25902 49138
rect 25954 49086 25956 49138
rect 25900 49074 25956 49086
rect 26124 48804 26180 50092
rect 26124 48738 26180 48748
rect 26236 50594 26292 50606
rect 26236 50542 26238 50594
rect 26290 50542 26292 50594
rect 26236 50372 26292 50542
rect 26012 48468 26068 48478
rect 26012 48130 26068 48412
rect 26012 48078 26014 48130
rect 26066 48078 26068 48130
rect 26012 48020 26068 48078
rect 26012 47954 26068 47964
rect 26012 47348 26068 47358
rect 26012 47254 26068 47292
rect 26124 47236 26180 47246
rect 26124 46898 26180 47180
rect 26124 46846 26126 46898
rect 26178 46846 26180 46898
rect 26124 46834 26180 46846
rect 25676 45276 25844 45332
rect 26012 45778 26068 45790
rect 26012 45726 26014 45778
rect 26066 45726 26068 45778
rect 25676 42756 25732 45276
rect 26012 45220 26068 45726
rect 26236 45668 26292 50316
rect 26348 49028 26404 51884
rect 26796 51604 26852 52780
rect 26796 51538 26852 51548
rect 27020 52836 27076 52892
rect 27020 51828 27076 52780
rect 27132 52500 27188 52510
rect 27132 52274 27188 52444
rect 27244 52388 27300 54684
rect 27692 54628 27748 54638
rect 27692 54534 27748 54572
rect 27916 54626 27972 54638
rect 27916 54574 27918 54626
rect 27970 54574 27972 54626
rect 27356 53620 27412 53630
rect 27356 53526 27412 53564
rect 27916 53284 27972 54574
rect 28028 54516 28084 55246
rect 28252 55300 28308 56030
rect 28476 56082 28532 56094
rect 28476 56030 28478 56082
rect 28530 56030 28532 56082
rect 28028 54514 28196 54516
rect 28028 54462 28030 54514
rect 28082 54462 28196 54514
rect 28028 54460 28196 54462
rect 28028 54450 28084 54460
rect 28028 53844 28084 53854
rect 28140 53844 28196 54460
rect 28252 53954 28308 55244
rect 28252 53902 28254 53954
rect 28306 53902 28308 53954
rect 28252 53890 28308 53902
rect 28364 55970 28420 55982
rect 28364 55918 28366 55970
rect 28418 55918 28420 55970
rect 28084 53788 28196 53844
rect 28028 53712 28084 53788
rect 28364 53732 28420 55918
rect 28476 55412 28532 56030
rect 29260 55972 29316 55982
rect 29260 55878 29316 55916
rect 31612 55970 31668 55982
rect 31612 55918 31614 55970
rect 31666 55918 31668 55970
rect 30940 55858 30996 55870
rect 30940 55806 30942 55858
rect 30994 55806 30996 55858
rect 30380 55522 30436 55534
rect 30380 55470 30382 55522
rect 30434 55470 30436 55522
rect 30380 55468 30436 55470
rect 28476 55318 28532 55356
rect 30268 55412 30436 55468
rect 30940 55522 30996 55806
rect 31612 55858 31668 55918
rect 31612 55806 31614 55858
rect 31666 55806 31668 55858
rect 31612 55794 31668 55806
rect 32172 55972 32228 55982
rect 30940 55470 30942 55522
rect 30994 55470 30996 55522
rect 30940 55458 30996 55470
rect 30604 55412 30660 55422
rect 29932 55300 29988 55310
rect 29932 55206 29988 55244
rect 30156 55188 30212 55198
rect 30156 55094 30212 55132
rect 28476 55076 28532 55086
rect 28476 53954 28532 55020
rect 28924 55076 28980 55086
rect 28924 55074 29652 55076
rect 28924 55022 28926 55074
rect 28978 55022 29652 55074
rect 28924 55020 29652 55022
rect 28924 55010 28980 55020
rect 28476 53902 28478 53954
rect 28530 53902 28532 53954
rect 28476 53890 28532 53902
rect 28588 54964 28644 54974
rect 28364 53666 28420 53676
rect 27916 53218 27972 53228
rect 27916 53060 27972 53070
rect 27972 53004 28196 53060
rect 27916 52966 27972 53004
rect 27356 52946 27412 52958
rect 27356 52894 27358 52946
rect 27410 52894 27412 52946
rect 27356 52724 27412 52894
rect 27804 52948 27860 52958
rect 27804 52854 27860 52892
rect 27916 52724 27972 52734
rect 27356 52722 27972 52724
rect 27356 52670 27918 52722
rect 27970 52670 27972 52722
rect 27356 52668 27972 52670
rect 27916 52658 27972 52668
rect 27468 52500 27524 52510
rect 27244 52332 27412 52388
rect 27132 52222 27134 52274
rect 27186 52222 27188 52274
rect 27132 52210 27188 52222
rect 27244 52162 27300 52174
rect 27244 52110 27246 52162
rect 27298 52110 27300 52162
rect 26572 51380 26628 51390
rect 26572 51378 26740 51380
rect 26572 51326 26574 51378
rect 26626 51326 26740 51378
rect 26572 51324 26740 51326
rect 26572 51314 26628 51324
rect 26684 51268 26740 51324
rect 27020 51268 27076 51772
rect 26684 51266 27076 51268
rect 26684 51214 27022 51266
rect 27074 51214 27076 51266
rect 26684 51212 27076 51214
rect 26572 51154 26628 51166
rect 26572 51102 26574 51154
rect 26626 51102 26628 51154
rect 26572 50818 26628 51102
rect 26572 50766 26574 50818
rect 26626 50766 26628 50818
rect 26572 50754 26628 50766
rect 27020 50484 27076 51212
rect 27132 52052 27188 52062
rect 27132 51380 27188 51996
rect 27244 51828 27300 52110
rect 27244 51762 27300 51772
rect 27132 50820 27188 51324
rect 27244 50820 27300 50830
rect 27132 50818 27300 50820
rect 27132 50766 27246 50818
rect 27298 50766 27300 50818
rect 27132 50764 27300 50766
rect 27244 50754 27300 50764
rect 27356 50596 27412 52332
rect 27468 52386 27524 52444
rect 27468 52334 27470 52386
rect 27522 52334 27524 52386
rect 27468 52322 27524 52334
rect 27692 52164 27748 52174
rect 27580 50708 27636 50718
rect 27356 50530 27412 50540
rect 27468 50594 27524 50606
rect 27468 50542 27470 50594
rect 27522 50542 27524 50594
rect 27468 50428 27524 50542
rect 27020 50418 27076 50428
rect 26460 50370 26516 50382
rect 26460 50318 26462 50370
rect 26514 50318 26516 50370
rect 26460 49924 26516 50318
rect 26460 49858 26516 49868
rect 27132 50372 27524 50428
rect 26684 49700 26740 49710
rect 26684 49698 26852 49700
rect 26684 49646 26686 49698
rect 26738 49646 26852 49698
rect 26684 49644 26852 49646
rect 26684 49634 26740 49644
rect 26348 48972 26516 49028
rect 26348 48804 26404 48814
rect 26348 48710 26404 48748
rect 26236 45602 26292 45612
rect 26348 48244 26404 48254
rect 26012 45154 26068 45164
rect 25788 45106 25844 45118
rect 25788 45054 25790 45106
rect 25842 45054 25844 45106
rect 25788 44546 25844 45054
rect 25900 45106 25956 45118
rect 25900 45054 25902 45106
rect 25954 45054 25956 45106
rect 25900 44660 25956 45054
rect 26124 45108 26180 45118
rect 26124 45014 26180 45052
rect 26236 45106 26292 45118
rect 26236 45054 26238 45106
rect 26290 45054 26292 45106
rect 25900 44594 25956 44604
rect 25788 44494 25790 44546
rect 25842 44494 25844 44546
rect 25788 44482 25844 44494
rect 25900 44436 25956 44446
rect 25900 44342 25956 44380
rect 26236 43876 26292 45054
rect 26348 44546 26404 48188
rect 26460 47236 26516 48972
rect 26796 48916 26852 49644
rect 26908 49588 26964 49598
rect 27132 49588 27188 50372
rect 27244 50036 27300 50046
rect 27580 50036 27636 50652
rect 27244 50034 27636 50036
rect 27244 49982 27246 50034
rect 27298 49982 27636 50034
rect 27244 49980 27636 49982
rect 27692 50484 27748 52108
rect 28140 51492 28196 53004
rect 28476 52836 28532 52846
rect 28476 52742 28532 52780
rect 27916 51378 27972 51390
rect 27916 51326 27918 51378
rect 27970 51326 27972 51378
rect 27916 50818 27972 51326
rect 27916 50766 27918 50818
rect 27970 50766 27972 50818
rect 27916 50754 27972 50766
rect 27804 50484 27860 50494
rect 28028 50484 28084 50494
rect 27692 50428 27804 50484
rect 27244 49970 27300 49980
rect 26908 49586 27188 49588
rect 26908 49534 26910 49586
rect 26962 49534 27188 49586
rect 26908 49532 27188 49534
rect 26908 49522 26964 49532
rect 26908 48916 26964 48926
rect 26796 48914 26964 48916
rect 26796 48862 26910 48914
rect 26962 48862 26964 48914
rect 26796 48860 26964 48862
rect 26684 48242 26740 48254
rect 26684 48190 26686 48242
rect 26738 48190 26740 48242
rect 26684 48132 26740 48190
rect 26684 48066 26740 48076
rect 26572 48020 26628 48030
rect 26572 47572 26628 47964
rect 26572 47458 26628 47516
rect 26572 47406 26574 47458
rect 26626 47406 26628 47458
rect 26572 47394 26628 47406
rect 26460 47180 26628 47236
rect 26348 44494 26350 44546
rect 26402 44494 26404 44546
rect 26348 44434 26404 44494
rect 26348 44382 26350 44434
rect 26402 44382 26404 44434
rect 26348 44370 26404 44382
rect 26460 44660 26516 44670
rect 26460 44212 26516 44604
rect 26460 44146 26516 44156
rect 26236 43820 26404 43876
rect 26348 43650 26404 43820
rect 26348 43598 26350 43650
rect 26402 43598 26404 43650
rect 26348 43586 26404 43598
rect 25900 43428 25956 43438
rect 25900 43334 25956 43372
rect 26348 43428 26404 43438
rect 26012 43314 26068 43326
rect 26236 43316 26292 43326
rect 26012 43262 26014 43314
rect 26066 43262 26068 43314
rect 26012 42868 26068 43262
rect 26012 42774 26068 42812
rect 26124 43314 26292 43316
rect 26124 43262 26238 43314
rect 26290 43262 26292 43314
rect 26124 43260 26292 43262
rect 25676 42690 25732 42700
rect 25788 42756 25844 42766
rect 25788 42754 25956 42756
rect 25788 42702 25790 42754
rect 25842 42702 25956 42754
rect 25788 42700 25956 42702
rect 25788 42690 25844 42700
rect 25900 42644 25956 42700
rect 26124 42644 26180 43260
rect 26236 43250 26292 43260
rect 26236 42980 26292 42990
rect 26348 42980 26404 43372
rect 26236 42978 26404 42980
rect 26236 42926 26238 42978
rect 26290 42926 26404 42978
rect 26236 42924 26404 42926
rect 26236 42914 26292 42924
rect 25900 42588 26180 42644
rect 25788 42082 25844 42094
rect 25788 42030 25790 42082
rect 25842 42030 25844 42082
rect 25676 41972 25732 41982
rect 25676 41878 25732 41916
rect 25788 41300 25844 42030
rect 25788 41234 25844 41244
rect 25788 41076 25844 41086
rect 25900 41076 25956 42588
rect 26460 42196 26516 42206
rect 26012 42084 26068 42094
rect 26012 41990 26068 42028
rect 26460 42082 26516 42140
rect 26460 42030 26462 42082
rect 26514 42030 26516 42082
rect 26460 42018 26516 42030
rect 26572 41748 26628 47180
rect 26684 46564 26740 46574
rect 26796 46564 26852 48860
rect 26908 48850 26964 48860
rect 26908 48132 26964 48142
rect 26908 46674 26964 48076
rect 27020 48020 27076 49532
rect 27692 49140 27748 50428
rect 27804 50352 27860 50428
rect 27916 50482 28084 50484
rect 27916 50430 28030 50482
rect 28082 50430 28084 50482
rect 27916 50428 28084 50430
rect 27804 49924 27860 49934
rect 27804 49830 27860 49868
rect 27244 49138 27748 49140
rect 27244 49086 27694 49138
rect 27746 49086 27748 49138
rect 27244 49084 27748 49086
rect 27916 49140 27972 50428
rect 28028 50418 28084 50428
rect 28028 50036 28084 50046
rect 28140 50036 28196 51436
rect 28476 52052 28532 52062
rect 28588 52052 28644 54908
rect 28700 54514 28756 54526
rect 28700 54462 28702 54514
rect 28754 54462 28756 54514
rect 28700 54404 28756 54462
rect 28700 54338 28756 54348
rect 29148 54514 29204 54526
rect 29148 54462 29150 54514
rect 29202 54462 29204 54514
rect 29148 54404 29204 54462
rect 29148 54338 29204 54348
rect 28700 53956 28756 53966
rect 28700 52722 28756 53900
rect 28924 53956 28980 53966
rect 28924 53862 28980 53900
rect 29596 53732 29652 55020
rect 29708 55074 29764 55086
rect 29708 55022 29710 55074
rect 29762 55022 29764 55074
rect 29708 54964 29764 55022
rect 30044 55076 30100 55086
rect 30044 54982 30100 55020
rect 29708 54898 29764 54908
rect 29932 54404 29988 54414
rect 29932 54310 29988 54348
rect 29820 53732 29876 53742
rect 29596 53730 29876 53732
rect 29596 53678 29822 53730
rect 29874 53678 29876 53730
rect 29596 53676 29876 53678
rect 29820 53666 29876 53676
rect 30156 53732 30212 53742
rect 30156 53638 30212 53676
rect 28700 52670 28702 52722
rect 28754 52670 28756 52722
rect 28700 52658 28756 52670
rect 28924 52834 28980 52846
rect 28924 52782 28926 52834
rect 28978 52782 28980 52834
rect 28924 52612 28980 52782
rect 29372 52836 29428 52846
rect 29372 52742 29428 52780
rect 29820 52834 29876 52846
rect 29820 52782 29822 52834
rect 29874 52782 29876 52834
rect 28924 52546 28980 52556
rect 29148 52722 29204 52734
rect 29148 52670 29150 52722
rect 29202 52670 29204 52722
rect 28476 52050 28644 52052
rect 28476 51998 28478 52050
rect 28530 51998 28644 52050
rect 28476 51996 28644 51998
rect 28476 51490 28532 51996
rect 28476 51438 28478 51490
rect 28530 51438 28532 51490
rect 28476 51426 28532 51438
rect 28812 51938 28868 51950
rect 28812 51886 28814 51938
rect 28866 51886 28868 51938
rect 28364 51380 28420 51390
rect 28364 51286 28420 51324
rect 28028 50034 28196 50036
rect 28028 49982 28030 50034
rect 28082 49982 28196 50034
rect 28028 49980 28196 49982
rect 28252 51266 28308 51278
rect 28252 51214 28254 51266
rect 28306 51214 28308 51266
rect 28252 50036 28308 51214
rect 28812 50708 28868 51886
rect 28812 50642 28868 50652
rect 28476 50484 28532 50494
rect 28476 50390 28532 50428
rect 28028 49970 28084 49980
rect 28252 49970 28308 49980
rect 28364 50372 28420 50382
rect 28364 50034 28420 50316
rect 28364 49982 28366 50034
rect 28418 49982 28420 50034
rect 28364 49970 28420 49982
rect 28252 49810 28308 49822
rect 28252 49758 28254 49810
rect 28306 49758 28308 49810
rect 28252 49476 28308 49758
rect 28364 49812 28420 49822
rect 28364 49698 28420 49756
rect 28364 49646 28366 49698
rect 28418 49646 28420 49698
rect 28364 49634 28420 49646
rect 28924 49698 28980 49710
rect 28924 49646 28926 49698
rect 28978 49646 28980 49698
rect 28252 49410 28308 49420
rect 28924 49476 28980 49646
rect 28252 49140 28308 49150
rect 27916 49084 28252 49140
rect 27244 48914 27300 49084
rect 27692 49074 27748 49084
rect 28252 49008 28308 49084
rect 28924 49028 28980 49420
rect 28924 48962 28980 48972
rect 29036 49140 29092 49150
rect 27244 48862 27246 48914
rect 27298 48862 27300 48914
rect 27132 48468 27188 48478
rect 27244 48468 27300 48862
rect 27132 48466 27300 48468
rect 27132 48414 27134 48466
rect 27186 48414 27300 48466
rect 27132 48412 27300 48414
rect 27468 48916 27524 48926
rect 27132 48244 27188 48412
rect 27132 48178 27188 48188
rect 27356 48242 27412 48254
rect 27356 48190 27358 48242
rect 27410 48190 27412 48242
rect 27244 48130 27300 48142
rect 27244 48078 27246 48130
rect 27298 48078 27300 48130
rect 27020 47964 27188 48020
rect 27132 47570 27188 47964
rect 27132 47518 27134 47570
rect 27186 47518 27188 47570
rect 27132 47506 27188 47518
rect 26908 46622 26910 46674
rect 26962 46622 26964 46674
rect 26908 46610 26964 46622
rect 27020 47458 27076 47470
rect 27020 47406 27022 47458
rect 27074 47406 27076 47458
rect 26684 46562 26852 46564
rect 26684 46510 26686 46562
rect 26738 46510 26852 46562
rect 26684 46508 26852 46510
rect 26684 46498 26740 46508
rect 26684 45332 26740 45342
rect 26684 45106 26740 45276
rect 26684 45054 26686 45106
rect 26738 45054 26740 45106
rect 26684 44436 26740 45054
rect 26684 44370 26740 44380
rect 26684 44212 26740 44222
rect 26684 44118 26740 44156
rect 26684 43652 26740 43662
rect 26684 42978 26740 43596
rect 26684 42926 26686 42978
rect 26738 42926 26740 42978
rect 26684 42914 26740 42926
rect 26796 42308 26852 46508
rect 27020 46452 27076 47406
rect 27244 47460 27300 48078
rect 27244 47394 27300 47404
rect 27356 47012 27412 48190
rect 27132 46956 27412 47012
rect 27132 46674 27188 46956
rect 27356 46788 27412 46956
rect 27356 46722 27412 46732
rect 27132 46622 27134 46674
rect 27186 46622 27188 46674
rect 27132 46610 27188 46622
rect 27020 46116 27076 46396
rect 27244 46340 27300 46350
rect 27020 46060 27188 46116
rect 27020 45668 27076 45678
rect 27020 45574 27076 45612
rect 27132 45332 27188 46060
rect 27020 45276 27188 45332
rect 26908 44996 26964 45006
rect 26908 44902 26964 44940
rect 27020 43652 27076 45276
rect 27132 45108 27188 45118
rect 27132 45014 27188 45052
rect 27132 44660 27188 44670
rect 27132 44434 27188 44604
rect 27132 44382 27134 44434
rect 27186 44382 27188 44434
rect 27132 44370 27188 44382
rect 27244 44212 27300 46284
rect 27356 45220 27412 45230
rect 27356 45126 27412 45164
rect 27020 43586 27076 43596
rect 27132 44156 27300 44212
rect 26796 42242 26852 42252
rect 27020 43316 27076 43326
rect 26684 42084 26740 42094
rect 26684 41990 26740 42028
rect 26908 42084 26964 42094
rect 26908 41990 26964 42028
rect 27020 42082 27076 43260
rect 27020 42030 27022 42082
rect 27074 42030 27076 42082
rect 26460 41692 26628 41748
rect 27020 41972 27076 42030
rect 26348 41300 26404 41310
rect 26460 41300 26516 41692
rect 27020 41412 27076 41916
rect 27020 41346 27076 41356
rect 26460 41244 26628 41300
rect 26348 41206 26404 41244
rect 25844 41020 25956 41076
rect 25788 40982 25844 41020
rect 26124 40740 26180 40750
rect 25900 40628 25956 40638
rect 25900 39730 25956 40572
rect 25900 39678 25902 39730
rect 25954 39678 25956 39730
rect 25900 39508 25956 39678
rect 25900 39442 25956 39452
rect 26012 40290 26068 40302
rect 26012 40238 26014 40290
rect 26066 40238 26068 40290
rect 25564 39228 25956 39284
rect 25676 39060 25732 39070
rect 25564 38724 25620 38734
rect 25564 38050 25620 38668
rect 25564 37998 25566 38050
rect 25618 37998 25620 38050
rect 25564 37986 25620 37998
rect 25452 37436 25620 37492
rect 25564 37156 25620 37436
rect 25676 37380 25732 39004
rect 25788 38836 25844 38846
rect 25788 38742 25844 38780
rect 25900 38668 25956 39228
rect 26012 38948 26068 40238
rect 26124 40178 26180 40684
rect 26348 40628 26404 40638
rect 26348 40534 26404 40572
rect 26124 40126 26126 40178
rect 26178 40126 26180 40178
rect 26124 40114 26180 40126
rect 26012 38882 26068 38892
rect 26460 39618 26516 39630
rect 26460 39566 26462 39618
rect 26514 39566 26516 39618
rect 26460 38836 26516 39566
rect 26460 38770 26516 38780
rect 26348 38722 26404 38734
rect 26348 38670 26350 38722
rect 26402 38670 26404 38722
rect 26348 38668 26404 38670
rect 25900 38612 26180 38668
rect 26348 38612 26516 38668
rect 26012 38388 26068 38398
rect 25788 37828 25844 37838
rect 25788 37734 25844 37772
rect 25676 37324 25844 37380
rect 25676 37156 25732 37166
rect 25564 37154 25732 37156
rect 25564 37102 25678 37154
rect 25730 37102 25732 37154
rect 25564 37100 25732 37102
rect 25676 36596 25732 37100
rect 25676 36530 25732 36540
rect 25452 36260 25508 36270
rect 25452 36166 25508 36204
rect 25564 35586 25620 35598
rect 25564 35534 25566 35586
rect 25618 35534 25620 35586
rect 25564 35476 25620 35534
rect 25564 35410 25620 35420
rect 25788 35140 25844 37324
rect 25228 34974 25230 35026
rect 25282 34974 25284 35026
rect 25228 34356 25284 34974
rect 25228 34290 25284 34300
rect 25340 35084 25844 35140
rect 26012 35922 26068 38332
rect 26012 35870 26014 35922
rect 26066 35870 26068 35922
rect 24892 33058 24948 33068
rect 25340 32788 25396 35084
rect 26012 35028 26068 35870
rect 25788 34972 26012 35028
rect 25788 34914 25844 34972
rect 26012 34962 26068 34972
rect 25788 34862 25790 34914
rect 25842 34862 25844 34914
rect 25788 34850 25844 34862
rect 25564 34356 25620 34366
rect 25564 34262 25620 34300
rect 26012 34018 26068 34030
rect 26012 33966 26014 34018
rect 26066 33966 26068 34018
rect 26012 33796 26068 33966
rect 26012 33730 26068 33740
rect 25228 32732 25396 32788
rect 25452 33346 25508 33358
rect 25452 33294 25454 33346
rect 25506 33294 25508 33346
rect 24556 30706 24612 30716
rect 25004 32340 25060 32350
rect 24332 28690 24388 28700
rect 24892 29988 24948 29998
rect 24892 29314 24948 29932
rect 24892 29262 24894 29314
rect 24946 29262 24948 29314
rect 23996 28030 23998 28082
rect 24050 28030 24052 28082
rect 23996 28018 24052 28030
rect 24780 27636 24836 27646
rect 24780 27542 24836 27580
rect 22540 24882 22596 24892
rect 22652 26852 23044 26908
rect 23772 26964 23828 26974
rect 22540 24276 22596 24286
rect 22540 24050 22596 24220
rect 22540 23998 22542 24050
rect 22594 23998 22596 24050
rect 22540 23986 22596 23998
rect 21756 23886 21758 23938
rect 21810 23886 21812 23938
rect 21756 23604 21812 23886
rect 21980 23716 22036 23726
rect 21980 23622 22036 23660
rect 21756 23538 21812 23548
rect 21308 23492 21364 23502
rect 21308 23266 21364 23436
rect 21308 23214 21310 23266
rect 21362 23214 21364 23266
rect 21308 23202 21364 23214
rect 22092 22260 22148 22270
rect 21980 22258 22148 22260
rect 21980 22206 22094 22258
rect 22146 22206 22148 22258
rect 21980 22204 22148 22206
rect 21756 21476 21812 21486
rect 21756 21382 21812 21420
rect 21756 20914 21812 20926
rect 21756 20862 21758 20914
rect 21810 20862 21812 20914
rect 21644 19124 21700 19134
rect 21644 19030 21700 19068
rect 21308 18900 21364 18910
rect 21196 18452 21252 18462
rect 21196 18358 21252 18396
rect 21308 17556 21364 18844
rect 21756 18676 21812 20862
rect 21532 18620 21812 18676
rect 21868 19122 21924 19134
rect 21868 19070 21870 19122
rect 21922 19070 21924 19122
rect 21196 17500 21364 17556
rect 21420 17668 21476 17678
rect 21196 13188 21252 17500
rect 21308 16884 21364 16894
rect 21308 16790 21364 16828
rect 21420 15426 21476 17612
rect 21532 16212 21588 18620
rect 21644 18452 21700 18462
rect 21868 18452 21924 19070
rect 21644 18450 21924 18452
rect 21644 18398 21646 18450
rect 21698 18398 21924 18450
rect 21644 18396 21924 18398
rect 21980 18452 22036 22204
rect 22092 22194 22148 22204
rect 22428 22260 22484 22270
rect 22652 22260 22708 26852
rect 22876 24834 22932 24846
rect 22876 24782 22878 24834
rect 22930 24782 22932 24834
rect 22428 22258 22708 22260
rect 22428 22206 22430 22258
rect 22482 22206 22708 22258
rect 22428 22204 22708 22206
rect 22764 24276 22820 24286
rect 22428 22194 22484 22204
rect 22652 21700 22708 21710
rect 22428 21588 22484 21598
rect 22428 21494 22484 21532
rect 22652 21586 22708 21644
rect 22652 21534 22654 21586
rect 22706 21534 22708 21586
rect 22652 21522 22708 21534
rect 22316 21476 22372 21486
rect 22204 20914 22260 20926
rect 22204 20862 22206 20914
rect 22258 20862 22260 20914
rect 22204 19908 22260 20862
rect 22204 19842 22260 19852
rect 22204 19122 22260 19134
rect 22204 19070 22206 19122
rect 22258 19070 22260 19122
rect 22092 19012 22148 19022
rect 22092 18918 22148 18956
rect 22092 18452 22148 18462
rect 21980 18450 22148 18452
rect 21980 18398 22094 18450
rect 22146 18398 22148 18450
rect 21980 18396 22148 18398
rect 21644 17554 21700 18396
rect 22092 18386 22148 18396
rect 22204 18452 22260 19070
rect 22204 18386 22260 18396
rect 21644 17502 21646 17554
rect 21698 17502 21700 17554
rect 21644 16882 21700 17502
rect 22092 17444 22148 17454
rect 21644 16830 21646 16882
rect 21698 16830 21700 16882
rect 21644 16818 21700 16830
rect 21868 16884 21924 16894
rect 21532 16080 21588 16156
rect 21420 15374 21422 15426
rect 21474 15374 21476 15426
rect 21420 15362 21476 15374
rect 21532 14644 21588 14654
rect 21532 14530 21588 14588
rect 21868 14642 21924 16828
rect 21980 15874 22036 15886
rect 21980 15822 21982 15874
rect 22034 15822 22036 15874
rect 21980 15764 22036 15822
rect 21980 15698 22036 15708
rect 21868 14590 21870 14642
rect 21922 14590 21924 14642
rect 21868 14578 21924 14590
rect 21532 14478 21534 14530
rect 21586 14478 21588 14530
rect 21532 14466 21588 14478
rect 21980 13746 22036 13758
rect 21980 13694 21982 13746
rect 22034 13694 22036 13746
rect 21980 13636 22036 13694
rect 21980 13570 22036 13580
rect 21196 13132 21588 13188
rect 21196 13076 21252 13132
rect 21196 13010 21252 13020
rect 21532 13074 21588 13132
rect 21532 13022 21534 13074
rect 21586 13022 21588 13074
rect 21532 13010 21588 13022
rect 21196 12628 21252 12638
rect 21196 12178 21252 12572
rect 21196 12126 21198 12178
rect 21250 12126 21252 12178
rect 21196 12114 21252 12126
rect 21868 12628 21924 12638
rect 21868 11506 21924 12572
rect 21980 12180 22036 12190
rect 21980 12086 22036 12124
rect 21868 11454 21870 11506
rect 21922 11454 21924 11506
rect 21868 11442 21924 11454
rect 21084 9940 21140 9950
rect 21084 9044 21140 9884
rect 21532 9940 21588 9950
rect 21532 9846 21588 9884
rect 21756 9940 21812 9950
rect 21084 8912 21140 8988
rect 21644 8034 21700 8046
rect 21644 7982 21646 8034
rect 21698 7982 21700 8034
rect 21644 7476 21700 7982
rect 21644 7410 21700 7420
rect 20972 6962 21028 6972
rect 21420 7362 21476 7374
rect 21420 7310 21422 7362
rect 21474 7310 21476 7362
rect 20636 6860 20916 6916
rect 20860 6804 20916 6860
rect 20972 6804 21028 6814
rect 20860 6802 21028 6804
rect 20860 6750 20974 6802
rect 21026 6750 21028 6802
rect 20860 6748 21028 6750
rect 20972 6738 21028 6748
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19628 6066 19684 6076
rect 20412 6018 20468 6636
rect 20636 6132 20692 6142
rect 20636 6038 20692 6076
rect 21420 6132 21476 7310
rect 21644 6804 21700 6814
rect 21756 6804 21812 9884
rect 21980 9268 22036 9278
rect 22092 9268 22148 17388
rect 22316 14532 22372 21420
rect 22540 21476 22596 21486
rect 22540 20802 22596 21420
rect 22540 20750 22542 20802
rect 22594 20750 22596 20802
rect 22540 20738 22596 20750
rect 22428 19906 22484 19918
rect 22428 19854 22430 19906
rect 22482 19854 22484 19906
rect 22428 19012 22484 19854
rect 22652 19012 22708 19022
rect 22428 19010 22708 19012
rect 22428 18958 22654 19010
rect 22706 18958 22708 19010
rect 22428 18956 22708 18958
rect 22652 18452 22708 18956
rect 22764 18564 22820 24220
rect 22876 24052 22932 24782
rect 23212 24276 23268 24286
rect 23100 24052 23156 24062
rect 22876 24050 23156 24052
rect 22876 23998 23102 24050
rect 23154 23998 23156 24050
rect 22876 23996 23156 23998
rect 23100 23986 23156 23996
rect 23212 23938 23268 24220
rect 23212 23886 23214 23938
rect 23266 23886 23268 23938
rect 23212 23874 23268 23886
rect 22988 23828 23044 23838
rect 22988 23734 23044 23772
rect 23548 23828 23604 23838
rect 23548 23826 23716 23828
rect 23548 23774 23550 23826
rect 23602 23774 23716 23826
rect 23548 23772 23716 23774
rect 23548 23762 23604 23772
rect 23100 23716 23156 23726
rect 22988 22146 23044 22158
rect 22988 22094 22990 22146
rect 23042 22094 23044 22146
rect 22988 21588 23044 22094
rect 23100 22036 23156 23660
rect 23660 23156 23716 23772
rect 23772 23378 23828 26908
rect 24556 26964 24612 27002
rect 24556 26898 24612 26908
rect 24444 26852 24500 26862
rect 24444 26514 24500 26796
rect 24892 26852 24948 29262
rect 25004 26908 25060 32284
rect 25116 28530 25172 28542
rect 25116 28478 25118 28530
rect 25170 28478 25172 28530
rect 25116 28084 25172 28478
rect 25116 28018 25172 28028
rect 25004 26852 25172 26908
rect 24892 26758 24948 26796
rect 24444 26462 24446 26514
rect 24498 26462 24500 26514
rect 24444 26450 24500 26462
rect 25004 26628 25060 26638
rect 25004 26514 25060 26572
rect 25004 26462 25006 26514
rect 25058 26462 25060 26514
rect 25004 26450 25060 26462
rect 24668 25394 24724 25406
rect 24668 25342 24670 25394
rect 24722 25342 24724 25394
rect 24108 25282 24164 25294
rect 24108 25230 24110 25282
rect 24162 25230 24164 25282
rect 24108 25172 24164 25230
rect 24108 23716 24164 25116
rect 24668 25172 24724 25342
rect 24668 25106 24724 25116
rect 24668 24836 24724 24846
rect 24668 24742 24724 24780
rect 24892 24612 24948 24622
rect 24332 24052 24388 24062
rect 24332 23958 24388 23996
rect 24108 23650 24164 23660
rect 23772 23326 23774 23378
rect 23826 23326 23828 23378
rect 23772 23314 23828 23326
rect 24668 23604 24724 23614
rect 24668 23378 24724 23548
rect 24668 23326 24670 23378
rect 24722 23326 24724 23378
rect 23660 23100 24612 23156
rect 24556 23042 24612 23100
rect 24556 22990 24558 23042
rect 24610 22990 24612 23042
rect 24556 22978 24612 22990
rect 23212 22484 23268 22494
rect 23212 22258 23268 22428
rect 23772 22484 23828 22494
rect 24668 22484 24724 23326
rect 24892 23266 24948 24556
rect 25116 24388 25172 26852
rect 25116 24322 25172 24332
rect 25228 24164 25284 32732
rect 25452 32676 25508 33294
rect 25900 33346 25956 33358
rect 25900 33294 25902 33346
rect 25954 33294 25956 33346
rect 25676 32676 25732 32686
rect 25452 32674 25732 32676
rect 25452 32622 25678 32674
rect 25730 32622 25732 32674
rect 25452 32620 25732 32622
rect 25676 32564 25732 32620
rect 25676 32498 25732 32508
rect 25900 31892 25956 33294
rect 26012 32676 26068 32686
rect 26012 32582 26068 32620
rect 25900 31826 25956 31836
rect 26124 29652 26180 38612
rect 26460 37826 26516 38612
rect 26572 38388 26628 41244
rect 27132 41188 27188 44156
rect 27244 43652 27300 43662
rect 27244 43558 27300 43596
rect 27356 43650 27412 43662
rect 27356 43598 27358 43650
rect 27410 43598 27412 43650
rect 27356 42980 27412 43598
rect 27468 43092 27524 48860
rect 28812 48804 28868 48814
rect 28700 48802 28868 48804
rect 28700 48750 28814 48802
rect 28866 48750 28868 48802
rect 28700 48748 28868 48750
rect 27916 48130 27972 48142
rect 27916 48078 27918 48130
rect 27970 48078 27972 48130
rect 27916 48020 27972 48078
rect 28588 48132 28644 48142
rect 28700 48132 28756 48748
rect 28812 48738 28868 48748
rect 29036 48468 29092 49084
rect 28588 48130 28756 48132
rect 28588 48078 28590 48130
rect 28642 48078 28756 48130
rect 28588 48076 28756 48078
rect 28588 48066 28644 48076
rect 27916 47954 27972 47964
rect 28700 48018 28756 48076
rect 28700 47966 28702 48018
rect 28754 47966 28756 48018
rect 28700 47954 28756 47966
rect 28812 48466 29092 48468
rect 28812 48414 29038 48466
rect 29090 48414 29092 48466
rect 28812 48412 29092 48414
rect 28588 47908 28644 47918
rect 28476 47796 28532 47806
rect 28476 47570 28532 47740
rect 28476 47518 28478 47570
rect 28530 47518 28532 47570
rect 28476 47506 28532 47518
rect 28140 47460 28196 47470
rect 28140 47366 28196 47404
rect 27580 47346 27636 47358
rect 27580 47294 27582 47346
rect 27634 47294 27636 47346
rect 27580 47124 27636 47294
rect 28476 47236 28532 47246
rect 27580 47058 27636 47068
rect 27692 47234 28532 47236
rect 27692 47182 28478 47234
rect 28530 47182 28532 47234
rect 27692 47180 28532 47182
rect 27580 46900 27636 46910
rect 27692 46900 27748 47180
rect 28476 47170 28532 47180
rect 27580 46898 27748 46900
rect 27580 46846 27582 46898
rect 27634 46846 27748 46898
rect 27580 46844 27748 46846
rect 28140 47012 28196 47022
rect 27580 46834 27636 46844
rect 28028 46788 28084 46798
rect 28028 46694 28084 46732
rect 28140 46674 28196 46956
rect 28588 46676 28644 47852
rect 28812 47460 28868 48412
rect 29036 48402 29092 48412
rect 28700 47404 28980 47460
rect 28700 47346 28756 47404
rect 28700 47294 28702 47346
rect 28754 47294 28756 47346
rect 28700 47282 28756 47294
rect 28140 46622 28142 46674
rect 28194 46622 28196 46674
rect 28140 46610 28196 46622
rect 28252 46674 28644 46676
rect 28252 46622 28590 46674
rect 28642 46622 28644 46674
rect 28252 46620 28644 46622
rect 28252 46116 28308 46620
rect 28588 46610 28644 46620
rect 28364 46452 28420 46462
rect 28364 46358 28420 46396
rect 27580 46060 28308 46116
rect 27580 46002 27636 46060
rect 27580 45950 27582 46002
rect 27634 45950 27636 46002
rect 27580 45938 27636 45950
rect 28140 45332 28196 46060
rect 28252 45666 28308 45678
rect 28252 45614 28254 45666
rect 28306 45614 28308 45666
rect 28252 45556 28308 45614
rect 28252 45490 28308 45500
rect 28700 45666 28756 45678
rect 28700 45614 28702 45666
rect 28754 45614 28756 45666
rect 28196 45276 28308 45332
rect 28140 45266 28196 45276
rect 28028 45220 28084 45230
rect 28028 45126 28084 45164
rect 27916 45106 27972 45118
rect 27916 45054 27918 45106
rect 27970 45054 27972 45106
rect 27916 44884 27972 45054
rect 28140 45108 28196 45118
rect 28140 45014 28196 45052
rect 28252 44884 28308 45276
rect 28588 45108 28644 45118
rect 28700 45108 28756 45614
rect 28588 45106 28756 45108
rect 28588 45054 28590 45106
rect 28642 45054 28756 45106
rect 28588 45052 28756 45054
rect 28588 45042 28644 45052
rect 27916 44828 28308 44884
rect 27692 44660 27748 44670
rect 27692 44210 27748 44604
rect 27692 44158 27694 44210
rect 27746 44158 27748 44210
rect 27692 43988 27748 44158
rect 27692 43922 27748 43932
rect 28028 44322 28084 44334
rect 28588 44324 28644 44334
rect 28028 44270 28030 44322
rect 28082 44270 28084 44322
rect 27580 43764 27636 43774
rect 28028 43764 28084 44270
rect 27580 43762 28084 43764
rect 27580 43710 27582 43762
rect 27634 43710 28030 43762
rect 28082 43710 28084 43762
rect 27580 43708 28084 43710
rect 27580 43698 27636 43708
rect 28028 43698 28084 43708
rect 28140 44322 28644 44324
rect 28140 44270 28590 44322
rect 28642 44270 28644 44322
rect 28140 44268 28644 44270
rect 28140 43650 28196 44268
rect 28588 44258 28644 44268
rect 28588 44100 28644 44110
rect 28476 44098 28644 44100
rect 28476 44046 28590 44098
rect 28642 44046 28644 44098
rect 28476 44044 28644 44046
rect 28252 43988 28308 43998
rect 28252 43762 28308 43932
rect 28252 43710 28254 43762
rect 28306 43710 28308 43762
rect 28252 43698 28308 43710
rect 28140 43598 28142 43650
rect 28194 43598 28196 43650
rect 28140 43586 28196 43598
rect 27468 43036 27972 43092
rect 27356 42978 27524 42980
rect 27356 42926 27358 42978
rect 27410 42926 27524 42978
rect 27356 42924 27524 42926
rect 27356 42914 27412 42924
rect 27020 41132 27188 41188
rect 27356 42530 27412 42542
rect 27356 42478 27358 42530
rect 27410 42478 27412 42530
rect 26796 40628 26852 40638
rect 26796 40534 26852 40572
rect 26684 39506 26740 39518
rect 26684 39454 26686 39506
rect 26738 39454 26740 39506
rect 26684 38948 26740 39454
rect 26684 38882 26740 38892
rect 26572 38322 26628 38332
rect 26684 38276 26740 38286
rect 26684 38182 26740 38220
rect 26572 38052 26628 38062
rect 26572 37958 26628 37996
rect 26460 37774 26462 37826
rect 26514 37774 26516 37826
rect 26236 37268 26292 37278
rect 26236 37174 26292 37212
rect 26460 37044 26516 37774
rect 26684 37828 26740 37838
rect 26684 37266 26740 37772
rect 26684 37214 26686 37266
rect 26738 37214 26740 37266
rect 26684 37156 26740 37214
rect 26684 37090 26740 37100
rect 26460 36978 26516 36988
rect 26908 37042 26964 37054
rect 26908 36990 26910 37042
rect 26962 36990 26964 37042
rect 26236 36932 26292 36942
rect 26236 36596 26292 36876
rect 26236 36502 26292 36540
rect 26908 36932 26964 36990
rect 26908 36482 26964 36876
rect 26908 36430 26910 36482
rect 26962 36430 26964 36482
rect 26908 36418 26964 36430
rect 26348 35252 26404 35262
rect 27020 35252 27076 41132
rect 26348 35026 26404 35196
rect 26348 34974 26350 35026
rect 26402 34974 26404 35026
rect 26348 34962 26404 34974
rect 26572 35196 27076 35252
rect 27132 40964 27188 40974
rect 27356 40964 27412 42478
rect 27468 41412 27524 42924
rect 27916 42644 27972 43036
rect 28028 42980 28084 42990
rect 28028 42978 28420 42980
rect 28028 42926 28030 42978
rect 28082 42926 28420 42978
rect 28028 42924 28420 42926
rect 28028 42914 28084 42924
rect 27916 42588 28196 42644
rect 27692 42530 27748 42542
rect 27692 42478 27694 42530
rect 27746 42478 27748 42530
rect 27580 42196 27636 42206
rect 27692 42196 27748 42478
rect 28028 42420 28084 42430
rect 27692 42140 27972 42196
rect 27580 42102 27636 42140
rect 27804 41972 27860 41982
rect 27692 41970 27860 41972
rect 27692 41918 27806 41970
rect 27858 41918 27860 41970
rect 27692 41916 27860 41918
rect 27580 41412 27636 41422
rect 27468 41410 27636 41412
rect 27468 41358 27582 41410
rect 27634 41358 27636 41410
rect 27468 41356 27636 41358
rect 27580 41346 27636 41356
rect 27692 41074 27748 41916
rect 27804 41906 27860 41916
rect 27916 41972 27972 42140
rect 27916 41906 27972 41916
rect 28028 41748 28084 42364
rect 27692 41022 27694 41074
rect 27746 41022 27748 41074
rect 27692 40964 27748 41022
rect 27132 40962 27748 40964
rect 27132 40910 27134 40962
rect 27186 40910 27748 40962
rect 27132 40908 27748 40910
rect 27804 41692 28084 41748
rect 26572 34914 26628 35196
rect 26908 35028 26964 35038
rect 26908 34934 26964 34972
rect 26572 34862 26574 34914
rect 26626 34862 26628 34914
rect 26572 33796 26628 34862
rect 26572 33730 26628 33740
rect 26908 34132 26964 34142
rect 26908 32786 26964 34076
rect 27132 33684 27188 40908
rect 27356 40740 27412 40750
rect 27356 40628 27412 40684
rect 27356 40626 27524 40628
rect 27356 40574 27358 40626
rect 27410 40574 27524 40626
rect 27356 40572 27524 40574
rect 27356 40562 27412 40572
rect 27244 40178 27300 40190
rect 27244 40126 27246 40178
rect 27298 40126 27300 40178
rect 27244 39618 27300 40126
rect 27244 39566 27246 39618
rect 27298 39566 27300 39618
rect 27244 39554 27300 39566
rect 27356 38836 27412 38846
rect 27356 38742 27412 38780
rect 27244 38276 27300 38286
rect 27244 37490 27300 38220
rect 27356 38052 27412 38062
rect 27356 37958 27412 37996
rect 27244 37438 27246 37490
rect 27298 37438 27300 37490
rect 27244 37426 27300 37438
rect 27468 37380 27524 40572
rect 27692 39618 27748 39630
rect 27692 39566 27694 39618
rect 27746 39566 27748 39618
rect 27692 39508 27748 39566
rect 27580 38948 27636 38958
rect 27580 38050 27636 38892
rect 27692 38834 27748 39452
rect 27804 39506 27860 41692
rect 27804 39454 27806 39506
rect 27858 39454 27860 39506
rect 27804 39442 27860 39454
rect 27916 41300 27972 41310
rect 27804 38948 27860 38958
rect 27916 38948 27972 41244
rect 28028 40628 28084 40638
rect 28028 40534 28084 40572
rect 27804 38946 27972 38948
rect 27804 38894 27806 38946
rect 27858 38894 27972 38946
rect 27804 38892 27972 38894
rect 27804 38882 27860 38892
rect 27692 38782 27694 38834
rect 27746 38782 27748 38834
rect 27692 38770 27748 38782
rect 28140 38724 28196 42588
rect 28252 42642 28308 42654
rect 28252 42590 28254 42642
rect 28306 42590 28308 42642
rect 28252 42420 28308 42590
rect 28364 42642 28420 42924
rect 28476 42756 28532 44044
rect 28588 44034 28644 44044
rect 28700 43876 28756 45052
rect 28700 43810 28756 43820
rect 28924 45330 28980 47404
rect 28924 45278 28926 45330
rect 28978 45278 28980 45330
rect 28924 43764 28980 45278
rect 29148 44772 29204 52670
rect 29820 52722 29876 52782
rect 29820 52670 29822 52722
rect 29874 52670 29876 52722
rect 29820 52658 29876 52670
rect 30268 52834 30324 55412
rect 30604 55318 30660 55356
rect 32172 55412 32228 55916
rect 32172 55346 32228 55356
rect 32956 55410 33012 56588
rect 33628 56308 33684 56700
rect 33628 56214 33684 56252
rect 33180 55970 33236 55982
rect 33180 55918 33182 55970
rect 33234 55918 33236 55970
rect 32956 55358 32958 55410
rect 33010 55358 33012 55410
rect 32956 55346 33012 55358
rect 33068 55524 33124 55534
rect 33180 55524 33236 55918
rect 33124 55468 33236 55524
rect 33292 55972 33348 55982
rect 30604 55188 30660 55198
rect 30604 54514 30660 55132
rect 31164 55188 31220 55198
rect 31164 55094 31220 55132
rect 30716 55076 30772 55086
rect 30716 54738 30772 55020
rect 31388 55076 31444 55086
rect 31388 54982 31444 55020
rect 31612 55074 31668 55086
rect 31612 55022 31614 55074
rect 31666 55022 31668 55074
rect 31164 54964 31220 54974
rect 30716 54686 30718 54738
rect 30770 54686 30772 54738
rect 30716 54674 30772 54686
rect 30940 54740 30996 54750
rect 30940 54646 30996 54684
rect 30604 54462 30606 54514
rect 30658 54462 30660 54514
rect 30492 54292 30548 54302
rect 30492 53954 30548 54236
rect 30492 53902 30494 53954
rect 30546 53902 30548 53954
rect 30492 53890 30548 53902
rect 30604 53956 30660 54462
rect 31164 54514 31220 54908
rect 31612 54964 31668 55022
rect 31612 54898 31668 54908
rect 31724 55074 31780 55086
rect 31724 55022 31726 55074
rect 31778 55022 31780 55074
rect 31164 54462 31166 54514
rect 31218 54462 31220 54514
rect 30604 53890 30660 53900
rect 30940 54404 30996 54414
rect 30380 53844 30436 53854
rect 30380 53618 30436 53788
rect 30828 53844 30884 53854
rect 30828 53750 30884 53788
rect 30380 53566 30382 53618
rect 30434 53566 30436 53618
rect 30380 53554 30436 53566
rect 30268 52782 30270 52834
rect 30322 52782 30324 52834
rect 30268 52724 30324 52782
rect 30268 52658 30324 52668
rect 30828 53396 30884 53406
rect 30716 52388 30772 52398
rect 29820 52276 29876 52286
rect 29820 52182 29876 52220
rect 30044 52162 30100 52174
rect 30044 52110 30046 52162
rect 30098 52110 30100 52162
rect 29708 51492 29764 51502
rect 29372 51268 29428 51278
rect 29148 44706 29204 44716
rect 29260 51266 29428 51268
rect 29260 51214 29374 51266
rect 29426 51214 29428 51266
rect 29260 51212 29428 51214
rect 28700 43540 28756 43550
rect 28924 43540 28980 43708
rect 28700 43538 28980 43540
rect 28700 43486 28702 43538
rect 28754 43486 28980 43538
rect 28700 43484 28980 43486
rect 28700 43474 28756 43484
rect 28476 42700 28980 42756
rect 28364 42590 28366 42642
rect 28418 42590 28420 42642
rect 28364 42578 28420 42590
rect 28588 42532 28644 42542
rect 28588 42530 28868 42532
rect 28588 42478 28590 42530
rect 28642 42478 28868 42530
rect 28588 42476 28868 42478
rect 28588 42466 28644 42476
rect 28252 42364 28532 42420
rect 28252 41860 28308 41870
rect 28252 41186 28308 41804
rect 28252 41134 28254 41186
rect 28306 41134 28308 41186
rect 28252 40628 28308 41134
rect 28364 41636 28420 41646
rect 28364 40628 28420 41580
rect 28476 41186 28532 42364
rect 28588 41972 28644 41982
rect 28588 41878 28644 41916
rect 28812 41970 28868 42476
rect 28812 41918 28814 41970
rect 28866 41918 28868 41970
rect 28812 41906 28868 41918
rect 28476 41134 28478 41186
rect 28530 41134 28532 41186
rect 28476 41076 28532 41134
rect 28924 41188 28980 42700
rect 28924 41122 28980 41132
rect 28476 41010 28532 41020
rect 28812 40964 28868 40974
rect 28812 40962 29092 40964
rect 28812 40910 28814 40962
rect 28866 40910 29092 40962
rect 28812 40908 29092 40910
rect 28812 40898 28868 40908
rect 28476 40628 28532 40638
rect 28924 40628 28980 40638
rect 28364 40626 28980 40628
rect 28364 40574 28478 40626
rect 28530 40574 28926 40626
rect 28978 40574 28980 40626
rect 28364 40572 28980 40574
rect 28252 40562 28308 40572
rect 28476 40562 28532 40572
rect 28924 40516 28980 40572
rect 28924 40450 28980 40460
rect 28364 39394 28420 39406
rect 28364 39342 28366 39394
rect 28418 39342 28420 39394
rect 28364 39060 28420 39342
rect 28364 38994 28420 39004
rect 28812 39394 28868 39406
rect 28812 39342 28814 39394
rect 28866 39342 28868 39394
rect 28700 38948 28756 38958
rect 28700 38854 28756 38892
rect 27580 37998 27582 38050
rect 27634 37998 27636 38050
rect 27580 37986 27636 37998
rect 27804 38612 28196 38668
rect 28364 38834 28420 38846
rect 28364 38782 28366 38834
rect 28418 38782 28420 38834
rect 27804 37490 27860 38612
rect 28364 38276 28420 38782
rect 28476 38836 28532 38846
rect 28476 38742 28532 38780
rect 28812 38834 28868 39342
rect 28812 38782 28814 38834
rect 28866 38782 28868 38834
rect 28812 38724 28868 38782
rect 28812 38658 28868 38668
rect 28364 38210 28420 38220
rect 28812 38500 28868 38510
rect 28812 38162 28868 38444
rect 28812 38110 28814 38162
rect 28866 38110 28868 38162
rect 28812 38098 28868 38110
rect 28252 37938 28308 37950
rect 28252 37886 28254 37938
rect 28306 37886 28308 37938
rect 28252 37604 28308 37886
rect 28252 37538 28308 37548
rect 27804 37438 27806 37490
rect 27858 37438 27860 37490
rect 27804 37426 27860 37438
rect 27468 37324 27636 37380
rect 27468 37156 27524 37166
rect 27132 33618 27188 33628
rect 27244 37044 27300 37054
rect 27244 35922 27300 36988
rect 27244 35870 27246 35922
rect 27298 35870 27300 35922
rect 26908 32734 26910 32786
rect 26962 32734 26964 32786
rect 26908 32722 26964 32734
rect 26460 32564 26516 32574
rect 27132 32564 27188 32574
rect 26236 29988 26292 29998
rect 26236 29894 26292 29932
rect 26124 29596 26292 29652
rect 25564 29540 25620 29550
rect 25564 29426 25620 29484
rect 26124 29428 26180 29438
rect 25564 29374 25566 29426
rect 25618 29374 25620 29426
rect 25564 29362 25620 29374
rect 25676 29426 26180 29428
rect 25676 29374 26126 29426
rect 26178 29374 26180 29426
rect 25676 29372 26180 29374
rect 25452 28532 25508 28542
rect 25676 28532 25732 29372
rect 26124 29362 26180 29372
rect 25900 28756 25956 28766
rect 25900 28662 25956 28700
rect 25452 28530 25732 28532
rect 25452 28478 25454 28530
rect 25506 28478 25732 28530
rect 25452 28476 25732 28478
rect 25452 28466 25508 28476
rect 25676 28084 25732 28094
rect 25676 27990 25732 28028
rect 26236 28084 26292 29596
rect 26460 29540 26516 32508
rect 27020 32562 27188 32564
rect 27020 32510 27134 32562
rect 27186 32510 27188 32562
rect 27020 32508 27188 32510
rect 27020 31948 27076 32508
rect 27132 32498 27188 32508
rect 26796 31892 27076 31948
rect 27244 31892 27300 35870
rect 27356 36594 27412 36606
rect 27356 36542 27358 36594
rect 27410 36542 27412 36594
rect 27356 35922 27412 36542
rect 27356 35870 27358 35922
rect 27410 35870 27412 35922
rect 27356 35858 27412 35870
rect 27468 35810 27524 37100
rect 27468 35758 27470 35810
rect 27522 35758 27524 35810
rect 27468 35746 27524 35758
rect 27356 31892 27412 31902
rect 26572 31556 26628 31566
rect 26796 31556 26852 31892
rect 27132 31890 27524 31892
rect 27132 31838 27358 31890
rect 27410 31838 27524 31890
rect 27132 31836 27524 31838
rect 26572 31554 26852 31556
rect 26572 31502 26574 31554
rect 26626 31502 26852 31554
rect 26572 31500 26852 31502
rect 27020 31668 27076 31678
rect 26572 29988 26628 31500
rect 27020 30210 27076 31612
rect 27132 31218 27188 31836
rect 27356 31826 27412 31836
rect 27468 31332 27524 31836
rect 27580 31556 27636 37324
rect 28140 37268 28196 37278
rect 27916 37044 27972 37054
rect 27692 36708 27748 36718
rect 27692 36614 27748 36652
rect 27916 35922 27972 36988
rect 28140 36260 28196 37212
rect 28476 37156 28532 37166
rect 28476 36706 28532 37100
rect 28476 36654 28478 36706
rect 28530 36654 28532 36706
rect 28476 36642 28532 36654
rect 28700 36820 28756 36830
rect 28700 36370 28756 36764
rect 28812 36594 28868 36606
rect 28812 36542 28814 36594
rect 28866 36542 28868 36594
rect 28812 36484 28868 36542
rect 28812 36418 28868 36428
rect 28700 36318 28702 36370
rect 28754 36318 28756 36370
rect 28700 36306 28756 36318
rect 29036 36372 29092 40908
rect 29148 37156 29204 37166
rect 29148 37062 29204 37100
rect 29260 36932 29316 51212
rect 29372 51202 29428 51212
rect 29372 50372 29428 50382
rect 29372 50034 29428 50316
rect 29372 49982 29374 50034
rect 29426 49982 29428 50034
rect 29372 49970 29428 49982
rect 29372 49028 29428 49038
rect 29372 44100 29428 48972
rect 29708 48916 29764 51436
rect 30044 51378 30100 52110
rect 30716 52050 30772 52332
rect 30716 51998 30718 52050
rect 30770 51998 30772 52050
rect 30716 51986 30772 51998
rect 30380 51492 30436 51502
rect 30380 51398 30436 51436
rect 30044 51326 30046 51378
rect 30098 51326 30100 51378
rect 29820 51268 29876 51278
rect 29820 50594 29876 51212
rect 29932 50708 29988 50718
rect 29932 50614 29988 50652
rect 29820 50542 29822 50594
rect 29874 50542 29876 50594
rect 29820 50530 29876 50542
rect 29820 49700 29876 49710
rect 29820 49698 29988 49700
rect 29820 49646 29822 49698
rect 29874 49646 29988 49698
rect 29820 49644 29988 49646
rect 29820 49634 29876 49644
rect 29820 48916 29876 48926
rect 29708 48914 29876 48916
rect 29708 48862 29822 48914
rect 29874 48862 29876 48914
rect 29708 48860 29876 48862
rect 29820 48850 29876 48860
rect 29932 48468 29988 49644
rect 29932 48402 29988 48412
rect 29708 48242 29764 48254
rect 29708 48190 29710 48242
rect 29762 48190 29764 48242
rect 29484 48020 29540 48030
rect 29708 48020 29764 48190
rect 29932 48244 29988 48254
rect 29932 48150 29988 48188
rect 29484 48018 29764 48020
rect 29484 47966 29486 48018
rect 29538 47966 29764 48018
rect 29484 47964 29764 47966
rect 29484 47954 29540 47964
rect 29484 47236 29540 47246
rect 29484 46674 29540 47180
rect 29484 46622 29486 46674
rect 29538 46622 29540 46674
rect 29484 46610 29540 46622
rect 29708 46450 29764 47964
rect 29820 48130 29876 48142
rect 29820 48078 29822 48130
rect 29874 48078 29876 48130
rect 29820 47572 29876 48078
rect 30044 48020 30100 51326
rect 30156 51268 30212 51278
rect 30156 50148 30212 51212
rect 30828 50596 30884 53340
rect 30940 52946 30996 54348
rect 31164 53844 31220 54462
rect 31612 54740 31668 54750
rect 31612 54516 31668 54684
rect 31724 54628 31780 55022
rect 32172 55074 32228 55086
rect 32172 55022 32174 55074
rect 32226 55022 32228 55074
rect 32172 54964 32228 55022
rect 32172 54898 32228 54908
rect 32620 55074 32676 55086
rect 32620 55022 32622 55074
rect 32674 55022 32676 55074
rect 32620 54964 32676 55022
rect 32620 54898 32676 54908
rect 33068 54740 33124 55468
rect 32284 54684 33124 54740
rect 31724 54572 32116 54628
rect 31612 54460 31892 54516
rect 31276 54404 31332 54414
rect 31276 54310 31332 54348
rect 31836 54402 31892 54460
rect 31836 54350 31838 54402
rect 31890 54350 31892 54402
rect 31164 53170 31220 53788
rect 31836 53730 31892 54350
rect 31836 53678 31838 53730
rect 31890 53678 31892 53730
rect 31836 53666 31892 53678
rect 31948 54402 32004 54414
rect 31948 54350 31950 54402
rect 32002 54350 32004 54402
rect 31948 53732 32004 54350
rect 32060 53842 32116 54572
rect 32060 53790 32062 53842
rect 32114 53790 32116 53842
rect 32060 53778 32116 53790
rect 31164 53118 31166 53170
rect 31218 53118 31220 53170
rect 31164 53106 31220 53118
rect 31948 53172 32004 53676
rect 31948 53106 32004 53116
rect 30940 52894 30942 52946
rect 30994 52894 30996 52946
rect 30940 52836 30996 52894
rect 31612 52836 31668 52846
rect 30940 52834 31668 52836
rect 30940 52782 31614 52834
rect 31666 52782 31668 52834
rect 30940 52780 31668 52782
rect 31276 52052 31332 52062
rect 31276 51938 31332 51996
rect 31276 51886 31278 51938
rect 31330 51886 31332 51938
rect 31276 51716 31332 51886
rect 31276 51650 31332 51660
rect 31052 51604 31108 51614
rect 31052 51510 31108 51548
rect 31612 51604 31668 52780
rect 32060 52836 32116 52846
rect 32060 52834 32228 52836
rect 32060 52782 32062 52834
rect 32114 52782 32228 52834
rect 32060 52780 32228 52782
rect 32060 52770 32116 52780
rect 32060 52276 32116 52286
rect 31836 52052 31892 52062
rect 31836 51958 31892 51996
rect 32060 52050 32116 52220
rect 32060 51998 32062 52050
rect 32114 51998 32116 52050
rect 32060 51986 32116 51998
rect 31612 51538 31668 51548
rect 31948 51938 32004 51950
rect 31948 51886 31950 51938
rect 32002 51886 32004 51938
rect 31724 51490 31780 51502
rect 31724 51438 31726 51490
rect 31778 51438 31780 51490
rect 31612 51380 31668 51390
rect 31612 51286 31668 51324
rect 31388 51156 31444 51166
rect 30828 50540 30996 50596
rect 30156 50082 30212 50092
rect 30604 50484 30660 50494
rect 30268 49698 30324 49710
rect 30268 49646 30270 49698
rect 30322 49646 30324 49698
rect 30268 49586 30324 49646
rect 30604 49700 30660 50428
rect 30716 50484 30772 50494
rect 30716 50482 30884 50484
rect 30716 50430 30718 50482
rect 30770 50430 30884 50482
rect 30716 50428 30884 50430
rect 30716 50418 30772 50428
rect 30828 49924 30884 50428
rect 30828 49858 30884 49868
rect 30716 49700 30772 49710
rect 30604 49698 30884 49700
rect 30604 49646 30718 49698
rect 30770 49646 30884 49698
rect 30604 49644 30884 49646
rect 30716 49634 30772 49644
rect 30268 49534 30270 49586
rect 30322 49534 30324 49586
rect 30268 49522 30324 49534
rect 29820 47506 29876 47516
rect 29932 47964 30100 48020
rect 30156 49026 30212 49038
rect 30156 48974 30158 49026
rect 30210 48974 30212 49026
rect 29932 46786 29988 47964
rect 30156 47684 30212 48974
rect 30604 49028 30660 49038
rect 30604 48934 30660 48972
rect 30380 48242 30436 48254
rect 30380 48190 30382 48242
rect 30434 48190 30436 48242
rect 30380 48132 30436 48190
rect 30716 48132 30772 48142
rect 30380 48130 30772 48132
rect 30380 48078 30718 48130
rect 30770 48078 30772 48130
rect 30380 48076 30772 48078
rect 30156 47618 30212 47628
rect 30268 47572 30324 47582
rect 30268 47478 30324 47516
rect 30156 47458 30212 47470
rect 30156 47406 30158 47458
rect 30210 47406 30212 47458
rect 30156 47236 30212 47406
rect 30156 47170 30212 47180
rect 30716 46900 30772 48076
rect 29932 46734 29934 46786
rect 29986 46734 29988 46786
rect 29932 46722 29988 46734
rect 30268 46898 30772 46900
rect 30268 46846 30718 46898
rect 30770 46846 30772 46898
rect 30268 46844 30772 46846
rect 30268 46786 30324 46844
rect 30268 46734 30270 46786
rect 30322 46734 30324 46786
rect 30268 46722 30324 46734
rect 29708 46398 29710 46450
rect 29762 46398 29764 46450
rect 29484 46228 29540 46238
rect 29708 46228 29764 46398
rect 29540 46172 29764 46228
rect 30044 46674 30100 46686
rect 30044 46622 30046 46674
rect 30098 46622 30100 46674
rect 29484 46002 29540 46172
rect 29484 45950 29486 46002
rect 29538 45950 29540 46002
rect 29484 45938 29540 45950
rect 29484 45556 29540 45566
rect 29484 44212 29540 45500
rect 29596 45106 29652 46172
rect 30044 45556 30100 46622
rect 30268 46114 30324 46126
rect 30268 46062 30270 46114
rect 30322 46062 30324 46114
rect 30268 46002 30324 46062
rect 30268 45950 30270 46002
rect 30322 45950 30324 46002
rect 30268 45938 30324 45950
rect 30044 45490 30100 45500
rect 29596 45054 29598 45106
rect 29650 45054 29652 45106
rect 29596 45042 29652 45054
rect 29932 45106 29988 45118
rect 29932 45054 29934 45106
rect 29986 45054 29988 45106
rect 29932 44322 29988 45054
rect 29932 44270 29934 44322
rect 29986 44270 29988 44322
rect 29932 44258 29988 44270
rect 29596 44212 29652 44222
rect 29484 44210 29652 44212
rect 29484 44158 29598 44210
rect 29650 44158 29652 44210
rect 29484 44156 29652 44158
rect 29372 44034 29428 44044
rect 29372 43764 29428 43774
rect 29372 43650 29428 43708
rect 29372 43598 29374 43650
rect 29426 43598 29428 43650
rect 29372 43586 29428 43598
rect 29484 42980 29540 42990
rect 29484 42866 29540 42924
rect 29484 42814 29486 42866
rect 29538 42814 29540 42866
rect 29484 42802 29540 42814
rect 29596 42420 29652 44156
rect 29708 44100 29764 44138
rect 30268 44100 30324 44110
rect 29708 44034 29764 44044
rect 30156 44098 30324 44100
rect 30156 44046 30270 44098
rect 30322 44046 30324 44098
rect 30156 44044 30324 44046
rect 29708 43876 29764 43886
rect 29708 43762 29764 43820
rect 30156 43764 30212 44044
rect 30268 44034 30324 44044
rect 29708 43710 29710 43762
rect 29762 43710 29764 43762
rect 29708 43698 29764 43710
rect 30044 43708 30156 43764
rect 29932 42980 29988 42990
rect 29932 42866 29988 42924
rect 29932 42814 29934 42866
rect 29986 42814 29988 42866
rect 29932 42802 29988 42814
rect 29596 42354 29652 42364
rect 29484 42196 29540 42206
rect 29484 42082 29540 42140
rect 30044 42194 30100 43708
rect 30156 43698 30212 43708
rect 30044 42142 30046 42194
rect 30098 42142 30100 42194
rect 30044 42130 30100 42142
rect 30156 43426 30212 43438
rect 30156 43374 30158 43426
rect 30210 43374 30212 43426
rect 30156 42644 30212 43374
rect 29484 42030 29486 42082
rect 29538 42030 29540 42082
rect 29484 42018 29540 42030
rect 29820 42084 29876 42094
rect 29820 41188 29876 42028
rect 29484 41186 29876 41188
rect 29484 41134 29822 41186
rect 29874 41134 29876 41186
rect 29484 41132 29876 41134
rect 29372 40964 29428 40974
rect 29372 40516 29428 40908
rect 29484 40516 29540 41132
rect 29820 41122 29876 41132
rect 29596 40964 29652 40974
rect 29596 40870 29652 40908
rect 29708 40962 29764 40974
rect 29708 40910 29710 40962
rect 29762 40910 29764 40962
rect 29708 40628 29764 40910
rect 30044 40964 30100 40974
rect 30044 40870 30100 40908
rect 29708 40572 29876 40628
rect 29484 40460 29652 40516
rect 29372 40422 29428 40460
rect 29596 40402 29652 40460
rect 29596 40350 29598 40402
rect 29650 40350 29652 40402
rect 29596 40338 29652 40350
rect 29820 40402 29876 40572
rect 29820 40350 29822 40402
rect 29874 40350 29876 40402
rect 29820 40338 29876 40350
rect 29484 40290 29540 40302
rect 29484 40238 29486 40290
rect 29538 40238 29540 40290
rect 29484 38164 29540 40238
rect 29932 39396 29988 39406
rect 29820 39394 29988 39396
rect 29820 39342 29934 39394
rect 29986 39342 29988 39394
rect 29820 39340 29988 39342
rect 29484 38098 29540 38108
rect 29596 38722 29652 38734
rect 29596 38670 29598 38722
rect 29650 38670 29652 38722
rect 29596 38052 29652 38670
rect 29820 38500 29876 39340
rect 29932 39330 29988 39340
rect 30044 39060 30100 39070
rect 30044 38668 30100 39004
rect 29820 38434 29876 38444
rect 29932 38612 30100 38668
rect 29596 37958 29652 37996
rect 29932 37492 29988 38612
rect 30044 38052 30100 38062
rect 30044 37958 30100 37996
rect 29932 37426 29988 37436
rect 28140 36194 28196 36204
rect 28812 36260 28868 36270
rect 27916 35870 27918 35922
rect 27970 35870 27972 35922
rect 27692 35476 27748 35486
rect 27692 31668 27748 35420
rect 27916 35028 27972 35870
rect 28588 35588 28644 35626
rect 28588 35522 28644 35532
rect 28812 35308 28868 36204
rect 29036 35698 29092 36316
rect 29036 35646 29038 35698
rect 29090 35646 29092 35698
rect 29036 35634 29092 35646
rect 29148 36876 29316 36932
rect 29596 37266 29652 37278
rect 29596 37214 29598 37266
rect 29650 37214 29652 37266
rect 28588 35252 28644 35262
rect 28588 35138 28644 35196
rect 28588 35086 28590 35138
rect 28642 35086 28644 35138
rect 28588 35074 28644 35086
rect 28700 35252 28868 35308
rect 28924 35588 28980 35598
rect 28924 35308 28980 35532
rect 28924 35252 29092 35308
rect 27916 35026 28532 35028
rect 27916 34974 27918 35026
rect 27970 34974 28532 35026
rect 27916 34972 28532 34974
rect 27916 34962 27972 34972
rect 28476 34914 28532 34972
rect 28476 34862 28478 34914
rect 28530 34862 28532 34914
rect 28476 34850 28532 34862
rect 28252 34356 28308 34366
rect 28700 34356 28756 35252
rect 28140 34300 28252 34356
rect 27804 34132 27860 34142
rect 27804 34038 27860 34076
rect 27804 33124 27860 33134
rect 27804 32676 27860 33068
rect 27804 32582 27860 32620
rect 28140 31892 28196 34300
rect 28252 34262 28308 34300
rect 28588 34300 28756 34356
rect 28364 34132 28420 34142
rect 28252 33122 28308 33134
rect 28252 33070 28254 33122
rect 28306 33070 28308 33122
rect 28252 32340 28308 33070
rect 28252 32274 28308 32284
rect 28364 31892 28420 34076
rect 28476 32564 28532 32574
rect 28476 32470 28532 32508
rect 28140 31826 28196 31836
rect 28252 31836 28420 31892
rect 28588 31892 28644 34300
rect 28700 34020 28756 34030
rect 28700 33926 28756 33964
rect 28924 33684 28980 33694
rect 28924 33570 28980 33628
rect 28924 33518 28926 33570
rect 28978 33518 28980 33570
rect 28924 33506 28980 33518
rect 28924 32450 28980 32462
rect 28924 32398 28926 32450
rect 28978 32398 28980 32450
rect 28924 32340 28980 32398
rect 28924 32274 28980 32284
rect 27692 31602 27748 31612
rect 27580 31490 27636 31500
rect 27468 31276 28196 31332
rect 27132 31166 27134 31218
rect 27186 31166 27188 31218
rect 27132 31154 27188 31166
rect 27580 30996 27636 31006
rect 27020 30158 27022 30210
rect 27074 30158 27076 30210
rect 27020 30146 27076 30158
rect 27468 30994 27636 30996
rect 27468 30942 27582 30994
rect 27634 30942 27636 30994
rect 27468 30940 27636 30942
rect 27468 30884 27524 30940
rect 27580 30930 27636 30940
rect 28140 30994 28196 31276
rect 28140 30942 28142 30994
rect 28194 30942 28196 30994
rect 28140 30930 28196 30942
rect 26572 29922 26628 29932
rect 27356 29988 27412 29998
rect 27244 29876 27300 29886
rect 27132 29652 27188 29662
rect 27244 29652 27300 29820
rect 27188 29596 27300 29652
rect 27132 29586 27188 29596
rect 26460 29474 26516 29484
rect 26460 28980 26516 28990
rect 26460 28754 26516 28924
rect 26460 28702 26462 28754
rect 26514 28702 26516 28754
rect 26460 28690 26516 28702
rect 27020 28980 27076 28990
rect 27020 28530 27076 28924
rect 27020 28478 27022 28530
rect 27074 28478 27076 28530
rect 26684 28084 26740 28094
rect 26236 28082 26740 28084
rect 26236 28030 26686 28082
rect 26738 28030 26740 28082
rect 26236 28028 26740 28030
rect 26236 27858 26292 28028
rect 26684 28018 26740 28028
rect 26236 27806 26238 27858
rect 26290 27806 26292 27858
rect 26012 27636 26068 27646
rect 26012 27542 26068 27580
rect 26124 27188 26180 27198
rect 26236 27188 26292 27806
rect 25676 27186 26292 27188
rect 25676 27134 26126 27186
rect 26178 27134 26292 27186
rect 25676 27132 26292 27134
rect 25676 27074 25732 27132
rect 26124 27122 26180 27132
rect 25676 27022 25678 27074
rect 25730 27022 25732 27074
rect 25676 27010 25732 27022
rect 26684 27076 26740 27086
rect 26684 26982 26740 27020
rect 26348 26964 26404 26974
rect 25228 24098 25284 24108
rect 25340 26850 25396 26862
rect 25340 26798 25342 26850
rect 25394 26798 25396 26850
rect 25340 23492 25396 26798
rect 25564 26850 25620 26862
rect 25564 26798 25566 26850
rect 25618 26798 25620 26850
rect 25564 26628 25620 26798
rect 25564 26562 25620 26572
rect 25676 26852 25732 26862
rect 25676 26514 25732 26796
rect 25676 26462 25678 26514
rect 25730 26462 25732 26514
rect 25676 26450 25732 26462
rect 26348 26514 26404 26908
rect 26348 26462 26350 26514
rect 26402 26462 26404 26514
rect 26348 26450 26404 26462
rect 26124 26066 26180 26078
rect 26124 26014 26126 26066
rect 26178 26014 26180 26066
rect 26012 25618 26068 25630
rect 26012 25566 26014 25618
rect 26066 25566 26068 25618
rect 25900 24948 25956 24958
rect 25900 24854 25956 24892
rect 25676 24724 25732 24734
rect 24892 23214 24894 23266
rect 24946 23214 24948 23266
rect 24892 23202 24948 23214
rect 25116 23436 25340 23492
rect 24780 22484 24836 22494
rect 24668 22482 24836 22484
rect 24668 22430 24782 22482
rect 24834 22430 24836 22482
rect 24668 22428 24836 22430
rect 23772 22390 23828 22428
rect 24780 22418 24836 22428
rect 25116 22484 25172 23436
rect 25340 23426 25396 23436
rect 25452 24668 25676 24724
rect 25116 22352 25172 22428
rect 23212 22206 23214 22258
rect 23266 22206 23268 22258
rect 23212 22194 23268 22206
rect 23324 22260 23380 22270
rect 23324 22258 23492 22260
rect 23324 22206 23326 22258
rect 23378 22206 23492 22258
rect 23324 22204 23492 22206
rect 23324 22194 23380 22204
rect 23100 21980 23268 22036
rect 22988 21522 23044 21532
rect 23100 21700 23156 21710
rect 23100 20242 23156 21644
rect 23212 21476 23268 21980
rect 23436 21812 23492 22204
rect 23548 21812 23604 21822
rect 23436 21810 23604 21812
rect 23436 21758 23550 21810
rect 23602 21758 23604 21810
rect 23436 21756 23604 21758
rect 23324 21700 23380 21710
rect 23324 21606 23380 21644
rect 23436 21476 23492 21486
rect 23212 21420 23380 21476
rect 23100 20190 23102 20242
rect 23154 20190 23156 20242
rect 23100 20178 23156 20190
rect 23212 18564 23268 18574
rect 22764 18508 22932 18564
rect 22652 17892 22708 18396
rect 22764 18340 22820 18350
rect 22764 18246 22820 18284
rect 22876 17892 22932 18508
rect 23212 18470 23268 18508
rect 22652 17836 22820 17892
rect 22652 17668 22708 17678
rect 22652 17574 22708 17612
rect 22764 16884 22820 17836
rect 22876 17826 22932 17836
rect 23212 17780 23268 17790
rect 23212 17666 23268 17724
rect 23212 17614 23214 17666
rect 23266 17614 23268 17666
rect 22988 17108 23044 17118
rect 22988 17014 23044 17052
rect 23212 16996 23268 17614
rect 23212 16930 23268 16940
rect 22988 16884 23044 16894
rect 22764 16828 22988 16884
rect 22988 16790 23044 16828
rect 23212 16212 23268 16222
rect 23212 16118 23268 16156
rect 22652 15314 22708 15326
rect 22652 15262 22654 15314
rect 22706 15262 22708 15314
rect 22316 13972 22372 14476
rect 22316 13746 22372 13916
rect 22540 15202 22596 15214
rect 22540 15150 22542 15202
rect 22594 15150 22596 15202
rect 22540 14642 22596 15150
rect 22540 14590 22542 14642
rect 22594 14590 22596 14642
rect 22540 13858 22596 14590
rect 22652 14532 22708 15262
rect 22652 14438 22708 14476
rect 22988 13972 23044 13982
rect 22988 13878 23044 13916
rect 22540 13806 22542 13858
rect 22594 13806 22596 13858
rect 22540 13794 22596 13806
rect 22316 13694 22318 13746
rect 22370 13694 22372 13746
rect 22316 13682 22372 13694
rect 22652 12178 22708 12190
rect 22652 12126 22654 12178
rect 22706 12126 22708 12178
rect 22652 10836 22708 12126
rect 22876 12066 22932 12078
rect 22876 12014 22878 12066
rect 22930 12014 22932 12066
rect 22876 11618 22932 12014
rect 23212 11844 23268 11854
rect 23212 11620 23268 11788
rect 22876 11566 22878 11618
rect 22930 11566 22932 11618
rect 22876 11396 22932 11566
rect 22876 11330 22932 11340
rect 22988 11564 23268 11620
rect 22652 10770 22708 10780
rect 22540 10610 22596 10622
rect 22540 10558 22542 10610
rect 22594 10558 22596 10610
rect 22540 9828 22596 10558
rect 22540 9762 22596 9772
rect 22876 10498 22932 10510
rect 22876 10446 22878 10498
rect 22930 10446 22932 10498
rect 22876 9492 22932 10446
rect 22988 10386 23044 11564
rect 23212 11506 23268 11564
rect 23212 11454 23214 11506
rect 23266 11454 23268 11506
rect 23212 11442 23268 11454
rect 22988 10334 22990 10386
rect 23042 10334 23044 10386
rect 22988 10322 23044 10334
rect 23100 11394 23156 11406
rect 23100 11342 23102 11394
rect 23154 11342 23156 11394
rect 23100 9938 23156 11342
rect 23100 9886 23102 9938
rect 23154 9886 23156 9938
rect 23100 9874 23156 9886
rect 22988 9828 23044 9838
rect 22988 9714 23044 9772
rect 22988 9662 22990 9714
rect 23042 9662 23044 9714
rect 22988 9650 23044 9662
rect 23212 9714 23268 9726
rect 23212 9662 23214 9714
rect 23266 9662 23268 9714
rect 22876 9426 22932 9436
rect 23212 9492 23268 9662
rect 23212 9426 23268 9436
rect 21980 9266 22148 9268
rect 21980 9214 21982 9266
rect 22034 9214 22148 9266
rect 21980 9212 22148 9214
rect 21980 8482 22036 9212
rect 21980 8430 21982 8482
rect 22034 8430 22036 8482
rect 21980 8372 22036 8430
rect 21980 8306 22036 8316
rect 22540 8932 22596 8942
rect 22988 8932 23044 8942
rect 22540 8930 23044 8932
rect 22540 8878 22542 8930
rect 22594 8878 22990 8930
rect 23042 8878 23044 8930
rect 22540 8876 23044 8878
rect 22204 8260 22260 8270
rect 22204 8148 22260 8204
rect 22540 8148 22596 8876
rect 22988 8866 23044 8876
rect 22764 8372 22820 8382
rect 22764 8278 22820 8316
rect 22204 8146 22596 8148
rect 22204 8094 22206 8146
rect 22258 8094 22596 8146
rect 22204 8092 22596 8094
rect 22204 8082 22260 8092
rect 22540 7924 22596 8092
rect 22540 7858 22596 7868
rect 23212 8034 23268 8046
rect 23212 7982 23214 8034
rect 23266 7982 23268 8034
rect 22092 7476 22148 7486
rect 22092 7382 22148 7420
rect 23212 7476 23268 7982
rect 23212 7410 23268 7420
rect 22316 7362 22372 7374
rect 22316 7310 22318 7362
rect 22370 7310 22372 7362
rect 22316 7140 22372 7310
rect 22988 7364 23044 7374
rect 22988 7362 23156 7364
rect 22988 7310 22990 7362
rect 23042 7310 23156 7362
rect 22988 7308 23156 7310
rect 22988 7298 23044 7308
rect 22316 7074 22372 7084
rect 22876 7140 22932 7150
rect 21644 6802 21812 6804
rect 21644 6750 21646 6802
rect 21698 6750 21812 6802
rect 21644 6748 21812 6750
rect 21644 6738 21700 6748
rect 22876 6690 22932 7084
rect 22876 6638 22878 6690
rect 22930 6638 22932 6690
rect 22876 6626 22932 6638
rect 21420 6066 21476 6076
rect 22988 6466 23044 6478
rect 22988 6414 22990 6466
rect 23042 6414 23044 6466
rect 20412 5966 20414 6018
rect 20466 5966 20468 6018
rect 20412 5954 20468 5966
rect 22092 5908 22148 5918
rect 22988 5908 23044 6414
rect 21980 5906 23044 5908
rect 21980 5854 22094 5906
rect 22146 5854 23044 5906
rect 21980 5852 23044 5854
rect 20748 5682 20804 5694
rect 20748 5630 20750 5682
rect 20802 5630 20804 5682
rect 20748 5236 20804 5630
rect 21644 5236 21700 5246
rect 20748 5234 21700 5236
rect 20748 5182 21646 5234
rect 21698 5182 21700 5234
rect 20748 5180 21700 5182
rect 20524 5124 20580 5134
rect 20524 5030 20580 5068
rect 20636 5122 20692 5134
rect 20636 5070 20638 5122
rect 20690 5070 20692 5122
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20636 4340 20692 5070
rect 20748 5010 20804 5180
rect 21644 5170 21700 5180
rect 21868 5124 21924 5134
rect 21868 5030 21924 5068
rect 20748 4958 20750 5010
rect 20802 4958 20804 5010
rect 20748 4946 20804 4958
rect 20636 4274 20692 4284
rect 21980 4788 22036 5852
rect 22092 5842 22148 5852
rect 22092 5682 22148 5694
rect 22092 5630 22094 5682
rect 22146 5630 22148 5682
rect 22092 5346 22148 5630
rect 22092 5294 22094 5346
rect 22146 5294 22148 5346
rect 22092 5282 22148 5294
rect 22428 5682 22484 5694
rect 22428 5630 22430 5682
rect 22482 5630 22484 5682
rect 21980 4338 22036 4732
rect 21980 4286 21982 4338
rect 22034 4286 22036 4338
rect 21980 4274 22036 4286
rect 22428 5012 22484 5630
rect 22428 4338 22484 4956
rect 23100 5012 23156 7308
rect 23212 7252 23268 7262
rect 23212 6690 23268 7196
rect 23212 6638 23214 6690
rect 23266 6638 23268 6690
rect 23212 6626 23268 6638
rect 23324 5572 23380 21420
rect 23436 21382 23492 21420
rect 23548 20804 23604 21756
rect 24780 21700 24836 21710
rect 24780 21606 24836 21644
rect 23996 21586 24052 21598
rect 23996 21534 23998 21586
rect 24050 21534 24052 21586
rect 23996 21476 24052 21534
rect 24332 21476 24388 21486
rect 23996 21474 24388 21476
rect 23996 21422 24334 21474
rect 24386 21422 24388 21474
rect 23996 21420 24388 21422
rect 24332 21362 24388 21420
rect 24332 21310 24334 21362
rect 24386 21310 24388 21362
rect 24332 21298 24388 21310
rect 24668 21362 24724 21374
rect 24668 21310 24670 21362
rect 24722 21310 24724 21362
rect 23772 20804 23828 20814
rect 23548 20802 23828 20804
rect 23548 20750 23774 20802
rect 23826 20750 23828 20802
rect 23548 20748 23828 20750
rect 23772 20738 23828 20748
rect 24108 20690 24164 20702
rect 24108 20638 24110 20690
rect 24162 20638 24164 20690
rect 23436 20580 23492 20590
rect 23436 20486 23492 20524
rect 23996 20580 24052 20590
rect 23996 20486 24052 20524
rect 24108 20468 24164 20638
rect 24668 20690 24724 21310
rect 25116 21364 25172 21374
rect 25452 21364 25508 24668
rect 25676 24630 25732 24668
rect 25788 24612 25844 24622
rect 25788 24518 25844 24556
rect 26012 24388 26068 25566
rect 26012 23828 26068 24332
rect 26124 24052 26180 26014
rect 26908 26066 26964 26078
rect 26908 26014 26910 26066
rect 26962 26014 26964 26066
rect 26460 25282 26516 25294
rect 26460 25230 26462 25282
rect 26514 25230 26516 25282
rect 26460 24948 26516 25230
rect 26908 25172 26964 26014
rect 27020 25620 27076 28478
rect 27244 28532 27300 29596
rect 27356 29652 27412 29932
rect 27356 29586 27412 29596
rect 27356 28532 27412 28542
rect 27244 28530 27412 28532
rect 27244 28478 27358 28530
rect 27410 28478 27412 28530
rect 27244 28476 27412 28478
rect 27356 28466 27412 28476
rect 27468 27076 27524 30828
rect 27916 29428 27972 29438
rect 27692 27860 27748 27870
rect 27244 26964 27300 27002
rect 27468 26982 27524 27020
rect 27580 27188 27636 27198
rect 27244 26898 27300 26908
rect 27580 25732 27636 27132
rect 27692 26514 27748 27804
rect 27916 26908 27972 29372
rect 28140 27972 28196 27982
rect 28140 27878 28196 27916
rect 28140 27188 28196 27198
rect 28252 27188 28308 31836
rect 28588 31666 28644 31836
rect 28588 31614 28590 31666
rect 28642 31614 28644 31666
rect 28588 31602 28644 31614
rect 28140 27186 28252 27188
rect 28140 27134 28142 27186
rect 28194 27134 28252 27186
rect 28140 27132 28252 27134
rect 28140 27122 28196 27132
rect 28028 27076 28084 27114
rect 28252 27056 28308 27132
rect 28364 31556 28420 31566
rect 28028 27010 28084 27020
rect 27916 26852 28308 26908
rect 27692 26462 27694 26514
rect 27746 26462 27748 26514
rect 27692 26450 27748 26462
rect 28140 25732 28196 25742
rect 28252 25732 28308 26852
rect 28364 25956 28420 31500
rect 29036 31332 29092 35252
rect 29148 32116 29204 36876
rect 29596 36820 29652 37214
rect 29596 36754 29652 36764
rect 30044 37154 30100 37166
rect 30044 37102 30046 37154
rect 30098 37102 30100 37154
rect 30044 36596 30100 37102
rect 29596 36540 30100 36596
rect 29596 36484 29652 36540
rect 29484 36482 29652 36484
rect 29484 36430 29598 36482
rect 29650 36430 29652 36482
rect 29484 36428 29652 36430
rect 29484 35698 29540 36428
rect 29596 36418 29652 36428
rect 29708 36372 29764 36382
rect 29708 36278 29764 36316
rect 29484 35646 29486 35698
rect 29538 35646 29540 35698
rect 29484 35634 29540 35646
rect 29596 36260 29652 36270
rect 29596 34802 29652 36204
rect 30044 35588 30100 35598
rect 29932 35532 30044 35588
rect 29932 35364 29988 35532
rect 30044 35494 30100 35532
rect 29932 34914 29988 35308
rect 29932 34862 29934 34914
rect 29986 34862 29988 34914
rect 29932 34850 29988 34862
rect 29596 34750 29598 34802
rect 29650 34750 29652 34802
rect 29260 34356 29316 34366
rect 29596 34356 29652 34750
rect 29708 34356 29764 34366
rect 29260 34354 29764 34356
rect 29260 34302 29262 34354
rect 29314 34302 29710 34354
rect 29762 34302 29764 34354
rect 29260 34300 29764 34302
rect 29260 34290 29316 34300
rect 29708 34290 29764 34300
rect 29932 34132 29988 34142
rect 29932 34038 29988 34076
rect 29372 34020 29428 34030
rect 29372 33684 29428 33964
rect 29372 33124 29428 33628
rect 29820 34018 29876 34030
rect 29820 33966 29822 34018
rect 29874 33966 29876 34018
rect 29708 33348 29764 33358
rect 29820 33348 29876 33966
rect 30156 33572 30212 42588
rect 30380 42196 30436 46844
rect 30716 46834 30772 46844
rect 30716 46114 30772 46126
rect 30716 46062 30718 46114
rect 30770 46062 30772 46114
rect 30716 45666 30772 46062
rect 30716 45614 30718 45666
rect 30770 45614 30772 45666
rect 30492 44994 30548 45006
rect 30492 44942 30494 44994
rect 30546 44942 30548 44994
rect 30492 44324 30548 44942
rect 30716 44546 30772 45614
rect 30716 44494 30718 44546
rect 30770 44494 30772 44546
rect 30716 44482 30772 44494
rect 30492 44258 30548 44268
rect 30716 44100 30772 44110
rect 30716 44006 30772 44044
rect 30604 43428 30660 43438
rect 30492 43372 30604 43428
rect 30492 42644 30548 43372
rect 30604 43296 30660 43372
rect 30492 42550 30548 42588
rect 30716 42980 30772 42990
rect 30716 42642 30772 42924
rect 30716 42590 30718 42642
rect 30770 42590 30772 42642
rect 30716 42578 30772 42590
rect 30268 42140 30436 42196
rect 30604 42530 30660 42542
rect 30604 42478 30606 42530
rect 30658 42478 30660 42530
rect 30268 35588 30324 42140
rect 30604 42084 30660 42478
rect 30604 42018 30660 42028
rect 30380 41970 30436 41982
rect 30380 41918 30382 41970
rect 30434 41918 30436 41970
rect 30380 40964 30436 41918
rect 30380 40898 30436 40908
rect 30604 40964 30660 40974
rect 30604 40870 30660 40908
rect 30828 40740 30884 49644
rect 30940 49028 30996 50540
rect 31164 50482 31220 50494
rect 31164 50430 31166 50482
rect 31218 50430 31220 50482
rect 31164 50372 31220 50430
rect 30940 48962 30996 48972
rect 31052 49586 31108 49598
rect 31052 49534 31054 49586
rect 31106 49534 31108 49586
rect 30940 48802 30996 48814
rect 30940 48750 30942 48802
rect 30994 48750 30996 48802
rect 30940 48468 30996 48750
rect 30940 48402 30996 48412
rect 30940 48020 30996 48030
rect 30940 47682 30996 47964
rect 30940 47630 30942 47682
rect 30994 47630 30996 47682
rect 30940 47618 30996 47630
rect 31052 45892 31108 49534
rect 31164 49252 31220 50316
rect 31276 50148 31332 50158
rect 31276 50034 31332 50092
rect 31276 49982 31278 50034
rect 31330 49982 31332 50034
rect 31276 49970 31332 49982
rect 31164 49186 31220 49196
rect 30604 40684 30884 40740
rect 30940 45836 31108 45892
rect 31164 48244 31220 48254
rect 31164 48130 31220 48188
rect 31164 48078 31166 48130
rect 31218 48078 31220 48130
rect 30380 39394 30436 39406
rect 30380 39342 30382 39394
rect 30434 39342 30436 39394
rect 30380 39060 30436 39342
rect 30492 39060 30548 39070
rect 30436 39058 30548 39060
rect 30436 39006 30494 39058
rect 30546 39006 30548 39058
rect 30436 39004 30548 39006
rect 30380 38928 30436 39004
rect 30492 38994 30548 39004
rect 30604 38668 30660 40684
rect 30940 40628 30996 45836
rect 31052 45668 31108 45678
rect 31052 45218 31108 45612
rect 31052 45166 31054 45218
rect 31106 45166 31108 45218
rect 31052 45154 31108 45166
rect 31164 45556 31220 48078
rect 31388 46900 31444 51100
rect 31724 50372 31780 51438
rect 31948 50820 32004 51886
rect 31948 50754 32004 50764
rect 32060 50484 32116 50494
rect 31724 50306 31780 50316
rect 31948 50482 32116 50484
rect 31948 50430 32062 50482
rect 32114 50430 32116 50482
rect 31948 50428 32116 50430
rect 31948 50034 32004 50428
rect 32060 50418 32116 50428
rect 32172 50484 32228 52780
rect 32172 50418 32228 50428
rect 31948 49982 31950 50034
rect 32002 49982 32004 50034
rect 31948 49970 32004 49982
rect 32060 50148 32116 50158
rect 32060 49922 32116 50092
rect 32060 49870 32062 49922
rect 32114 49870 32116 49922
rect 31836 49700 31892 49710
rect 31836 49606 31892 49644
rect 31836 49028 31892 49038
rect 31500 48916 31556 48926
rect 31500 48822 31556 48860
rect 31836 48466 31892 48972
rect 31836 48414 31838 48466
rect 31890 48414 31892 48466
rect 31836 48356 31892 48414
rect 31836 48290 31892 48300
rect 31948 47572 32004 47582
rect 31948 47478 32004 47516
rect 31500 47236 31556 47246
rect 31500 47142 31556 47180
rect 31388 46834 31444 46844
rect 32060 46788 32116 49870
rect 32284 49140 32340 54684
rect 32620 54514 32676 54526
rect 32620 54462 32622 54514
rect 32674 54462 32676 54514
rect 32620 53172 32676 54462
rect 33292 53732 33348 55916
rect 33404 55074 33460 55086
rect 33404 55022 33406 55074
rect 33458 55022 33460 55074
rect 33404 54068 33460 55022
rect 33852 55076 33908 58156
rect 34972 56196 35028 59200
rect 38220 58548 38276 58558
rect 36540 56420 36596 56430
rect 35196 56196 35252 56206
rect 34972 56194 35252 56196
rect 34972 56142 35198 56194
rect 35250 56142 35252 56194
rect 34972 56140 35252 56142
rect 35196 56130 35252 56140
rect 34412 56084 34468 56094
rect 34412 55990 34468 56028
rect 36092 56082 36148 56094
rect 36092 56030 36094 56082
rect 36146 56030 36148 56082
rect 33964 55970 34020 55982
rect 33964 55918 33966 55970
rect 34018 55918 34020 55970
rect 33964 55412 34020 55918
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 36092 55468 36148 56030
rect 33964 55346 34020 55356
rect 35756 55412 36148 55468
rect 34300 55300 34356 55310
rect 34300 55206 34356 55244
rect 35756 55186 35812 55412
rect 36540 55410 36596 56364
rect 36988 55972 37044 55982
rect 36988 55878 37044 55916
rect 37548 55970 37604 55982
rect 37548 55918 37550 55970
rect 37602 55918 37604 55970
rect 37548 55468 37604 55918
rect 37996 55970 38052 55982
rect 37996 55918 37998 55970
rect 38050 55918 38052 55970
rect 37996 55748 38052 55918
rect 37996 55682 38052 55692
rect 36540 55358 36542 55410
rect 36594 55358 36596 55410
rect 36540 55346 36596 55358
rect 37100 55412 37604 55468
rect 38220 55468 38276 58492
rect 40124 58324 40180 58334
rect 38668 57876 38724 57886
rect 38332 57652 38388 57662
rect 38332 56306 38388 57596
rect 38332 56254 38334 56306
rect 38386 56254 38388 56306
rect 38332 56242 38388 56254
rect 37884 55412 37940 55422
rect 38220 55412 38388 55468
rect 35756 55134 35758 55186
rect 35810 55134 35812 55186
rect 35756 55122 35812 55134
rect 36092 55188 36148 55198
rect 36092 55094 36148 55132
rect 33964 55076 34020 55086
rect 33852 55074 34020 55076
rect 33852 55022 33966 55074
rect 34018 55022 34020 55074
rect 33852 55020 34020 55022
rect 33852 54516 33908 55020
rect 33964 55010 34020 55020
rect 34860 55074 34916 55086
rect 34860 55022 34862 55074
rect 34914 55022 34916 55074
rect 33852 54450 33908 54460
rect 34412 54626 34468 54638
rect 34412 54574 34414 54626
rect 34466 54574 34468 54626
rect 33516 54402 33572 54414
rect 33516 54350 33518 54402
rect 33570 54350 33572 54402
rect 33516 54180 33572 54350
rect 34076 54404 34132 54414
rect 33516 54124 33796 54180
rect 33404 54002 33460 54012
rect 33180 53676 33348 53732
rect 33404 53842 33460 53854
rect 33404 53790 33406 53842
rect 33458 53790 33460 53842
rect 33404 53732 33460 53790
rect 32732 53618 32788 53630
rect 32732 53566 32734 53618
rect 32786 53566 32788 53618
rect 32732 53284 32788 53566
rect 32732 53218 32788 53228
rect 32620 53106 32676 53116
rect 32620 52836 32676 52846
rect 32396 52834 32676 52836
rect 32396 52782 32622 52834
rect 32674 52782 32676 52834
rect 32396 52780 32676 52782
rect 32396 52052 32452 52780
rect 32620 52770 32676 52780
rect 33068 52388 33124 52398
rect 32508 52386 33124 52388
rect 32508 52334 33070 52386
rect 33122 52334 33124 52386
rect 32508 52332 33124 52334
rect 32508 52162 32564 52332
rect 33068 52322 33124 52332
rect 32508 52110 32510 52162
rect 32562 52110 32564 52162
rect 32508 52098 32564 52110
rect 32396 51986 32452 51996
rect 32956 52052 33012 52062
rect 32956 51958 33012 51996
rect 33068 51938 33124 51950
rect 33068 51886 33070 51938
rect 33122 51886 33124 51938
rect 32396 51828 32452 51838
rect 32396 51154 32452 51772
rect 33068 51828 33124 51886
rect 33068 51762 33124 51772
rect 32396 51102 32398 51154
rect 32450 51102 32452 51154
rect 32396 50594 32452 51102
rect 32396 50542 32398 50594
rect 32450 50542 32452 50594
rect 32396 49250 32452 50542
rect 32508 51380 32564 51390
rect 32508 50370 32564 51324
rect 32732 51156 32788 51166
rect 32732 51062 32788 51100
rect 32732 50594 32788 50606
rect 32732 50542 32734 50594
rect 32786 50542 32788 50594
rect 32508 50318 32510 50370
rect 32562 50318 32564 50370
rect 32508 50306 32564 50318
rect 32620 50372 32676 50382
rect 32396 49198 32398 49250
rect 32450 49198 32452 49250
rect 32396 49186 32452 49198
rect 32620 50034 32676 50316
rect 32620 49982 32622 50034
rect 32674 49982 32676 50034
rect 31948 46732 32116 46788
rect 32172 49084 32340 49140
rect 31276 46676 31332 46686
rect 31276 46582 31332 46620
rect 31724 46562 31780 46574
rect 31724 46510 31726 46562
rect 31778 46510 31780 46562
rect 31724 46452 31780 46510
rect 31388 45890 31444 45902
rect 31388 45838 31390 45890
rect 31442 45838 31444 45890
rect 31388 45668 31444 45838
rect 31388 45602 31444 45612
rect 31612 45890 31668 45902
rect 31612 45838 31614 45890
rect 31666 45838 31668 45890
rect 31164 44434 31220 45500
rect 31612 45108 31668 45838
rect 31724 45892 31780 46396
rect 31948 46340 32004 46732
rect 32060 46564 32116 46574
rect 32060 46470 32116 46508
rect 31948 46284 32116 46340
rect 31724 45826 31780 45836
rect 31836 45890 31892 45902
rect 31836 45838 31838 45890
rect 31890 45838 31892 45890
rect 31388 45052 31668 45108
rect 31724 45666 31780 45678
rect 31724 45614 31726 45666
rect 31778 45614 31780 45666
rect 31388 44994 31444 45052
rect 31388 44942 31390 44994
rect 31442 44942 31444 44994
rect 31276 44884 31332 44894
rect 31276 44790 31332 44828
rect 31164 44382 31166 44434
rect 31218 44382 31220 44434
rect 31164 44370 31220 44382
rect 31388 44546 31444 44942
rect 31388 44494 31390 44546
rect 31442 44494 31444 44546
rect 31164 43428 31220 43438
rect 31052 43426 31220 43428
rect 31052 43374 31166 43426
rect 31218 43374 31220 43426
rect 31052 43372 31220 43374
rect 31052 41858 31108 43372
rect 31164 43362 31220 43372
rect 31052 41806 31054 41858
rect 31106 41806 31108 41858
rect 31052 41524 31108 41806
rect 31052 41458 31108 41468
rect 31052 40964 31108 40974
rect 31052 40870 31108 40908
rect 30268 35522 30324 35532
rect 30380 38612 30660 38668
rect 30716 40572 30996 40628
rect 30380 34356 30436 38612
rect 30604 38052 30660 38062
rect 30604 37266 30660 37996
rect 30604 37214 30606 37266
rect 30658 37214 30660 37266
rect 30604 37202 30660 37214
rect 30492 36484 30548 36522
rect 30492 36418 30548 36428
rect 30604 36260 30660 36270
rect 30604 36166 30660 36204
rect 30716 35812 30772 40572
rect 31164 40516 31220 40526
rect 30828 40460 31164 40516
rect 30828 39506 30884 40460
rect 31164 40384 31220 40460
rect 31388 40292 31444 44494
rect 31612 44772 31668 44782
rect 31500 43428 31556 43438
rect 31500 43334 31556 43372
rect 31164 40236 31444 40292
rect 31500 42754 31556 42766
rect 31500 42702 31502 42754
rect 31554 42702 31556 42754
rect 30940 39844 30996 39854
rect 30940 39750 30996 39788
rect 30828 39454 30830 39506
rect 30882 39454 30884 39506
rect 30828 38948 30884 39454
rect 30828 38892 30996 38948
rect 30828 38724 30884 38734
rect 30828 38050 30884 38668
rect 30828 37998 30830 38050
rect 30882 37998 30884 38050
rect 30828 37940 30884 37998
rect 30828 37874 30884 37884
rect 30828 37042 30884 37054
rect 30828 36990 30830 37042
rect 30882 36990 30884 37042
rect 30828 36596 30884 36990
rect 30828 36530 30884 36540
rect 30716 35756 30884 35812
rect 30716 35588 30772 35598
rect 30716 35494 30772 35532
rect 30604 34690 30660 34702
rect 30604 34638 30606 34690
rect 30658 34638 30660 34690
rect 29708 33346 29876 33348
rect 29708 33294 29710 33346
rect 29762 33294 29876 33346
rect 29708 33292 29876 33294
rect 29932 33516 30212 33572
rect 30268 34300 30436 34356
rect 30492 34468 30548 34478
rect 30268 33572 30324 34300
rect 30380 34132 30436 34142
rect 30380 34038 30436 34076
rect 29708 33282 29764 33292
rect 29820 33124 29876 33134
rect 29372 33122 29876 33124
rect 29372 33070 29822 33122
rect 29874 33070 29876 33122
rect 29372 33068 29876 33070
rect 29372 32786 29428 33068
rect 29820 33058 29876 33068
rect 29932 32900 29988 33516
rect 30268 33506 30324 33516
rect 30044 33348 30100 33358
rect 30380 33348 30436 33358
rect 30044 33346 30436 33348
rect 30044 33294 30046 33346
rect 30098 33294 30382 33346
rect 30434 33294 30436 33346
rect 30044 33292 30436 33294
rect 30044 33282 30100 33292
rect 30380 33282 30436 33292
rect 30492 33124 30548 34412
rect 30604 33684 30660 34638
rect 30604 33618 30660 33628
rect 30828 33348 30884 35756
rect 30940 34356 30996 38892
rect 31052 38834 31108 38846
rect 31052 38782 31054 38834
rect 31106 38782 31108 38834
rect 31052 38724 31108 38782
rect 31052 38658 31108 38668
rect 31052 38500 31108 38510
rect 31052 38274 31108 38444
rect 31052 38222 31054 38274
rect 31106 38222 31108 38274
rect 31052 38210 31108 38222
rect 31164 37268 31220 40236
rect 31500 39844 31556 42702
rect 31612 42644 31668 44716
rect 31724 44436 31780 45614
rect 31836 44884 31892 45838
rect 31836 44818 31892 44828
rect 31724 44380 32004 44436
rect 31948 44322 32004 44380
rect 31948 44270 31950 44322
rect 32002 44270 32004 44322
rect 31948 44258 32004 44270
rect 32060 44212 32116 46284
rect 32172 45668 32228 49084
rect 32284 48914 32340 48926
rect 32284 48862 32286 48914
rect 32338 48862 32340 48914
rect 32284 48692 32340 48862
rect 32620 48916 32676 49982
rect 32732 49700 32788 50542
rect 32732 49634 32788 49644
rect 32620 48850 32676 48860
rect 32732 49140 32788 49150
rect 33180 49140 33236 53676
rect 33404 53666 33460 53676
rect 33628 53730 33684 53742
rect 33628 53678 33630 53730
rect 33682 53678 33684 53730
rect 33404 53396 33460 53406
rect 33404 52500 33460 53340
rect 33404 52434 33460 52444
rect 33628 52722 33684 53678
rect 33740 53396 33796 54124
rect 33964 53956 34020 53966
rect 34076 53956 34132 54348
rect 34188 54402 34244 54414
rect 34188 54350 34190 54402
rect 34242 54350 34244 54402
rect 34188 54292 34244 54350
rect 34188 54226 34244 54236
rect 34188 53956 34244 53966
rect 34076 53954 34244 53956
rect 34076 53902 34190 53954
rect 34242 53902 34244 53954
rect 34076 53900 34244 53902
rect 33964 53842 34020 53900
rect 34188 53890 34244 53900
rect 33964 53790 33966 53842
rect 34018 53790 34020 53842
rect 33964 53778 34020 53790
rect 33740 53330 33796 53340
rect 33964 53618 34020 53630
rect 33964 53566 33966 53618
rect 34018 53566 34020 53618
rect 33740 53172 33796 53182
rect 33740 53078 33796 53116
rect 33628 52670 33630 52722
rect 33682 52670 33684 52722
rect 33292 52276 33348 52286
rect 33292 50148 33348 52220
rect 33292 50082 33348 50092
rect 33404 51492 33460 51502
rect 33404 50482 33460 51436
rect 33404 50430 33406 50482
rect 33458 50430 33460 50482
rect 33180 49084 33348 49140
rect 32396 48804 32452 48814
rect 32396 48802 32564 48804
rect 32396 48750 32398 48802
rect 32450 48750 32564 48802
rect 32396 48748 32564 48750
rect 32396 48738 32452 48748
rect 32284 48580 32340 48636
rect 32284 48524 32452 48580
rect 32284 48356 32340 48366
rect 32284 48262 32340 48300
rect 32396 47236 32452 48524
rect 32508 47796 32564 48748
rect 32732 48466 32788 49084
rect 33068 49028 33124 49038
rect 33068 48934 33124 48972
rect 33180 48916 33236 48926
rect 33180 48822 33236 48860
rect 32732 48414 32734 48466
rect 32786 48414 32788 48466
rect 32732 48402 32788 48414
rect 32844 48692 32900 48702
rect 32844 48354 32900 48636
rect 32844 48302 32846 48354
rect 32898 48302 32900 48354
rect 32844 48290 32900 48302
rect 32620 48244 32676 48254
rect 32620 48150 32676 48188
rect 32508 47740 32900 47796
rect 32844 47460 32900 47740
rect 32844 47328 32900 47404
rect 33180 47348 33236 47358
rect 33180 47254 33236 47292
rect 32396 47180 32676 47236
rect 32620 47068 32676 47180
rect 32844 47124 32900 47134
rect 32508 47012 32564 47022
rect 32620 47012 32788 47068
rect 32508 46898 32564 46956
rect 32508 46846 32510 46898
rect 32562 46846 32564 46898
rect 32508 46834 32564 46846
rect 32284 45668 32340 45678
rect 32172 45666 32340 45668
rect 32172 45614 32286 45666
rect 32338 45614 32340 45666
rect 32172 45612 32340 45614
rect 32284 44212 32340 45612
rect 32620 45106 32676 45118
rect 32620 45054 32622 45106
rect 32674 45054 32676 45106
rect 32620 44772 32676 45054
rect 32732 44882 32788 47012
rect 32732 44830 32734 44882
rect 32786 44830 32788 44882
rect 32732 44818 32788 44830
rect 32060 44210 32228 44212
rect 32060 44158 32062 44210
rect 32114 44158 32228 44210
rect 32060 44156 32228 44158
rect 32060 44146 32116 44156
rect 32172 44100 32228 44156
rect 32284 44146 32340 44156
rect 32396 44716 32676 44772
rect 31724 43652 31780 43662
rect 31724 42866 31780 43596
rect 31724 42814 31726 42866
rect 31778 42814 31780 42866
rect 31724 42802 31780 42814
rect 31836 43428 31892 43438
rect 31836 42754 31892 43372
rect 31836 42702 31838 42754
rect 31890 42702 31892 42754
rect 31836 42690 31892 42702
rect 32060 43426 32116 43438
rect 32060 43374 32062 43426
rect 32114 43374 32116 43426
rect 32060 42980 32116 43374
rect 32060 42754 32116 42924
rect 32060 42702 32062 42754
rect 32114 42702 32116 42754
rect 32060 42690 32116 42702
rect 31612 42588 31780 42644
rect 31500 39618 31556 39788
rect 31500 39566 31502 39618
rect 31554 39566 31556 39618
rect 31500 39554 31556 39566
rect 31612 41970 31668 41982
rect 31612 41918 31614 41970
rect 31666 41918 31668 41970
rect 31388 38722 31444 38734
rect 31388 38670 31390 38722
rect 31442 38670 31444 38722
rect 31276 38610 31332 38622
rect 31276 38558 31278 38610
rect 31330 38558 31332 38610
rect 31276 38500 31332 38558
rect 31276 38434 31332 38444
rect 31388 37940 31444 38670
rect 31500 38276 31556 38286
rect 31612 38276 31668 41918
rect 31500 38274 31668 38276
rect 31500 38222 31502 38274
rect 31554 38222 31668 38274
rect 31500 38220 31668 38222
rect 31500 38210 31556 38220
rect 31388 37874 31444 37884
rect 30940 34290 30996 34300
rect 31052 37212 31220 37268
rect 31052 33796 31108 37212
rect 31164 37044 31220 37054
rect 31164 37042 31444 37044
rect 31164 36990 31166 37042
rect 31218 36990 31444 37042
rect 31164 36988 31444 36990
rect 31164 36978 31220 36988
rect 31276 36820 31332 36830
rect 31276 36706 31332 36764
rect 31276 36654 31278 36706
rect 31330 36654 31332 36706
rect 31276 36642 31332 36654
rect 31388 36594 31444 36988
rect 31388 36542 31390 36594
rect 31442 36542 31444 36594
rect 31388 36530 31444 36542
rect 31388 35588 31444 35598
rect 31388 34914 31444 35532
rect 31724 34916 31780 42588
rect 32172 42532 32228 44044
rect 32284 43428 32340 43438
rect 32284 43334 32340 43372
rect 32060 42476 32228 42532
rect 31836 42082 31892 42094
rect 31836 42030 31838 42082
rect 31890 42030 31892 42082
rect 31836 41524 31892 42030
rect 31948 42084 32004 42122
rect 31948 42018 32004 42028
rect 31836 41458 31892 41468
rect 31836 39508 31892 39518
rect 31836 39414 31892 39452
rect 32060 39284 32116 42476
rect 32396 42308 32452 44716
rect 32620 44324 32676 44334
rect 32844 44324 32900 47068
rect 33068 47124 33124 47134
rect 32956 46004 33012 46014
rect 32956 45910 33012 45948
rect 32956 44548 33012 44558
rect 32956 44454 33012 44492
rect 32620 44322 32900 44324
rect 32620 44270 32622 44322
rect 32674 44270 32900 44322
rect 32620 44268 32900 44270
rect 32620 43652 32676 44268
rect 32620 43586 32676 43596
rect 32620 43428 32676 43438
rect 32620 43334 32676 43372
rect 33068 43204 33124 47068
rect 33180 47012 33236 47022
rect 33180 45444 33236 46956
rect 33180 45378 33236 45388
rect 33292 44548 33348 49084
rect 33404 46004 33460 50430
rect 33516 49698 33572 49710
rect 33516 49646 33518 49698
rect 33570 49646 33572 49698
rect 33516 49028 33572 49646
rect 33628 49138 33684 52670
rect 33964 52946 34020 53566
rect 34412 53396 34468 54574
rect 34636 54628 34692 54638
rect 34636 53844 34692 54572
rect 34860 54292 34916 55022
rect 35196 55076 35252 55086
rect 35196 54982 35252 55020
rect 35868 55076 35924 55086
rect 34860 54226 34916 54236
rect 35644 54514 35700 54526
rect 35644 54462 35646 54514
rect 35698 54462 35700 54514
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 34636 53730 34692 53788
rect 34636 53678 34638 53730
rect 34690 53678 34692 53730
rect 34636 53666 34692 53678
rect 34412 53330 34468 53340
rect 34748 53508 34804 53518
rect 33964 52894 33966 52946
rect 34018 52894 34020 52946
rect 33740 52050 33796 52062
rect 33740 51998 33742 52050
rect 33794 51998 33796 52050
rect 33740 51828 33796 51998
rect 33740 51762 33796 51772
rect 33852 51938 33908 51950
rect 33852 51886 33854 51938
rect 33906 51886 33908 51938
rect 33852 51492 33908 51886
rect 33852 51398 33908 51436
rect 33740 51380 33796 51390
rect 33740 51286 33796 51324
rect 33964 51268 34020 52894
rect 34524 52834 34580 52846
rect 34524 52782 34526 52834
rect 34578 52782 34580 52834
rect 34412 52276 34468 52286
rect 34412 52182 34468 52220
rect 34076 51938 34132 51950
rect 34076 51886 34078 51938
rect 34130 51886 34132 51938
rect 34076 51380 34132 51886
rect 34524 51492 34580 52782
rect 34748 51602 34804 53452
rect 35084 53506 35140 53518
rect 35084 53454 35086 53506
rect 35138 53454 35140 53506
rect 35084 53396 35140 53454
rect 35644 53508 35700 54462
rect 35868 53730 35924 55020
rect 36988 55076 37044 55086
rect 36204 54740 36260 54750
rect 36204 54646 36260 54684
rect 36988 54738 37044 55020
rect 36988 54686 36990 54738
rect 37042 54686 37044 54738
rect 36988 54674 37044 54686
rect 36876 54514 36932 54526
rect 36876 54462 36878 54514
rect 36930 54462 36932 54514
rect 35868 53678 35870 53730
rect 35922 53678 35924 53730
rect 35868 53666 35924 53678
rect 35980 54292 36036 54302
rect 35644 53414 35700 53452
rect 35756 53506 35812 53518
rect 35756 53454 35758 53506
rect 35810 53454 35812 53506
rect 35084 53330 35140 53340
rect 35756 53284 35812 53454
rect 35980 53284 36036 54236
rect 36092 53506 36148 53518
rect 36092 53454 36094 53506
rect 36146 53454 36148 53506
rect 36092 53396 36148 53454
rect 36092 53330 36148 53340
rect 36764 53506 36820 53518
rect 36764 53454 36766 53506
rect 36818 53454 36820 53506
rect 36764 53396 36820 53454
rect 36876 53508 36932 54462
rect 36988 54292 37044 54302
rect 36988 54198 37044 54236
rect 36876 53442 36932 53452
rect 36764 53330 36820 53340
rect 35644 53228 35812 53284
rect 35868 53228 36036 53284
rect 35644 53058 35700 53228
rect 35644 53006 35646 53058
rect 35698 53006 35700 53058
rect 35644 52994 35700 53006
rect 35756 53060 35812 53070
rect 35868 53060 35924 53228
rect 36764 53172 36820 53182
rect 36764 53078 36820 53116
rect 35756 53058 35924 53060
rect 35756 53006 35758 53058
rect 35810 53006 35924 53058
rect 35756 53004 35924 53006
rect 36540 53060 36596 53070
rect 35756 52994 35812 53004
rect 35980 52948 36036 52958
rect 36428 52948 36484 52958
rect 35980 52854 36036 52892
rect 36316 52946 36484 52948
rect 36316 52894 36430 52946
rect 36482 52894 36484 52946
rect 36316 52892 36484 52894
rect 35196 52836 35252 52846
rect 34748 51550 34750 51602
rect 34802 51550 34804 51602
rect 34748 51538 34804 51550
rect 35084 52834 35252 52836
rect 35084 52782 35198 52834
rect 35250 52782 35252 52834
rect 35084 52780 35252 52782
rect 34524 51426 34580 51436
rect 34076 51314 34132 51324
rect 34860 51378 34916 51390
rect 34860 51326 34862 51378
rect 34914 51326 34916 51378
rect 33964 51202 34020 51212
rect 34860 51268 34916 51326
rect 34860 51202 34916 51212
rect 35084 51156 35140 52780
rect 35196 52770 35252 52780
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35532 52274 35588 52286
rect 35532 52222 35534 52274
rect 35586 52222 35588 52274
rect 35532 52164 35588 52222
rect 35532 52098 35588 52108
rect 35868 52276 35924 52286
rect 35868 52162 35924 52220
rect 35868 52110 35870 52162
rect 35922 52110 35924 52162
rect 35868 51604 35924 52110
rect 36316 52162 36372 52892
rect 36428 52882 36484 52892
rect 36540 52388 36596 53004
rect 36316 52110 36318 52162
rect 36370 52110 36372 52162
rect 36316 52098 36372 52110
rect 36428 52332 36596 52388
rect 35980 51604 36036 51614
rect 35868 51602 36036 51604
rect 35868 51550 35982 51602
rect 36034 51550 36036 51602
rect 35868 51548 36036 51550
rect 35980 51538 36036 51548
rect 35644 51380 35700 51390
rect 35644 51286 35700 51324
rect 35420 51266 35476 51278
rect 35420 51214 35422 51266
rect 35474 51214 35476 51266
rect 35420 51156 35476 51214
rect 35084 51100 35476 51156
rect 36092 51156 36148 51166
rect 34188 50820 34244 50830
rect 34188 50726 34244 50764
rect 34524 50820 34580 50830
rect 34524 50726 34580 50764
rect 34524 50596 34580 50606
rect 34524 50502 34580 50540
rect 35084 50482 35140 51100
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35532 50708 35588 50718
rect 35084 50430 35086 50482
rect 35138 50430 35140 50482
rect 35084 50428 35140 50430
rect 34748 50372 35140 50428
rect 35196 50596 35252 50606
rect 33964 49700 34020 49710
rect 33964 49606 34020 49644
rect 34748 49698 34804 50372
rect 35196 49700 35252 50540
rect 35532 50594 35588 50652
rect 36092 50706 36148 51100
rect 36092 50654 36094 50706
rect 36146 50654 36148 50706
rect 36092 50642 36148 50654
rect 36428 50708 36484 52332
rect 36764 52164 36820 52174
rect 36764 52070 36820 52108
rect 36764 51490 36820 51502
rect 36764 51438 36766 51490
rect 36818 51438 36820 51490
rect 36652 51268 36708 51278
rect 36540 51154 36596 51166
rect 36540 51102 36542 51154
rect 36594 51102 36596 51154
rect 36540 50820 36596 51102
rect 36540 50754 36596 50764
rect 36428 50642 36484 50652
rect 35532 50542 35534 50594
rect 35586 50542 35588 50594
rect 35532 50428 35588 50542
rect 36204 50596 36260 50606
rect 36204 50502 36260 50540
rect 36540 50484 36596 50494
rect 35532 50372 35812 50428
rect 36540 50390 36596 50428
rect 34748 49646 34750 49698
rect 34802 49646 34804 49698
rect 34748 49588 34804 49646
rect 34300 49532 34804 49588
rect 35084 49698 35252 49700
rect 35084 49646 35198 49698
rect 35250 49646 35252 49698
rect 35084 49644 35252 49646
rect 33628 49086 33630 49138
rect 33682 49086 33684 49138
rect 33628 49074 33684 49086
rect 33852 49140 33908 49150
rect 33852 49046 33908 49084
rect 33516 48962 33572 48972
rect 34188 49028 34244 49038
rect 34188 48934 34244 48972
rect 33852 48692 33908 48702
rect 33852 48356 33908 48636
rect 33740 48354 33908 48356
rect 33740 48302 33854 48354
rect 33906 48302 33908 48354
rect 33740 48300 33908 48302
rect 33628 48244 33684 48254
rect 33628 47348 33684 48188
rect 33740 47458 33796 48300
rect 33852 48290 33908 48300
rect 33964 48580 34020 48590
rect 33964 48354 34020 48524
rect 33964 48302 33966 48354
rect 34018 48302 34020 48354
rect 33964 48290 34020 48302
rect 34300 48020 34356 49532
rect 34972 49140 35028 49150
rect 34860 48580 34916 48590
rect 34860 48466 34916 48524
rect 34860 48414 34862 48466
rect 34914 48414 34916 48466
rect 33964 47964 34356 48020
rect 34412 48020 34468 48030
rect 34412 48018 34804 48020
rect 34412 47966 34414 48018
rect 34466 47966 34804 48018
rect 34412 47964 34804 47966
rect 33740 47406 33742 47458
rect 33794 47406 33796 47458
rect 33740 47394 33796 47406
rect 33852 47460 33908 47470
rect 33852 47366 33908 47404
rect 33628 47282 33684 47292
rect 33628 47124 33684 47134
rect 33628 46898 33684 47068
rect 33628 46846 33630 46898
rect 33682 46846 33684 46898
rect 33628 46834 33684 46846
rect 33964 46900 34020 47964
rect 34412 47954 34468 47964
rect 34300 47684 34356 47694
rect 34300 47458 34356 47628
rect 34300 47406 34302 47458
rect 34354 47406 34356 47458
rect 34076 47348 34132 47358
rect 34132 47292 34244 47348
rect 34076 47216 34132 47292
rect 33964 46844 34132 46900
rect 33964 46562 34020 46574
rect 33964 46510 33966 46562
rect 34018 46510 34020 46562
rect 33460 45948 33684 46004
rect 33404 45938 33460 45948
rect 33516 45778 33572 45790
rect 33516 45726 33518 45778
rect 33570 45726 33572 45778
rect 32620 43148 33124 43204
rect 33180 44492 33348 44548
rect 33404 45444 33460 45454
rect 32284 42252 32452 42308
rect 32508 42420 32564 42430
rect 32284 41970 32340 42252
rect 32284 41918 32286 41970
rect 32338 41918 32340 41970
rect 32172 41524 32228 41534
rect 32172 41186 32228 41468
rect 32172 41134 32174 41186
rect 32226 41134 32228 41186
rect 32172 41122 32228 41134
rect 32284 41074 32340 41918
rect 32396 42084 32452 42094
rect 32396 41858 32452 42028
rect 32396 41806 32398 41858
rect 32450 41806 32452 41858
rect 32396 41794 32452 41806
rect 32508 41186 32564 42364
rect 32508 41134 32510 41186
rect 32562 41134 32564 41186
rect 32508 41122 32564 41134
rect 32284 41022 32286 41074
rect 32338 41022 32340 41074
rect 32284 39508 32340 41022
rect 32620 40964 32676 43148
rect 33068 42642 33124 42654
rect 33068 42590 33070 42642
rect 33122 42590 33124 42642
rect 32844 41972 32900 41982
rect 32284 39442 32340 39452
rect 32508 40908 32676 40964
rect 32732 41916 32844 41972
rect 32396 39394 32452 39406
rect 32396 39342 32398 39394
rect 32450 39342 32452 39394
rect 32396 39284 32452 39342
rect 32060 39228 32452 39284
rect 32172 39060 32228 39070
rect 31948 38162 32004 38174
rect 31948 38110 31950 38162
rect 32002 38110 32004 38162
rect 31948 37266 32004 38110
rect 32060 37940 32116 37950
rect 32060 37846 32116 37884
rect 31948 37214 31950 37266
rect 32002 37214 32004 37266
rect 31948 37202 32004 37214
rect 31948 36596 32004 36606
rect 31948 36502 32004 36540
rect 32060 35700 32116 35710
rect 32060 35026 32116 35644
rect 32060 34974 32062 35026
rect 32114 34974 32116 35026
rect 32060 34962 32116 34974
rect 31388 34862 31390 34914
rect 31442 34862 31444 34914
rect 31388 34850 31444 34862
rect 31500 34860 31780 34916
rect 31836 34914 31892 34926
rect 31836 34862 31838 34914
rect 31890 34862 31892 34914
rect 31276 34356 31332 34366
rect 31164 34020 31220 34030
rect 31164 33926 31220 33964
rect 31052 33740 31220 33796
rect 30828 33282 30884 33292
rect 31052 33572 31108 33582
rect 31052 33346 31108 33516
rect 31052 33294 31054 33346
rect 31106 33294 31108 33346
rect 31052 33282 31108 33294
rect 30828 33124 30884 33134
rect 29372 32734 29374 32786
rect 29426 32734 29428 32786
rect 29372 32722 29428 32734
rect 29596 32844 29988 32900
rect 30156 33068 30548 33124
rect 30716 33122 30884 33124
rect 30716 33070 30830 33122
rect 30882 33070 30884 33122
rect 30716 33068 30884 33070
rect 29148 32050 29204 32060
rect 28700 31276 29092 31332
rect 29260 31892 29316 31902
rect 28476 29652 28532 29662
rect 28476 29558 28532 29596
rect 28476 27970 28532 27982
rect 28476 27918 28478 27970
rect 28530 27918 28532 27970
rect 28476 26292 28532 27918
rect 28588 27188 28644 27198
rect 28588 27094 28644 27132
rect 28700 26516 28756 31276
rect 29036 29988 29092 29998
rect 28812 29540 28868 29550
rect 28812 28754 28868 29484
rect 28812 28702 28814 28754
rect 28866 28702 28868 28754
rect 28812 28690 28868 28702
rect 28700 26450 28756 26460
rect 28476 26226 28532 26236
rect 28364 25890 28420 25900
rect 27580 25676 27748 25732
rect 27020 25618 27636 25620
rect 27020 25566 27022 25618
rect 27074 25566 27636 25618
rect 27020 25564 27636 25566
rect 27020 25554 27076 25564
rect 27580 25506 27636 25564
rect 27580 25454 27582 25506
rect 27634 25454 27636 25506
rect 27580 25442 27636 25454
rect 26908 25116 27188 25172
rect 26460 24882 26516 24892
rect 27020 24948 27076 24958
rect 26908 24836 26964 24846
rect 26908 24742 26964 24780
rect 27020 24834 27076 24892
rect 27020 24782 27022 24834
rect 27074 24782 27076 24834
rect 27020 24770 27076 24782
rect 26348 24724 26404 24734
rect 26684 24724 26740 24734
rect 26348 24722 26740 24724
rect 26348 24670 26350 24722
rect 26402 24670 26686 24722
rect 26738 24670 26740 24722
rect 26348 24668 26740 24670
rect 26348 24658 26404 24668
rect 26124 23986 26180 23996
rect 26124 23828 26180 23838
rect 26012 23826 26180 23828
rect 26012 23774 26126 23826
rect 26178 23774 26180 23826
rect 26012 23772 26180 23774
rect 26124 23762 26180 23772
rect 26236 23604 26292 23614
rect 26124 23492 26180 23502
rect 25676 23156 25732 23166
rect 25676 23062 25732 23100
rect 26012 23156 26068 23166
rect 26012 22594 26068 23100
rect 26012 22542 26014 22594
rect 26066 22542 26068 22594
rect 26012 22530 26068 22542
rect 26124 23154 26180 23436
rect 26124 23102 26126 23154
rect 26178 23102 26180 23154
rect 25116 21362 25508 21364
rect 25116 21310 25118 21362
rect 25170 21310 25508 21362
rect 25116 21308 25508 21310
rect 25676 22146 25732 22158
rect 25676 22094 25678 22146
rect 25730 22094 25732 22146
rect 25116 21298 25172 21308
rect 24668 20638 24670 20690
rect 24722 20638 24724 20690
rect 24108 20402 24164 20412
rect 24444 20580 24500 20590
rect 24332 20132 24388 20142
rect 24332 20038 24388 20076
rect 23548 19908 23604 19918
rect 23548 19814 23604 19852
rect 24220 19794 24276 19806
rect 24220 19742 24222 19794
rect 24274 19742 24276 19794
rect 24108 19234 24164 19246
rect 24108 19182 24110 19234
rect 24162 19182 24164 19234
rect 23548 19012 23604 19022
rect 23548 19010 23716 19012
rect 23548 18958 23550 19010
rect 23602 18958 23716 19010
rect 23548 18956 23716 18958
rect 23548 18946 23604 18956
rect 23548 18562 23604 18574
rect 23548 18510 23550 18562
rect 23602 18510 23604 18562
rect 23548 16100 23604 18510
rect 23660 16996 23716 18956
rect 24108 18338 24164 19182
rect 24220 18674 24276 19742
rect 24444 19348 24500 20524
rect 24444 19234 24500 19292
rect 24444 19182 24446 19234
rect 24498 19182 24500 19234
rect 24444 19170 24500 19182
rect 24668 18788 24724 20638
rect 25004 20692 25060 20702
rect 25004 20598 25060 20636
rect 25564 20692 25620 20702
rect 25564 20598 25620 20636
rect 24220 18622 24222 18674
rect 24274 18622 24276 18674
rect 24220 18564 24276 18622
rect 24220 18498 24276 18508
rect 24332 18732 24724 18788
rect 24780 20468 24836 20478
rect 24780 20242 24836 20412
rect 24780 20190 24782 20242
rect 24834 20190 24836 20242
rect 24108 18286 24110 18338
rect 24162 18286 24164 18338
rect 24108 18274 24164 18286
rect 24332 18340 24388 18732
rect 24780 18676 24836 20190
rect 25564 20132 25620 20142
rect 25564 20038 25620 20076
rect 25004 19124 25060 19134
rect 25004 19122 25172 19124
rect 25004 19070 25006 19122
rect 25058 19070 25172 19122
rect 25004 19068 25172 19070
rect 25004 19058 25060 19068
rect 24892 18676 24948 18686
rect 24444 18674 24948 18676
rect 24444 18622 24894 18674
rect 24946 18622 24948 18674
rect 24444 18620 24948 18622
rect 24444 18562 24500 18620
rect 24892 18610 24948 18620
rect 24444 18510 24446 18562
rect 24498 18510 24500 18562
rect 24444 18498 24500 18510
rect 24332 17780 24388 18284
rect 23884 17668 23940 17678
rect 23884 17574 23940 17612
rect 24108 17668 24164 17678
rect 24332 17668 24388 17724
rect 24108 17666 24388 17668
rect 24108 17614 24110 17666
rect 24162 17614 24388 17666
rect 24108 17612 24388 17614
rect 24556 18228 24612 18238
rect 24556 17666 24612 18172
rect 24556 17614 24558 17666
rect 24610 17614 24612 17666
rect 24108 17602 24164 17612
rect 24556 17602 24612 17614
rect 24892 17780 24948 17790
rect 24892 17666 24948 17724
rect 24892 17614 24894 17666
rect 24946 17614 24948 17666
rect 24668 17556 24724 17566
rect 23996 17444 24052 17454
rect 23996 17350 24052 17388
rect 23660 16930 23716 16940
rect 24220 16996 24276 17006
rect 24220 16902 24276 16940
rect 24668 16882 24724 17500
rect 24892 17220 24948 17614
rect 24892 17154 24948 17164
rect 24668 16830 24670 16882
rect 24722 16830 24724 16882
rect 24668 16818 24724 16830
rect 24668 16660 24724 16670
rect 23548 16034 23604 16044
rect 24108 16100 24164 16110
rect 23772 15874 23828 15886
rect 23772 15822 23774 15874
rect 23826 15822 23828 15874
rect 23772 15540 23828 15822
rect 24108 15652 24164 16044
rect 24668 15988 24724 16604
rect 24892 16212 24948 16222
rect 24892 16098 24948 16156
rect 24892 16046 24894 16098
rect 24946 16046 24948 16098
rect 24892 16034 24948 16046
rect 24108 15586 24164 15596
rect 24556 15986 24724 15988
rect 24556 15934 24670 15986
rect 24722 15934 24724 15986
rect 24556 15932 24724 15934
rect 23772 15474 23828 15484
rect 24556 15314 24612 15932
rect 24668 15922 24724 15932
rect 24556 15262 24558 15314
rect 24610 15262 24612 15314
rect 24556 15250 24612 15262
rect 24444 15204 24500 15242
rect 24444 15138 24500 15148
rect 23772 15090 23828 15102
rect 23772 15038 23774 15090
rect 23826 15038 23828 15090
rect 23436 14306 23492 14318
rect 23436 14254 23438 14306
rect 23490 14254 23492 14306
rect 23436 13972 23492 14254
rect 23436 13906 23492 13916
rect 23436 13636 23492 13646
rect 23436 11732 23492 13580
rect 23772 11844 23828 15038
rect 24220 14532 24276 14542
rect 24220 14438 24276 14476
rect 24780 14530 24836 14542
rect 24780 14478 24782 14530
rect 24834 14478 24836 14530
rect 24108 14420 24164 14430
rect 24108 14326 24164 14364
rect 24332 14308 24388 14318
rect 24332 14306 24500 14308
rect 24332 14254 24334 14306
rect 24386 14254 24500 14306
rect 24332 14252 24500 14254
rect 24332 14242 24388 14252
rect 24444 13972 24500 14252
rect 24780 14084 24836 14478
rect 24780 14018 24836 14028
rect 24556 13972 24612 13982
rect 24444 13916 24556 13972
rect 24556 13840 24612 13916
rect 24892 13858 24948 13870
rect 24892 13806 24894 13858
rect 24946 13806 24948 13858
rect 24892 13636 24948 13806
rect 24892 13570 24948 13580
rect 25116 13188 25172 19068
rect 25564 19010 25620 19022
rect 25564 18958 25566 19010
rect 25618 18958 25620 19010
rect 25564 18452 25620 18958
rect 25676 18788 25732 22094
rect 26124 21812 26180 23102
rect 26236 22484 26292 23548
rect 26460 23042 26516 24668
rect 26684 24658 26740 24668
rect 27132 23940 27188 25116
rect 27580 24948 27636 24958
rect 27692 24948 27748 25676
rect 28140 25730 28308 25732
rect 28140 25678 28142 25730
rect 28194 25678 28308 25730
rect 28140 25676 28308 25678
rect 28140 25666 28196 25676
rect 27804 25506 27860 25518
rect 27804 25454 27806 25506
rect 27858 25454 27860 25506
rect 27804 25284 27860 25454
rect 27804 25218 27860 25228
rect 28028 25506 28084 25518
rect 28028 25454 28030 25506
rect 28082 25454 28084 25506
rect 27636 24892 27748 24948
rect 27580 24816 27636 24892
rect 27804 24836 27860 24846
rect 27804 24388 27860 24780
rect 27916 24724 27972 24734
rect 27916 24630 27972 24668
rect 27804 24052 27860 24332
rect 27916 24052 27972 24062
rect 27804 24050 27972 24052
rect 27804 23998 27918 24050
rect 27970 23998 27972 24050
rect 27804 23996 27972 23998
rect 27916 23986 27972 23996
rect 26460 22990 26462 23042
rect 26514 22990 26516 23042
rect 26460 22978 26516 22990
rect 27020 23884 27188 23940
rect 26796 22484 26852 22494
rect 26236 22482 26852 22484
rect 26236 22430 26238 22482
rect 26290 22430 26798 22482
rect 26850 22430 26852 22482
rect 26236 22428 26852 22430
rect 26236 22418 26292 22428
rect 26796 22418 26852 22428
rect 25900 21810 26180 21812
rect 25900 21758 26126 21810
rect 26178 21758 26180 21810
rect 25900 21756 26180 21758
rect 25900 20802 25956 21756
rect 26124 21746 26180 21756
rect 25900 20750 25902 20802
rect 25954 20750 25956 20802
rect 25900 20132 25956 20750
rect 26684 20802 26740 20814
rect 26684 20750 26686 20802
rect 26738 20750 26740 20802
rect 26124 20692 26180 20702
rect 25900 20066 25956 20076
rect 26012 20580 26068 20590
rect 25900 19460 25956 19470
rect 26012 19460 26068 20524
rect 25900 19458 26068 19460
rect 25900 19406 25902 19458
rect 25954 19406 26068 19458
rect 25900 19404 26068 19406
rect 25900 19394 25956 19404
rect 26124 19346 26180 20636
rect 26460 20692 26516 20702
rect 26460 20242 26516 20636
rect 26684 20692 26740 20750
rect 26684 20626 26740 20636
rect 26460 20190 26462 20242
rect 26514 20190 26516 20242
rect 26460 20178 26516 20190
rect 26684 20020 26740 20030
rect 26684 19926 26740 19964
rect 26572 19908 26628 19918
rect 26124 19294 26126 19346
rect 26178 19294 26180 19346
rect 26124 19282 26180 19294
rect 26460 19906 26628 19908
rect 26460 19854 26574 19906
rect 26626 19854 26628 19906
rect 26460 19852 26628 19854
rect 26460 18900 26516 19852
rect 26572 19842 26628 19852
rect 26572 19684 26628 19694
rect 26572 19348 26628 19628
rect 26572 19254 26628 19292
rect 26460 18834 26516 18844
rect 26572 18788 26628 18798
rect 25676 18732 26068 18788
rect 25788 18562 25844 18574
rect 25788 18510 25790 18562
rect 25842 18510 25844 18562
rect 25788 18452 25844 18510
rect 25452 18396 25844 18452
rect 25900 18562 25956 18574
rect 25900 18510 25902 18562
rect 25954 18510 25956 18562
rect 25340 17554 25396 17566
rect 25340 17502 25342 17554
rect 25394 17502 25396 17554
rect 25004 13132 25172 13188
rect 25228 17442 25284 17454
rect 25228 17390 25230 17442
rect 25282 17390 25284 17442
rect 24668 12964 24724 12974
rect 24668 12870 24724 12908
rect 24892 12964 24948 12974
rect 24892 12402 24948 12908
rect 24892 12350 24894 12402
rect 24946 12350 24948 12402
rect 24892 12338 24948 12350
rect 23772 11778 23828 11788
rect 23436 11666 23492 11676
rect 23996 11396 24052 11406
rect 23996 11302 24052 11340
rect 25004 11394 25060 13132
rect 25116 12964 25172 12974
rect 25116 12870 25172 12908
rect 25228 11620 25284 17390
rect 25340 17108 25396 17502
rect 25340 17042 25396 17052
rect 25452 16660 25508 18396
rect 25788 18228 25844 18238
rect 25788 18134 25844 18172
rect 25900 18116 25956 18510
rect 25900 17668 25956 18060
rect 25900 17602 25956 17612
rect 25564 17556 25620 17566
rect 25564 17554 25844 17556
rect 25564 17502 25566 17554
rect 25618 17502 25844 17554
rect 25564 17500 25844 17502
rect 25564 17490 25620 17500
rect 25452 16594 25508 16604
rect 25564 17220 25620 17230
rect 25564 16210 25620 17164
rect 25788 17106 25844 17500
rect 25788 17054 25790 17106
rect 25842 17054 25844 17106
rect 25788 17042 25844 17054
rect 25900 17108 25956 17118
rect 25900 17014 25956 17052
rect 25788 16884 25844 16894
rect 25676 16660 25732 16670
rect 25676 16566 25732 16604
rect 25564 16158 25566 16210
rect 25618 16158 25620 16210
rect 25564 16146 25620 16158
rect 25564 15316 25620 15326
rect 25788 15316 25844 16828
rect 25564 15314 25844 15316
rect 25564 15262 25566 15314
rect 25618 15262 25844 15314
rect 25564 15260 25844 15262
rect 25564 15250 25620 15260
rect 25788 15148 25844 15260
rect 25676 15092 25732 15102
rect 25788 15092 25956 15148
rect 25564 14980 25620 14990
rect 25340 14306 25396 14318
rect 25340 14254 25342 14306
rect 25394 14254 25396 14306
rect 25340 14084 25396 14254
rect 25564 14308 25620 14924
rect 25676 14642 25732 15036
rect 25676 14590 25678 14642
rect 25730 14590 25732 14642
rect 25676 14578 25732 14590
rect 25788 14532 25844 14542
rect 25788 14438 25844 14476
rect 25900 14308 25956 15092
rect 25564 14306 25732 14308
rect 25564 14254 25566 14306
rect 25618 14254 25732 14306
rect 25564 14252 25732 14254
rect 25564 14242 25620 14252
rect 25340 14018 25396 14028
rect 25564 14084 25620 14094
rect 25452 13972 25508 13982
rect 25452 12850 25508 13916
rect 25452 12798 25454 12850
rect 25506 12798 25508 12850
rect 25452 12786 25508 12798
rect 25564 13746 25620 14028
rect 25564 13694 25566 13746
rect 25618 13694 25620 13746
rect 25228 11564 25396 11620
rect 25004 11342 25006 11394
rect 25058 11342 25060 11394
rect 24108 11170 24164 11182
rect 24108 11118 24110 11170
rect 24162 11118 24164 11170
rect 24108 10836 24164 11118
rect 24108 10770 24164 10780
rect 24332 11170 24388 11182
rect 24332 11118 24334 11170
rect 24386 11118 24388 11170
rect 23996 10724 24052 10734
rect 23996 10630 24052 10668
rect 24332 10610 24388 11118
rect 24892 10836 24948 10846
rect 25004 10836 25060 11342
rect 24892 10834 25060 10836
rect 24892 10782 24894 10834
rect 24946 10782 25060 10834
rect 24892 10780 25060 10782
rect 24892 10770 24948 10780
rect 24332 10558 24334 10610
rect 24386 10558 24388 10610
rect 24332 10546 24388 10558
rect 25004 10612 25060 10780
rect 25004 10546 25060 10556
rect 25228 11394 25284 11406
rect 25228 11342 25230 11394
rect 25282 11342 25284 11394
rect 25228 10276 25284 11342
rect 25228 10210 25284 10220
rect 25340 10052 25396 11564
rect 25564 10388 25620 13694
rect 25676 13636 25732 14252
rect 25676 13570 25732 13580
rect 25788 14252 25956 14308
rect 25676 13412 25732 13422
rect 25676 11618 25732 13356
rect 25676 11566 25678 11618
rect 25730 11566 25732 11618
rect 25676 11554 25732 11566
rect 25564 10322 25620 10332
rect 25676 10498 25732 10510
rect 25676 10446 25678 10498
rect 25730 10446 25732 10498
rect 25004 9996 25396 10052
rect 25452 10164 25508 10174
rect 24108 9828 24164 9838
rect 24108 9734 24164 9772
rect 23772 9602 23828 9614
rect 23772 9550 23774 9602
rect 23826 9550 23828 9602
rect 23772 9492 23828 9550
rect 23772 9426 23828 9436
rect 24892 9602 24948 9614
rect 24892 9550 24894 9602
rect 24946 9550 24948 9602
rect 24892 9492 24948 9550
rect 24892 9426 24948 9436
rect 25004 9266 25060 9996
rect 25228 9828 25284 9838
rect 25452 9828 25508 10108
rect 25284 9772 25508 9828
rect 25564 9828 25620 9838
rect 25676 9828 25732 10446
rect 25788 10276 25844 14252
rect 26012 14196 26068 18732
rect 26460 18564 26516 18574
rect 26460 18470 26516 18508
rect 26124 18452 26180 18462
rect 26124 17892 26180 18396
rect 26124 17778 26180 17836
rect 26124 17726 26126 17778
rect 26178 17726 26180 17778
rect 26124 17332 26180 17726
rect 26124 17266 26180 17276
rect 26460 17108 26516 17118
rect 26572 17108 26628 18732
rect 26908 18676 26964 18686
rect 27020 18676 27076 23884
rect 27468 23826 27524 23838
rect 27468 23774 27470 23826
rect 27522 23774 27524 23826
rect 27132 23714 27188 23726
rect 27132 23662 27134 23714
rect 27186 23662 27188 23714
rect 27132 23604 27188 23662
rect 27132 23538 27188 23548
rect 27132 23380 27188 23390
rect 27132 22372 27188 23324
rect 27356 23268 27412 23278
rect 27468 23268 27524 23774
rect 28028 23380 28084 25454
rect 28028 23314 28084 23324
rect 28140 25284 28196 25294
rect 27356 23266 27524 23268
rect 27356 23214 27358 23266
rect 27410 23214 27524 23266
rect 27356 23212 27524 23214
rect 27356 23202 27412 23212
rect 27244 23156 27300 23166
rect 27244 23062 27300 23100
rect 27468 22482 27524 23212
rect 27580 23156 27636 23166
rect 28140 23156 28196 25228
rect 28588 25284 28644 25294
rect 28588 25190 28644 25228
rect 27580 23154 27860 23156
rect 27580 23102 27582 23154
rect 27634 23102 27860 23154
rect 27580 23100 27860 23102
rect 27580 23090 27636 23100
rect 27468 22430 27470 22482
rect 27522 22430 27524 22482
rect 27468 22418 27524 22430
rect 27580 22482 27636 22494
rect 27580 22430 27582 22482
rect 27634 22430 27636 22482
rect 27244 22372 27300 22382
rect 27132 22370 27300 22372
rect 27132 22318 27246 22370
rect 27298 22318 27300 22370
rect 27132 22316 27300 22318
rect 27580 22372 27636 22430
rect 27692 22372 27748 22382
rect 27580 22370 27748 22372
rect 27580 22318 27694 22370
rect 27746 22318 27748 22370
rect 27580 22316 27748 22318
rect 27132 20690 27188 22316
rect 27244 22306 27300 22316
rect 27692 22306 27748 22316
rect 27132 20638 27134 20690
rect 27186 20638 27188 20690
rect 27132 20244 27188 20638
rect 27244 20580 27300 20590
rect 27244 20486 27300 20524
rect 27356 20578 27412 20590
rect 27356 20526 27358 20578
rect 27410 20526 27412 20578
rect 27132 20178 27188 20188
rect 27132 20020 27188 20030
rect 27356 20020 27412 20526
rect 27132 20018 27412 20020
rect 27132 19966 27134 20018
rect 27186 19966 27412 20018
rect 27132 19964 27412 19966
rect 27468 20578 27524 20590
rect 27468 20526 27470 20578
rect 27522 20526 27524 20578
rect 27132 19954 27188 19964
rect 27468 19908 27524 20526
rect 27692 19908 27748 19918
rect 27468 19906 27748 19908
rect 27468 19854 27694 19906
rect 27746 19854 27748 19906
rect 27468 19852 27748 19854
rect 27692 19684 27748 19852
rect 27692 19618 27748 19628
rect 27244 19010 27300 19022
rect 27244 18958 27246 19010
rect 27298 18958 27300 19010
rect 27244 18676 27300 18958
rect 27804 18788 27860 23100
rect 27916 23100 28196 23156
rect 28476 24500 28532 24510
rect 28476 23154 28532 24444
rect 28924 23716 28980 23726
rect 28924 23622 28980 23660
rect 28476 23102 28478 23154
rect 28530 23102 28532 23154
rect 27916 22370 27972 23100
rect 28476 23090 28532 23102
rect 27916 22318 27918 22370
rect 27970 22318 27972 22370
rect 27916 22260 27972 22318
rect 28140 22930 28196 22942
rect 28140 22878 28142 22930
rect 28194 22878 28196 22930
rect 28028 22260 28084 22270
rect 27916 22258 28084 22260
rect 27916 22206 28030 22258
rect 28082 22206 28084 22258
rect 27916 22204 28084 22206
rect 28028 22194 28084 22204
rect 28140 21700 28196 22878
rect 28924 22372 28980 22382
rect 28924 22278 28980 22316
rect 28140 21644 28532 21700
rect 28252 21476 28308 21486
rect 28028 21474 28308 21476
rect 28028 21422 28254 21474
rect 28306 21422 28308 21474
rect 28028 21420 28308 21422
rect 28028 20690 28084 21420
rect 28252 21410 28308 21420
rect 28476 20802 28532 21644
rect 28700 21476 28756 21486
rect 28476 20750 28478 20802
rect 28530 20750 28532 20802
rect 28476 20738 28532 20750
rect 28588 21474 28756 21476
rect 28588 21422 28702 21474
rect 28754 21422 28756 21474
rect 28588 21420 28756 21422
rect 28028 20638 28030 20690
rect 28082 20638 28084 20690
rect 27916 20580 27972 20590
rect 27916 20486 27972 20524
rect 28028 19796 28084 20638
rect 28252 20580 28308 20590
rect 28588 20580 28644 21420
rect 28700 21410 28756 21420
rect 28252 20578 28644 20580
rect 28252 20526 28254 20578
rect 28306 20526 28644 20578
rect 28252 20524 28644 20526
rect 28700 20690 28756 20702
rect 28700 20638 28702 20690
rect 28754 20638 28756 20690
rect 28252 20468 28308 20524
rect 28140 20132 28196 20142
rect 28140 20038 28196 20076
rect 28028 19730 28084 19740
rect 27804 18732 28084 18788
rect 27020 18620 27188 18676
rect 26908 18564 26964 18620
rect 26908 18508 27076 18564
rect 26796 18450 26852 18462
rect 26796 18398 26798 18450
rect 26850 18398 26852 18450
rect 26796 17668 26852 18398
rect 27020 18450 27076 18508
rect 27020 18398 27022 18450
rect 27074 18398 27076 18450
rect 27020 18386 27076 18398
rect 26908 18338 26964 18350
rect 26908 18286 26910 18338
rect 26962 18286 26964 18338
rect 26908 17668 26964 18286
rect 26908 17612 27076 17668
rect 26796 17602 26852 17612
rect 26684 17444 26740 17454
rect 26684 17350 26740 17388
rect 26796 17442 26852 17454
rect 26796 17390 26798 17442
rect 26850 17390 26852 17442
rect 26516 17052 26628 17108
rect 26236 16996 26292 17006
rect 26236 15876 26292 16940
rect 26348 16212 26404 16222
rect 26460 16212 26516 17052
rect 26348 16210 26516 16212
rect 26348 16158 26350 16210
rect 26402 16158 26516 16210
rect 26348 16156 26516 16158
rect 26348 16146 26404 16156
rect 26684 15876 26740 15886
rect 26236 15874 26740 15876
rect 26236 15822 26686 15874
rect 26738 15822 26740 15874
rect 26236 15820 26740 15822
rect 26236 15314 26292 15326
rect 26236 15262 26238 15314
rect 26290 15262 26292 15314
rect 26236 14980 26292 15262
rect 26236 14914 26292 14924
rect 25900 14140 26068 14196
rect 26124 14308 26180 14318
rect 25900 12964 25956 14140
rect 25900 12178 25956 12908
rect 26012 13972 26068 13982
rect 26012 12962 26068 13916
rect 26124 13970 26180 14252
rect 26124 13918 26126 13970
rect 26178 13918 26180 13970
rect 26124 13906 26180 13918
rect 26236 13972 26292 13982
rect 26236 13878 26292 13916
rect 26348 13412 26404 15820
rect 26684 15810 26740 15820
rect 26572 15428 26628 15438
rect 26796 15428 26852 17390
rect 26572 15426 26852 15428
rect 26572 15374 26574 15426
rect 26626 15374 26852 15426
rect 26572 15372 26852 15374
rect 26908 17442 26964 17454
rect 26908 17390 26910 17442
rect 26962 17390 26964 17442
rect 26908 17332 26964 17390
rect 26572 15362 26628 15372
rect 26348 13346 26404 13356
rect 26460 15202 26516 15214
rect 26460 15150 26462 15202
rect 26514 15150 26516 15202
rect 26012 12910 26014 12962
rect 26066 12910 26068 12962
rect 26012 12898 26068 12910
rect 26460 12964 26516 15150
rect 26796 14532 26852 14542
rect 26796 14438 26852 14476
rect 26684 14308 26740 14318
rect 26684 14214 26740 14252
rect 26908 14308 26964 17276
rect 27020 15148 27076 17612
rect 27132 16884 27188 18620
rect 27244 18610 27300 18620
rect 27580 18676 27636 18686
rect 27580 18582 27636 18620
rect 28028 18674 28084 18732
rect 28028 18622 28030 18674
rect 28082 18622 28084 18674
rect 27692 18564 27748 18574
rect 27692 18470 27748 18508
rect 27804 18452 27860 18462
rect 27804 18358 27860 18396
rect 28028 18340 28084 18622
rect 28028 18274 28084 18284
rect 28252 18116 28308 20412
rect 28364 20130 28420 20142
rect 28364 20078 28366 20130
rect 28418 20078 28420 20130
rect 28364 20020 28420 20078
rect 28700 20132 28756 20638
rect 29036 20244 29092 29932
rect 29260 29650 29316 31836
rect 29484 31892 29540 31902
rect 29484 31798 29540 31836
rect 29596 30324 29652 32844
rect 29260 29598 29262 29650
rect 29314 29598 29316 29650
rect 29260 29586 29316 29598
rect 29484 30268 29652 30324
rect 29372 27970 29428 27982
rect 29372 27918 29374 27970
rect 29426 27918 29428 27970
rect 29372 27860 29428 27918
rect 29372 27300 29428 27804
rect 29372 27234 29428 27244
rect 29484 26908 29540 30268
rect 29596 30098 29652 30110
rect 29596 30046 29598 30098
rect 29650 30046 29652 30098
rect 29596 29764 29652 30046
rect 29708 30100 29764 30110
rect 29708 30006 29764 30044
rect 29932 29988 29988 29998
rect 29596 29092 29652 29708
rect 29596 29026 29652 29036
rect 29820 29986 29988 29988
rect 29820 29934 29934 29986
rect 29986 29934 29988 29986
rect 29820 29932 29988 29934
rect 29820 29204 29876 29932
rect 29932 29922 29988 29932
rect 29820 28754 29876 29148
rect 29820 28702 29822 28754
rect 29874 28702 29876 28754
rect 29820 28690 29876 28702
rect 30044 29652 30100 29662
rect 30044 28644 30100 29596
rect 30044 28578 30100 28588
rect 29708 28084 29764 28094
rect 30156 28084 30212 33068
rect 30716 33012 30772 33068
rect 30828 33058 30884 33068
rect 30940 33122 30996 33134
rect 30940 33070 30942 33122
rect 30994 33070 30996 33122
rect 30716 32946 30772 32956
rect 30380 32676 30436 32686
rect 30380 32582 30436 32620
rect 30940 32676 30996 33070
rect 30940 32610 30996 32620
rect 30380 32340 30436 32350
rect 30268 31668 30324 31678
rect 30268 30210 30324 31612
rect 30268 30158 30270 30210
rect 30322 30158 30324 30210
rect 30268 30100 30324 30158
rect 30268 28980 30324 30044
rect 30380 31108 30436 32284
rect 30492 31108 30548 31118
rect 30380 31052 30492 31108
rect 30380 28980 30436 31052
rect 30492 30976 30548 31052
rect 30716 30100 30772 30110
rect 30716 29652 30772 30044
rect 30828 29986 30884 29998
rect 30828 29934 30830 29986
rect 30882 29934 30884 29986
rect 30828 29764 30884 29934
rect 30828 29698 30884 29708
rect 30716 29520 30772 29596
rect 31164 29540 31220 33740
rect 31276 31218 31332 34300
rect 31388 33012 31444 33022
rect 31388 31890 31444 32956
rect 31388 31838 31390 31890
rect 31442 31838 31444 31890
rect 31388 31826 31444 31838
rect 31276 31166 31278 31218
rect 31330 31166 31332 31218
rect 31276 31154 31332 31166
rect 31276 29988 31332 29998
rect 31276 29894 31332 29932
rect 30828 29484 31220 29540
rect 30828 29428 30884 29484
rect 30716 29372 30884 29428
rect 30604 29314 30660 29326
rect 30604 29262 30606 29314
rect 30658 29262 30660 29314
rect 30492 29204 30548 29214
rect 30492 29110 30548 29148
rect 30380 28924 30548 28980
rect 30268 28914 30324 28924
rect 29708 28082 30212 28084
rect 29708 28030 29710 28082
rect 29762 28030 30212 28082
rect 29708 28028 30212 28030
rect 29708 28018 29764 28028
rect 30044 27186 30100 28028
rect 30156 27748 30212 28028
rect 30268 28530 30324 28542
rect 30268 28478 30270 28530
rect 30322 28478 30324 28530
rect 30268 27972 30324 28478
rect 30268 27906 30324 27916
rect 30268 27748 30324 27758
rect 30156 27746 30324 27748
rect 30156 27694 30270 27746
rect 30322 27694 30324 27746
rect 30156 27692 30324 27694
rect 30268 27682 30324 27692
rect 30044 27134 30046 27186
rect 30098 27134 30100 27186
rect 30044 27122 30100 27134
rect 30380 27412 30436 27422
rect 30380 27186 30436 27356
rect 30492 27300 30548 28924
rect 30604 28756 30660 29262
rect 30604 28690 30660 28700
rect 30492 27234 30548 27244
rect 30604 28532 30660 28542
rect 30380 27134 30382 27186
rect 30434 27134 30436 27186
rect 29484 26852 29652 26908
rect 29148 23268 29204 23278
rect 29148 23174 29204 23212
rect 29260 23154 29316 23166
rect 29260 23102 29262 23154
rect 29314 23102 29316 23154
rect 29260 22372 29316 23102
rect 29596 22708 29652 26852
rect 29932 26292 29988 26302
rect 29932 26198 29988 26236
rect 30044 25282 30100 25294
rect 30044 25230 30046 25282
rect 30098 25230 30100 25282
rect 29708 25172 29764 25182
rect 29708 24946 29764 25116
rect 29708 24894 29710 24946
rect 29762 24894 29764 24946
rect 29708 24882 29764 24894
rect 29820 24948 29876 24958
rect 29820 24834 29876 24892
rect 30044 24948 30100 25230
rect 30044 24882 30100 24892
rect 30268 25172 30324 25182
rect 30268 24946 30324 25116
rect 30268 24894 30270 24946
rect 30322 24894 30324 24946
rect 30268 24882 30324 24894
rect 29820 24782 29822 24834
rect 29874 24782 29876 24834
rect 29708 24500 29764 24510
rect 29708 24406 29764 24444
rect 29820 23940 29876 24782
rect 29932 23940 29988 23950
rect 29820 23938 29988 23940
rect 29820 23886 29934 23938
rect 29986 23886 29988 23938
rect 29820 23884 29988 23886
rect 29932 23874 29988 23884
rect 30044 23716 30100 23726
rect 30044 23622 30100 23660
rect 30268 23714 30324 23726
rect 30268 23662 30270 23714
rect 30322 23662 30324 23714
rect 30268 23380 30324 23662
rect 30380 23604 30436 27134
rect 30604 27076 30660 28476
rect 30492 27020 30660 27076
rect 30492 23716 30548 27020
rect 30604 26908 30660 26918
rect 30604 26290 30660 26852
rect 30604 26238 30606 26290
rect 30658 26238 30660 26290
rect 30604 26226 30660 26238
rect 30604 24948 30660 24958
rect 30604 24050 30660 24892
rect 30604 23998 30606 24050
rect 30658 23998 30660 24050
rect 30604 23986 30660 23998
rect 30492 23660 30660 23716
rect 30380 23548 30548 23604
rect 30380 23380 30436 23390
rect 30268 23378 30436 23380
rect 30268 23326 30382 23378
rect 30434 23326 30436 23378
rect 30268 23324 30436 23326
rect 30380 23314 30436 23324
rect 29596 22642 29652 22652
rect 29820 23268 29876 23278
rect 29820 23156 29876 23212
rect 29932 23156 29988 23166
rect 29820 23154 29988 23156
rect 29820 23102 29934 23154
rect 29986 23102 29988 23154
rect 29820 23100 29988 23102
rect 29260 22306 29316 22316
rect 29708 22372 29764 22382
rect 29708 22278 29764 22316
rect 29484 22148 29540 22158
rect 28364 19954 28420 19964
rect 28476 20018 28532 20030
rect 28476 19966 28478 20018
rect 28530 19966 28532 20018
rect 28476 19012 28532 19966
rect 28700 19908 28756 20076
rect 28700 19842 28756 19852
rect 28812 20242 29092 20244
rect 28812 20190 29038 20242
rect 29090 20190 29092 20242
rect 28812 20188 29092 20190
rect 28700 19012 28756 19022
rect 28476 18956 28700 19012
rect 28476 18788 28532 18956
rect 28700 18918 28756 18956
rect 28476 18722 28532 18732
rect 28812 18564 28868 20188
rect 29036 20178 29092 20188
rect 29148 21698 29204 21710
rect 29148 21646 29150 21698
rect 29202 21646 29204 21698
rect 29148 20020 29204 21646
rect 29484 21698 29540 22092
rect 29820 21924 29876 23100
rect 29932 23090 29988 23100
rect 30156 23154 30212 23166
rect 30156 23102 30158 23154
rect 30210 23102 30212 23154
rect 30044 23042 30100 23054
rect 30044 22990 30046 23042
rect 30098 22990 30100 23042
rect 29932 22148 29988 22158
rect 29932 22054 29988 22092
rect 29820 21858 29876 21868
rect 29484 21646 29486 21698
rect 29538 21646 29540 21698
rect 29484 21634 29540 21646
rect 30044 21700 30100 22990
rect 30156 22148 30212 23102
rect 30156 22082 30212 22092
rect 30380 22596 30436 22606
rect 30044 21634 30100 21644
rect 30156 21924 30212 21934
rect 30044 21476 30100 21486
rect 30156 21476 30212 21868
rect 30044 21474 30212 21476
rect 30044 21422 30046 21474
rect 30098 21422 30212 21474
rect 30044 21420 30212 21422
rect 30044 21410 30100 21420
rect 29932 20804 29988 20814
rect 29932 20710 29988 20748
rect 30156 20578 30212 20590
rect 30156 20526 30158 20578
rect 30210 20526 30212 20578
rect 30044 20356 30100 20366
rect 29932 20132 29988 20142
rect 29932 20038 29988 20076
rect 29372 20020 29428 20030
rect 29148 20018 29428 20020
rect 29148 19966 29374 20018
rect 29426 19966 29428 20018
rect 29148 19964 29428 19966
rect 29372 19012 29428 19964
rect 29820 19908 29876 19918
rect 29596 19012 29652 19022
rect 29372 19010 29652 19012
rect 29372 18958 29598 19010
rect 29650 18958 29652 19010
rect 29372 18956 29652 18958
rect 27804 18060 28308 18116
rect 28588 18508 28868 18564
rect 27580 17780 27636 17790
rect 27244 17666 27300 17678
rect 27244 17614 27246 17666
rect 27298 17614 27300 17666
rect 27244 17106 27300 17614
rect 27244 17054 27246 17106
rect 27298 17054 27300 17106
rect 27244 17042 27300 17054
rect 27468 17556 27524 17566
rect 27468 16994 27524 17500
rect 27468 16942 27470 16994
rect 27522 16942 27524 16994
rect 27132 16828 27300 16884
rect 27132 15874 27188 15886
rect 27132 15822 27134 15874
rect 27186 15822 27188 15874
rect 27132 15652 27188 15822
rect 27132 15428 27188 15596
rect 27132 15362 27188 15372
rect 27020 15092 27188 15148
rect 26908 14306 27076 14308
rect 26908 14254 26910 14306
rect 26962 14254 27076 14306
rect 26908 14252 27076 14254
rect 26908 14242 26964 14252
rect 27020 13748 27076 14252
rect 27020 13682 27076 13692
rect 26460 12908 26740 12964
rect 26348 12740 26404 12750
rect 25900 12126 25902 12178
rect 25954 12126 25956 12178
rect 25900 12114 25956 12126
rect 26236 12738 26404 12740
rect 26236 12686 26350 12738
rect 26402 12686 26404 12738
rect 26236 12684 26404 12686
rect 26124 11956 26180 11966
rect 26236 11956 26292 12684
rect 26348 12674 26404 12684
rect 26460 12738 26516 12750
rect 26460 12686 26462 12738
rect 26514 12686 26516 12738
rect 26348 12516 26404 12526
rect 26348 12178 26404 12460
rect 26348 12126 26350 12178
rect 26402 12126 26404 12178
rect 26348 12114 26404 12126
rect 26124 11954 26292 11956
rect 26124 11902 26126 11954
rect 26178 11902 26292 11954
rect 26124 11900 26292 11902
rect 26124 11620 26180 11900
rect 26124 11554 26180 11564
rect 26348 11394 26404 11406
rect 26348 11342 26350 11394
rect 26402 11342 26404 11394
rect 25900 10612 25956 10622
rect 25900 10518 25956 10556
rect 26124 10610 26180 10622
rect 26124 10558 26126 10610
rect 26178 10558 26180 10610
rect 25788 10210 25844 10220
rect 26124 10052 26180 10558
rect 26124 9986 26180 9996
rect 26236 10388 26292 10398
rect 26012 9828 26068 9838
rect 25676 9772 25844 9828
rect 25228 9696 25284 9772
rect 25004 9214 25006 9266
rect 25058 9214 25060 9266
rect 24444 8484 24500 8494
rect 23548 8372 23604 8382
rect 23548 8278 23604 8316
rect 24220 8372 24276 8382
rect 23772 8148 23828 8158
rect 23660 8146 23828 8148
rect 23660 8094 23774 8146
rect 23826 8094 23828 8146
rect 23660 8092 23828 8094
rect 23436 7476 23492 7486
rect 23436 7382 23492 7420
rect 23660 7476 23716 8092
rect 23772 8082 23828 8092
rect 23884 8148 23940 8158
rect 23660 7252 23716 7420
rect 23436 7196 23716 7252
rect 23884 7474 23940 8092
rect 23884 7422 23886 7474
rect 23938 7422 23940 7474
rect 23436 6690 23492 7196
rect 23436 6638 23438 6690
rect 23490 6638 23492 6690
rect 23436 6626 23492 6638
rect 23884 6692 23940 7422
rect 23996 6692 24052 6702
rect 23884 6690 24052 6692
rect 23884 6638 23998 6690
rect 24050 6638 24052 6690
rect 23884 6636 24052 6638
rect 23996 6626 24052 6636
rect 24220 6690 24276 8316
rect 24444 8370 24500 8428
rect 24444 8318 24446 8370
rect 24498 8318 24500 8370
rect 24444 8306 24500 8318
rect 24892 8372 24948 8382
rect 24892 7586 24948 8316
rect 25004 8260 25060 9214
rect 25004 8166 25060 8204
rect 25116 9604 25172 9614
rect 25116 8484 25172 9548
rect 25564 8428 25620 9772
rect 25788 9714 25844 9772
rect 26012 9734 26068 9772
rect 25788 9662 25790 9714
rect 25842 9662 25844 9714
rect 25676 9604 25732 9614
rect 25788 9604 25844 9662
rect 25788 9548 26068 9604
rect 25676 9266 25732 9548
rect 25676 9214 25678 9266
rect 25730 9214 25732 9266
rect 25676 9202 25732 9214
rect 25900 9042 25956 9054
rect 25900 8990 25902 9042
rect 25954 8990 25956 9042
rect 25788 8930 25844 8942
rect 25788 8878 25790 8930
rect 25842 8878 25844 8930
rect 25116 8258 25172 8428
rect 25340 8372 25396 8382
rect 25340 8278 25396 8316
rect 25452 8372 25620 8428
rect 25676 8482 25732 8494
rect 25676 8430 25678 8482
rect 25730 8430 25732 8482
rect 25116 8206 25118 8258
rect 25170 8206 25172 8258
rect 25116 8194 25172 8206
rect 25452 7700 25508 8372
rect 25564 8260 25620 8270
rect 25676 8260 25732 8430
rect 25564 8258 25732 8260
rect 25564 8206 25566 8258
rect 25618 8206 25732 8258
rect 25564 8204 25732 8206
rect 25564 8194 25620 8204
rect 25676 8036 25732 8204
rect 25676 7970 25732 7980
rect 25452 7644 25620 7700
rect 24892 7534 24894 7586
rect 24946 7534 24948 7586
rect 24892 7522 24948 7534
rect 24556 7476 24612 7514
rect 24556 7410 24612 7420
rect 24668 7364 24724 7374
rect 24556 7252 24612 7262
rect 24556 7158 24612 7196
rect 24220 6638 24222 6690
rect 24274 6638 24276 6690
rect 24220 6626 24276 6638
rect 24668 6690 24724 7308
rect 24668 6638 24670 6690
rect 24722 6638 24724 6690
rect 24668 6626 24724 6638
rect 24108 6466 24164 6478
rect 24108 6414 24110 6466
rect 24162 6414 24164 6466
rect 24108 6020 24164 6414
rect 24556 6244 24612 6254
rect 24556 6130 24612 6188
rect 24556 6078 24558 6130
rect 24610 6078 24612 6130
rect 24332 6020 24388 6030
rect 24108 6018 24388 6020
rect 24108 5966 24334 6018
rect 24386 5966 24388 6018
rect 24108 5964 24388 5966
rect 23324 5506 23380 5516
rect 24108 5124 24164 5134
rect 24108 5030 24164 5068
rect 24220 5122 24276 5964
rect 24332 5954 24388 5964
rect 24220 5070 24222 5122
rect 24274 5070 24276 5122
rect 24220 5058 24276 5070
rect 24556 5124 24612 6078
rect 24668 5684 24724 5694
rect 24668 5682 24948 5684
rect 24668 5630 24670 5682
rect 24722 5630 24948 5682
rect 24668 5628 24948 5630
rect 24668 5618 24724 5628
rect 24556 5058 24612 5068
rect 24892 5122 24948 5628
rect 24892 5070 24894 5122
rect 24946 5070 24948 5122
rect 24892 5058 24948 5070
rect 23100 4946 23156 4956
rect 23772 5012 23828 5022
rect 23772 4918 23828 4956
rect 23996 5012 24052 5022
rect 23996 4918 24052 4956
rect 25116 5010 25172 5022
rect 25116 4958 25118 5010
rect 25170 4958 25172 5010
rect 22540 4900 22596 4910
rect 22540 4806 22596 4844
rect 23884 4898 23940 4910
rect 23884 4846 23886 4898
rect 23938 4846 23940 4898
rect 23884 4788 23940 4846
rect 25116 4900 25172 4958
rect 25452 5012 25508 5022
rect 25452 4918 25508 4956
rect 25116 4834 25172 4844
rect 25340 4900 25396 4910
rect 25340 4806 25396 4844
rect 23884 4722 23940 4732
rect 23660 4452 23716 4462
rect 22428 4286 22430 4338
rect 22482 4286 22484 4338
rect 22428 4274 22484 4286
rect 23100 4340 23156 4350
rect 23100 4246 23156 4284
rect 19292 3666 19460 3668
rect 19292 3614 19294 3666
rect 19346 3614 19460 3666
rect 19292 3612 19460 3614
rect 12236 3554 12740 3556
rect 12236 3502 12238 3554
rect 12290 3502 12740 3554
rect 12236 3500 12740 3502
rect 18732 3556 18788 3566
rect 19292 3556 19348 3612
rect 18732 3554 19348 3556
rect 18732 3502 18734 3554
rect 18786 3502 19348 3554
rect 18732 3500 19348 3502
rect 23660 3554 23716 4396
rect 23660 3502 23662 3554
rect 23714 3502 23716 3554
rect 12236 3490 12292 3500
rect 18732 3490 18788 3500
rect 23660 3490 23716 3502
rect 23884 4226 23940 4238
rect 23884 4174 23886 4226
rect 23938 4174 23940 4226
rect 3164 2594 3220 2604
rect 5068 3444 5124 3454
rect 5068 2212 5124 3388
rect 5852 3444 5908 3454
rect 11116 3444 11172 3454
rect 5852 3350 5908 3388
rect 10780 3442 11172 3444
rect 10780 3390 11118 3442
rect 11170 3390 11172 3442
rect 10780 3388 11172 3390
rect 5068 2156 5460 2212
rect 1932 1810 1988 1820
rect 5404 800 5460 2156
rect 10780 800 10836 3388
rect 11116 3378 11172 3388
rect 16828 3444 16884 3454
rect 16828 800 16884 3388
rect 17612 3444 17668 3454
rect 22540 3442 22596 3454
rect 22540 3390 22542 3442
rect 22594 3390 22596 3442
rect 22540 3388 22596 3390
rect 17612 3350 17668 3388
rect 22204 3332 22596 3388
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 22204 800 22260 3332
rect 23884 2772 23940 4174
rect 25564 4228 25620 7644
rect 25676 7476 25732 7486
rect 25676 7382 25732 7420
rect 25788 7364 25844 8878
rect 25900 8482 25956 8990
rect 25900 8430 25902 8482
rect 25954 8430 25956 8482
rect 25900 8418 25956 8430
rect 25900 8260 25956 8270
rect 25900 8166 25956 8204
rect 26012 7476 26068 9548
rect 26236 9602 26292 10332
rect 26348 10050 26404 11342
rect 26460 10724 26516 12686
rect 26572 12738 26628 12750
rect 26572 12686 26574 12738
rect 26626 12686 26628 12738
rect 26572 12516 26628 12686
rect 26572 12450 26628 12460
rect 26684 11396 26740 12908
rect 27132 12292 27188 15092
rect 27244 12516 27300 16828
rect 27468 15540 27524 16942
rect 27580 17444 27636 17724
rect 27580 16994 27636 17388
rect 27580 16942 27582 16994
rect 27634 16942 27636 16994
rect 27580 16930 27636 16942
rect 27468 15474 27524 15484
rect 27356 15202 27412 15214
rect 27356 15150 27358 15202
rect 27410 15150 27412 15202
rect 27356 15148 27412 15150
rect 27804 15148 27860 18060
rect 28028 17780 28084 17790
rect 28028 17778 28196 17780
rect 28028 17726 28030 17778
rect 28082 17726 28196 17778
rect 28028 17724 28196 17726
rect 28028 17714 28084 17724
rect 28028 17332 28084 17342
rect 28028 15986 28084 17276
rect 28028 15934 28030 15986
rect 28082 15934 28084 15986
rect 28028 15922 28084 15934
rect 27916 15540 27972 15550
rect 27916 15446 27972 15484
rect 28140 15428 28196 17724
rect 28252 17556 28308 17566
rect 28252 17462 28308 17500
rect 28476 17556 28532 17566
rect 28476 17106 28532 17500
rect 28476 17054 28478 17106
rect 28530 17054 28532 17106
rect 28476 17042 28532 17054
rect 28588 17554 28644 18508
rect 29260 18452 29316 18462
rect 29260 18358 29316 18396
rect 28812 18340 28868 18350
rect 28868 18284 29092 18340
rect 28812 18246 28868 18284
rect 28588 17502 28590 17554
rect 28642 17502 28644 17554
rect 28588 17108 28644 17502
rect 28812 17444 28868 17454
rect 28700 17108 28756 17118
rect 28588 17106 28756 17108
rect 28588 17054 28702 17106
rect 28754 17054 28756 17106
rect 28588 17052 28756 17054
rect 28812 17108 28868 17388
rect 28924 17108 28980 17118
rect 28812 17106 28980 17108
rect 28812 17054 28926 17106
rect 28978 17054 28980 17106
rect 28812 17052 28980 17054
rect 28700 16884 28756 17052
rect 28924 17042 28980 17052
rect 28700 16322 28756 16828
rect 28700 16270 28702 16322
rect 28754 16270 28756 16322
rect 28700 16258 28756 16270
rect 28812 16770 28868 16782
rect 28812 16718 28814 16770
rect 28866 16718 28868 16770
rect 28364 15988 28420 15998
rect 28812 15988 28868 16718
rect 28924 16322 28980 16334
rect 28924 16270 28926 16322
rect 28978 16270 28980 16322
rect 28924 16210 28980 16270
rect 28924 16158 28926 16210
rect 28978 16158 28980 16210
rect 28924 16146 28980 16158
rect 28364 15894 28420 15932
rect 28588 15932 28868 15988
rect 28476 15652 28532 15662
rect 28252 15540 28308 15550
rect 28252 15446 28308 15484
rect 28028 15372 28196 15428
rect 28028 15204 28084 15372
rect 27356 15092 27524 15148
rect 27356 14532 27412 14542
rect 27356 14438 27412 14476
rect 27468 14308 27524 15092
rect 27468 14242 27524 14252
rect 27692 15092 27860 15148
rect 27916 15148 28084 15204
rect 28364 15316 28420 15326
rect 27244 12460 27524 12516
rect 27244 12292 27300 12302
rect 27132 12290 27300 12292
rect 27132 12238 27246 12290
rect 27298 12238 27300 12290
rect 27132 12236 27300 12238
rect 27244 12226 27300 12236
rect 27356 12066 27412 12078
rect 27356 12014 27358 12066
rect 27410 12014 27412 12066
rect 26460 10658 26516 10668
rect 26572 11340 26740 11396
rect 26796 11954 26852 11966
rect 26796 11902 26798 11954
rect 26850 11902 26852 11954
rect 26348 9998 26350 10050
rect 26402 9998 26404 10050
rect 26348 9986 26404 9998
rect 26236 9550 26238 9602
rect 26290 9550 26292 9602
rect 26236 9538 26292 9550
rect 26460 9828 26516 9838
rect 26124 9042 26180 9054
rect 26124 8990 26126 9042
rect 26178 8990 26180 9042
rect 26124 8260 26180 8990
rect 26460 8260 26516 9772
rect 26572 9156 26628 11340
rect 26684 11170 26740 11182
rect 26684 11118 26686 11170
rect 26738 11118 26740 11170
rect 26684 10612 26740 11118
rect 26684 10546 26740 10556
rect 26684 10052 26740 10062
rect 26684 9602 26740 9996
rect 26796 9828 26852 11902
rect 27356 11956 27412 12014
rect 27356 11890 27412 11900
rect 27468 11060 27524 12460
rect 27132 11004 27524 11060
rect 27580 12178 27636 12190
rect 27580 12126 27582 12178
rect 27634 12126 27636 12178
rect 27580 11282 27636 12126
rect 27580 11230 27582 11282
rect 27634 11230 27636 11282
rect 27132 9828 27188 11004
rect 27580 10948 27636 11230
rect 27356 10892 27636 10948
rect 27244 10388 27300 10398
rect 27244 10294 27300 10332
rect 27132 9772 27300 9828
rect 26796 9762 26852 9772
rect 26684 9550 26686 9602
rect 26738 9550 26740 9602
rect 26684 9380 26740 9550
rect 26684 9314 26740 9324
rect 27132 9602 27188 9614
rect 27132 9550 27134 9602
rect 27186 9550 27188 9602
rect 27132 9380 27188 9550
rect 27132 9314 27188 9324
rect 26684 9156 26740 9166
rect 26572 9154 26740 9156
rect 26572 9102 26686 9154
rect 26738 9102 26740 9154
rect 26572 9100 26740 9102
rect 26684 9090 26740 9100
rect 26908 9156 26964 9194
rect 26908 9090 26964 9100
rect 26908 8930 26964 8942
rect 26908 8878 26910 8930
rect 26962 8878 26964 8930
rect 26908 8708 26964 8878
rect 26852 8652 26964 8708
rect 26852 8596 26908 8652
rect 26796 8540 26908 8596
rect 26572 8260 26628 8270
rect 26460 8258 26628 8260
rect 26460 8206 26574 8258
rect 26626 8206 26628 8258
rect 26460 8204 26628 8206
rect 26124 8194 26180 8204
rect 26572 8194 26628 8204
rect 26796 8148 26852 8540
rect 27020 8370 27076 8382
rect 27020 8318 27022 8370
rect 27074 8318 27076 8370
rect 26908 8260 26964 8270
rect 26908 8166 26964 8204
rect 26796 8082 26852 8092
rect 26572 7476 26628 7486
rect 26012 7474 26628 7476
rect 26012 7422 26574 7474
rect 26626 7422 26628 7474
rect 26012 7420 26628 7422
rect 26572 7410 26628 7420
rect 27020 7474 27076 8318
rect 27020 7422 27022 7474
rect 27074 7422 27076 7474
rect 27020 7410 27076 7422
rect 27132 8034 27188 8046
rect 27132 7982 27134 8034
rect 27186 7982 27188 8034
rect 25788 7270 25844 7308
rect 27132 6580 27188 7982
rect 27132 6020 27188 6524
rect 27244 6244 27300 9772
rect 27356 9156 27412 10892
rect 27580 10724 27636 10734
rect 27580 10610 27636 10668
rect 27580 10558 27582 10610
rect 27634 10558 27636 10610
rect 27468 9604 27524 9614
rect 27468 9266 27524 9548
rect 27468 9214 27470 9266
rect 27522 9214 27524 9266
rect 27468 9202 27524 9214
rect 27356 9090 27412 9100
rect 27580 8932 27636 10558
rect 27692 9156 27748 15092
rect 27804 14418 27860 14430
rect 27804 14366 27806 14418
rect 27858 14366 27860 14418
rect 27804 13972 27860 14366
rect 27804 13906 27860 13916
rect 27804 13748 27860 13758
rect 27804 13654 27860 13692
rect 27916 11394 27972 15148
rect 28252 14644 28308 14654
rect 28252 13188 28308 14588
rect 28364 13858 28420 15260
rect 28476 14530 28532 15596
rect 28476 14478 28478 14530
rect 28530 14478 28532 14530
rect 28476 14466 28532 14478
rect 28364 13806 28366 13858
rect 28418 13806 28420 13858
rect 28364 13794 28420 13806
rect 28476 13748 28532 13758
rect 28476 13654 28532 13692
rect 28588 13412 28644 15932
rect 28700 15540 28756 15550
rect 28700 14644 28756 15484
rect 28700 14512 28756 14588
rect 28812 15092 28868 15102
rect 28812 13748 28868 15036
rect 28812 13682 28868 13692
rect 27916 11342 27918 11394
rect 27970 11342 27972 11394
rect 27916 11330 27972 11342
rect 28140 13186 28308 13188
rect 28140 13134 28254 13186
rect 28306 13134 28308 13186
rect 28140 13132 28308 13134
rect 28028 11170 28084 11182
rect 28028 11118 28030 11170
rect 28082 11118 28084 11170
rect 27804 10498 27860 10510
rect 27804 10446 27806 10498
rect 27858 10446 27860 10498
rect 27804 9492 27860 10446
rect 28028 9940 28084 11118
rect 28028 9874 28084 9884
rect 28140 9828 28196 13132
rect 28252 13122 28308 13132
rect 28476 13356 28644 13412
rect 28700 13636 28756 13646
rect 28252 12292 28308 12302
rect 28476 12292 28532 13356
rect 28588 13076 28644 13086
rect 28588 12982 28644 13020
rect 28252 12290 28532 12292
rect 28252 12238 28254 12290
rect 28306 12238 28532 12290
rect 28252 12236 28532 12238
rect 28588 12740 28644 12750
rect 28588 12290 28644 12684
rect 28588 12238 28590 12290
rect 28642 12238 28644 12290
rect 28252 12226 28308 12236
rect 28588 12226 28644 12238
rect 28700 12178 28756 13580
rect 28924 13634 28980 13646
rect 28924 13582 28926 13634
rect 28978 13582 28980 13634
rect 28812 12852 28868 12862
rect 28812 12758 28868 12796
rect 28700 12126 28702 12178
rect 28754 12126 28756 12178
rect 28700 12114 28756 12126
rect 28364 12066 28420 12078
rect 28364 12014 28366 12066
rect 28418 12014 28420 12066
rect 28252 11396 28308 11406
rect 28364 11396 28420 12014
rect 28252 11394 28420 11396
rect 28252 11342 28254 11394
rect 28306 11342 28420 11394
rect 28252 11340 28420 11342
rect 28812 11618 28868 11630
rect 28812 11566 28814 11618
rect 28866 11566 28868 11618
rect 28812 11506 28868 11566
rect 28812 11454 28814 11506
rect 28866 11454 28868 11506
rect 28252 11330 28308 11340
rect 28364 10836 28420 10846
rect 28364 10742 28420 10780
rect 28140 9762 28196 9772
rect 28812 9938 28868 11454
rect 28924 10498 28980 13582
rect 29036 11620 29092 18284
rect 29596 18228 29652 18956
rect 29820 18676 29876 19852
rect 29820 18450 29876 18620
rect 29820 18398 29822 18450
rect 29874 18398 29876 18450
rect 29820 18386 29876 18398
rect 29484 17556 29540 17566
rect 29484 17462 29540 17500
rect 29596 17108 29652 18172
rect 29820 18226 29876 18238
rect 29820 18174 29822 18226
rect 29874 18174 29876 18226
rect 29820 17666 29876 18174
rect 29820 17614 29822 17666
rect 29874 17614 29876 17666
rect 29820 17602 29876 17614
rect 29708 17556 29764 17566
rect 29708 17462 29764 17500
rect 29932 17556 29988 17566
rect 29596 17106 29876 17108
rect 29596 17054 29598 17106
rect 29650 17054 29876 17106
rect 29596 17052 29876 17054
rect 29596 17042 29652 17052
rect 29484 16884 29540 16894
rect 29484 16212 29540 16828
rect 29596 16212 29652 16222
rect 29484 16210 29652 16212
rect 29484 16158 29598 16210
rect 29650 16158 29652 16210
rect 29484 16156 29652 16158
rect 29820 16212 29876 17052
rect 29932 17106 29988 17500
rect 29932 17054 29934 17106
rect 29986 17054 29988 17106
rect 29932 17042 29988 17054
rect 29932 16212 29988 16222
rect 29820 16210 29988 16212
rect 29820 16158 29934 16210
rect 29986 16158 29988 16210
rect 29820 16156 29988 16158
rect 29596 16146 29652 16156
rect 29932 16146 29988 16156
rect 29148 15988 29204 15998
rect 29148 15316 29204 15932
rect 30044 15652 30100 20300
rect 30156 19124 30212 20526
rect 30380 19796 30436 22540
rect 30492 21028 30548 23548
rect 30604 21698 30660 23660
rect 30716 22932 30772 29372
rect 30828 28980 30884 28990
rect 30828 27188 30884 28924
rect 30940 28644 30996 28654
rect 30940 28550 30996 28588
rect 31276 27972 31332 27982
rect 31164 27970 31332 27972
rect 31164 27918 31278 27970
rect 31330 27918 31332 27970
rect 31164 27916 31332 27918
rect 31164 27412 31220 27916
rect 31276 27906 31332 27916
rect 31500 27748 31556 34860
rect 31724 34692 31780 34702
rect 31724 34354 31780 34636
rect 31724 34302 31726 34354
rect 31778 34302 31780 34354
rect 31724 34290 31780 34302
rect 31836 34132 31892 34862
rect 31612 34018 31668 34030
rect 31612 33966 31614 34018
rect 31666 33966 31668 34018
rect 31612 33684 31668 33966
rect 31612 33618 31668 33628
rect 31724 33572 31780 33582
rect 31836 33572 31892 34076
rect 31724 33570 31892 33572
rect 31724 33518 31726 33570
rect 31778 33518 31892 33570
rect 31724 33516 31892 33518
rect 31724 33506 31780 33516
rect 31724 33236 31780 33246
rect 31724 33122 31780 33180
rect 31836 33236 31892 33246
rect 31836 33234 32116 33236
rect 31836 33182 31838 33234
rect 31890 33182 32116 33234
rect 31836 33180 32116 33182
rect 31836 33170 31892 33180
rect 31724 33070 31726 33122
rect 31778 33070 31780 33122
rect 31612 32564 31668 32574
rect 31612 30884 31668 32508
rect 31724 31108 31780 33070
rect 32060 32786 32116 33180
rect 32060 32734 32062 32786
rect 32114 32734 32116 32786
rect 32060 32722 32116 32734
rect 32172 32788 32228 39004
rect 32284 38668 32340 39228
rect 32508 39172 32564 40908
rect 32508 39106 32564 39116
rect 32620 39844 32676 39854
rect 32620 39618 32676 39788
rect 32620 39566 32622 39618
rect 32674 39566 32676 39618
rect 32508 38948 32564 38958
rect 32508 38854 32564 38892
rect 32620 38834 32676 39566
rect 32620 38782 32622 38834
rect 32674 38782 32676 38834
rect 32620 38770 32676 38782
rect 32732 38668 32788 41916
rect 32844 41878 32900 41916
rect 32844 41524 32900 41534
rect 33068 41524 33124 42590
rect 32900 41468 33124 41524
rect 32844 41298 32900 41468
rect 32844 41246 32846 41298
rect 32898 41246 32900 41298
rect 32844 41234 32900 41246
rect 32956 39508 33012 39518
rect 32284 38612 32452 38668
rect 32732 38612 32900 38668
rect 32284 38500 32340 38510
rect 32284 38274 32340 38444
rect 32284 38222 32286 38274
rect 32338 38222 32340 38274
rect 32284 38210 32340 38222
rect 32396 37492 32452 38612
rect 32284 37436 32452 37492
rect 32732 37826 32788 37838
rect 32732 37774 32734 37826
rect 32786 37774 32788 37826
rect 32284 33012 32340 37436
rect 32396 37268 32452 37278
rect 32732 37268 32788 37774
rect 32844 37380 32900 38612
rect 32956 37938 33012 39452
rect 33068 38052 33124 38062
rect 33068 37958 33124 37996
rect 32956 37886 32958 37938
rect 33010 37886 33012 37938
rect 32956 37874 33012 37886
rect 32844 37324 33012 37380
rect 32396 37266 32788 37268
rect 32396 37214 32398 37266
rect 32450 37214 32788 37266
rect 32396 37212 32788 37214
rect 32396 37202 32452 37212
rect 32844 37154 32900 37166
rect 32844 37102 32846 37154
rect 32898 37102 32900 37154
rect 32844 36484 32900 37102
rect 32844 36418 32900 36428
rect 32956 35922 33012 37324
rect 33180 36708 33236 44492
rect 33068 36652 33236 36708
rect 33292 44212 33348 44222
rect 33068 36148 33124 36652
rect 33180 36372 33236 36382
rect 33180 36278 33236 36316
rect 33068 36082 33124 36092
rect 32956 35870 32958 35922
rect 33010 35870 33012 35922
rect 32956 35858 33012 35870
rect 32732 35812 32788 35822
rect 32620 35700 32676 35710
rect 32620 35606 32676 35644
rect 32508 34916 32564 34926
rect 32564 34860 32676 34916
rect 32508 34822 32564 34860
rect 32620 34242 32676 34860
rect 32732 34692 32788 35756
rect 32788 34636 32900 34692
rect 32732 34626 32788 34636
rect 32732 34356 32788 34366
rect 32732 34262 32788 34300
rect 32620 34190 32622 34242
rect 32674 34190 32676 34242
rect 32620 34178 32676 34190
rect 32732 33348 32788 33358
rect 32844 33348 32900 34636
rect 32732 33346 32900 33348
rect 32732 33294 32734 33346
rect 32786 33294 32900 33346
rect 32732 33292 32900 33294
rect 32956 34130 33012 34142
rect 32956 34078 32958 34130
rect 33010 34078 33012 34130
rect 32732 33282 32788 33292
rect 32396 33124 32452 33134
rect 32396 33030 32452 33068
rect 32284 32946 32340 32956
rect 32172 32732 32452 32788
rect 32172 31220 32228 31230
rect 31724 31042 31780 31052
rect 32060 31108 32116 31118
rect 32060 31014 32116 31052
rect 31612 30790 31668 30828
rect 31948 30324 32004 30334
rect 31948 30210 32004 30268
rect 32172 30212 32228 31164
rect 31948 30158 31950 30210
rect 32002 30158 32004 30210
rect 31948 30146 32004 30158
rect 32060 30156 32228 30212
rect 31836 29988 31892 29998
rect 32060 29988 32116 30156
rect 32284 30098 32340 30110
rect 32284 30046 32286 30098
rect 32338 30046 32340 30098
rect 31836 29426 31892 29932
rect 31836 29374 31838 29426
rect 31890 29374 31892 29426
rect 31836 29362 31892 29374
rect 31948 29932 32116 29988
rect 32172 29986 32228 29998
rect 32172 29934 32174 29986
rect 32226 29934 32228 29986
rect 31724 28756 31780 28766
rect 31724 28642 31780 28700
rect 31724 28590 31726 28642
rect 31778 28590 31780 28642
rect 31724 28578 31780 28590
rect 31164 27346 31220 27356
rect 31276 27692 31556 27748
rect 30940 27188 30996 27198
rect 30828 27186 30996 27188
rect 30828 27134 30942 27186
rect 30994 27134 30996 27186
rect 30828 27132 30996 27134
rect 30828 26964 30884 27132
rect 30940 27122 30996 27132
rect 31164 27188 31220 27198
rect 30828 26898 30884 26908
rect 31164 25508 31220 27132
rect 31276 26068 31332 27692
rect 31948 27524 32004 29932
rect 32172 29428 32228 29934
rect 32060 29372 32228 29428
rect 32060 29314 32116 29372
rect 32284 29316 32340 30046
rect 32060 29262 32062 29314
rect 32114 29262 32116 29314
rect 32060 28754 32116 29262
rect 32060 28702 32062 28754
rect 32114 28702 32116 28754
rect 32060 28690 32116 28702
rect 32172 29260 32340 29316
rect 32172 28532 32228 29260
rect 32172 28466 32228 28476
rect 32284 28644 32340 28654
rect 32284 28530 32340 28588
rect 32284 28478 32286 28530
rect 32338 28478 32340 28530
rect 32284 28466 32340 28478
rect 32060 28420 32116 28430
rect 32060 28326 32116 28364
rect 31948 27458 32004 27468
rect 31388 27300 31444 27310
rect 31388 27186 31444 27244
rect 31388 27134 31390 27186
rect 31442 27134 31444 27186
rect 31388 27122 31444 27134
rect 32396 26908 32452 32732
rect 32956 32004 33012 34078
rect 33292 33796 33348 44156
rect 32956 31938 33012 31948
rect 33068 33740 33348 33796
rect 32620 30882 32676 30894
rect 32620 30830 32622 30882
rect 32674 30830 32676 30882
rect 32620 30324 32676 30830
rect 32620 30268 33012 30324
rect 32844 30098 32900 30110
rect 32844 30046 32846 30098
rect 32898 30046 32900 30098
rect 32844 29988 32900 30046
rect 32508 29932 32900 29988
rect 32508 29538 32564 29932
rect 32956 29652 33012 30268
rect 33068 30212 33124 33740
rect 33404 33684 33460 45388
rect 33516 44548 33572 45726
rect 33628 45780 33684 45948
rect 33628 45778 33796 45780
rect 33628 45726 33630 45778
rect 33682 45726 33796 45778
rect 33628 45724 33796 45726
rect 33628 45714 33684 45724
rect 33628 45108 33684 45118
rect 33628 45014 33684 45052
rect 33516 44482 33572 44492
rect 33516 44100 33572 44110
rect 33516 44006 33572 44044
rect 33516 43426 33572 43438
rect 33516 43374 33518 43426
rect 33570 43374 33572 43426
rect 33516 42980 33572 43374
rect 33516 42914 33572 42924
rect 33740 42082 33796 45724
rect 33852 45668 33908 45706
rect 33852 45602 33908 45612
rect 33740 42030 33742 42082
rect 33794 42030 33796 42082
rect 33740 41972 33796 42030
rect 33740 41906 33796 41916
rect 33852 45444 33908 45454
rect 33852 40740 33908 45388
rect 33964 45108 34020 46510
rect 33964 45042 34020 45052
rect 33964 42084 34020 42094
rect 33964 41990 34020 42028
rect 33852 40674 33908 40684
rect 33964 40516 34020 40526
rect 33964 40422 34020 40460
rect 33852 40404 33908 40414
rect 33628 40402 33908 40404
rect 33628 40350 33854 40402
rect 33906 40350 33908 40402
rect 33628 40348 33908 40350
rect 33628 39730 33684 40348
rect 33852 40338 33908 40348
rect 33964 40180 34020 40190
rect 34076 40180 34132 46844
rect 34188 45890 34244 47292
rect 34300 47124 34356 47406
rect 34748 47460 34804 47964
rect 34860 47684 34916 48414
rect 34972 48132 35028 49084
rect 35084 49028 35140 49644
rect 35196 49634 35252 49644
rect 35644 49698 35700 49710
rect 35644 49646 35646 49698
rect 35698 49646 35700 49698
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35084 48804 35140 48972
rect 35532 48804 35588 48814
rect 35084 48802 35476 48804
rect 35084 48750 35086 48802
rect 35138 48750 35476 48802
rect 35084 48748 35476 48750
rect 35084 48738 35140 48748
rect 35308 48132 35364 48142
rect 34972 48076 35140 48132
rect 34860 47618 34916 47628
rect 34972 47460 35028 47470
rect 34748 47458 35028 47460
rect 34748 47406 34974 47458
rect 35026 47406 35028 47458
rect 34748 47404 35028 47406
rect 34972 47394 35028 47404
rect 34300 47058 34356 47068
rect 35084 47012 35140 48076
rect 35308 48038 35364 48076
rect 35420 48018 35476 48748
rect 35532 48710 35588 48748
rect 35420 47966 35422 48018
rect 35474 47966 35476 48018
rect 35420 47954 35476 47966
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35196 47460 35252 47470
rect 35196 47366 35252 47404
rect 35420 47458 35476 47470
rect 35420 47406 35422 47458
rect 35474 47406 35476 47458
rect 35420 47236 35476 47406
rect 35532 47460 35588 47470
rect 35532 47366 35588 47404
rect 35420 47170 35476 47180
rect 35084 46946 35140 46956
rect 34412 46900 34468 46910
rect 34412 46806 34468 46844
rect 34636 46900 34692 46910
rect 34524 45892 34580 45902
rect 34188 45838 34190 45890
rect 34242 45838 34244 45890
rect 34188 45826 34244 45838
rect 34300 45890 34580 45892
rect 34300 45838 34526 45890
rect 34578 45838 34580 45890
rect 34300 45836 34580 45838
rect 34300 45218 34356 45836
rect 34524 45826 34580 45836
rect 34524 45666 34580 45678
rect 34524 45614 34526 45666
rect 34578 45614 34580 45666
rect 34524 45332 34580 45614
rect 34636 45444 34692 46844
rect 34860 46562 34916 46574
rect 34860 46510 34862 46562
rect 34914 46510 34916 46562
rect 34860 46004 34916 46510
rect 35308 46564 35364 46574
rect 35308 46470 35364 46508
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 34860 45938 34916 45948
rect 34636 45378 34692 45388
rect 34860 45778 34916 45790
rect 34860 45726 34862 45778
rect 34914 45726 34916 45778
rect 34524 45266 34580 45276
rect 34300 45166 34302 45218
rect 34354 45166 34356 45218
rect 34300 43538 34356 45166
rect 34860 45220 34916 45726
rect 35308 45780 35364 45790
rect 35308 45686 35364 45724
rect 34860 45154 34916 45164
rect 34412 45106 34468 45118
rect 34412 45054 34414 45106
rect 34466 45054 34468 45106
rect 34412 43652 34468 45054
rect 34524 45108 34580 45118
rect 34524 45014 34580 45052
rect 34972 45108 35028 45118
rect 34972 45014 35028 45052
rect 35532 45108 35588 45118
rect 35532 45014 35588 45052
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35644 44660 35700 49646
rect 35756 46788 35812 50372
rect 36540 50036 36596 50046
rect 36652 50036 36708 51212
rect 36540 50034 36708 50036
rect 36540 49982 36542 50034
rect 36594 49982 36708 50034
rect 36540 49980 36708 49982
rect 36540 49970 36596 49980
rect 36316 49924 36372 49934
rect 36316 49138 36372 49868
rect 36316 49086 36318 49138
rect 36370 49086 36372 49138
rect 36316 49028 36372 49086
rect 36316 48962 36372 48972
rect 35868 48468 35924 48478
rect 35868 48374 35924 48412
rect 36428 48468 36484 48478
rect 36428 48244 36484 48412
rect 36652 48356 36708 49980
rect 36764 49810 36820 51438
rect 36876 51156 36932 51166
rect 36876 51062 36932 51100
rect 36764 49758 36766 49810
rect 36818 49758 36820 49810
rect 36764 49476 36820 49758
rect 36764 49410 36820 49420
rect 37100 49140 37156 55412
rect 37548 55410 37940 55412
rect 37548 55358 37886 55410
rect 37938 55358 37940 55410
rect 37548 55356 37940 55358
rect 37884 55346 37940 55356
rect 37436 55076 37492 55086
rect 37324 55074 37492 55076
rect 37324 55022 37438 55074
rect 37490 55022 37492 55074
rect 37324 55020 37492 55022
rect 37324 53732 37380 55020
rect 37436 55010 37492 55020
rect 37772 54628 37828 54638
rect 37772 54534 37828 54572
rect 37660 54404 37716 54414
rect 37548 54402 37716 54404
rect 37548 54350 37662 54402
rect 37714 54350 37716 54402
rect 37548 54348 37716 54350
rect 37324 53666 37380 53676
rect 37436 53844 37492 53854
rect 37324 53396 37380 53406
rect 37324 52948 37380 53340
rect 37436 53172 37492 53788
rect 37548 53842 37604 54348
rect 37660 54338 37716 54348
rect 37548 53790 37550 53842
rect 37602 53790 37604 53842
rect 37548 53778 37604 53790
rect 37660 53730 37716 53742
rect 37996 53732 38052 53742
rect 37660 53678 37662 53730
rect 37714 53678 37716 53730
rect 37660 53396 37716 53678
rect 37660 53330 37716 53340
rect 37772 53730 38052 53732
rect 37772 53678 37998 53730
rect 38050 53678 38052 53730
rect 37772 53676 38052 53678
rect 37548 53172 37604 53182
rect 37436 53170 37604 53172
rect 37436 53118 37550 53170
rect 37602 53118 37604 53170
rect 37436 53116 37604 53118
rect 37548 53106 37604 53116
rect 37772 53172 37828 53676
rect 37996 53666 38052 53676
rect 37436 52948 37492 52958
rect 37324 52946 37492 52948
rect 37324 52894 37438 52946
rect 37490 52894 37492 52946
rect 37324 52892 37492 52894
rect 37436 52836 37492 52892
rect 37772 52946 37828 53116
rect 38220 53060 38276 53070
rect 38220 52966 38276 53004
rect 37772 52894 37774 52946
rect 37826 52894 37828 52946
rect 37772 52882 37828 52894
rect 37436 52770 37492 52780
rect 37548 52388 37604 52398
rect 37548 52274 37604 52332
rect 37548 52222 37550 52274
rect 37602 52222 37604 52274
rect 37548 52210 37604 52222
rect 37660 52052 37716 52062
rect 37660 51938 37716 51996
rect 37660 51886 37662 51938
rect 37714 51886 37716 51938
rect 37212 51604 37268 51614
rect 37212 50428 37268 51548
rect 37324 51266 37380 51278
rect 37324 51214 37326 51266
rect 37378 51214 37380 51266
rect 37324 50596 37380 51214
rect 37660 51156 37716 51886
rect 38108 51940 38164 51950
rect 38108 51490 38164 51884
rect 38108 51438 38110 51490
rect 38162 51438 38164 51490
rect 37884 51156 37940 51166
rect 37660 51154 37940 51156
rect 37660 51102 37886 51154
rect 37938 51102 37940 51154
rect 37660 51100 37940 51102
rect 37436 50708 37492 50718
rect 37436 50614 37492 50652
rect 37884 50596 37940 51100
rect 38108 50932 38164 51438
rect 38220 51380 38276 51390
rect 38220 51266 38276 51324
rect 38220 51214 38222 51266
rect 38274 51214 38276 51266
rect 38220 51202 38276 51214
rect 38332 50932 38388 55412
rect 38556 55188 38612 55198
rect 38444 55186 38612 55188
rect 38444 55134 38558 55186
rect 38610 55134 38612 55186
rect 38444 55132 38612 55134
rect 38444 55076 38500 55132
rect 38556 55122 38612 55132
rect 38444 54514 38500 55020
rect 38444 54462 38446 54514
rect 38498 54462 38500 54514
rect 38444 54450 38500 54462
rect 38668 53060 38724 57820
rect 39228 57764 39284 57774
rect 38780 56420 38836 56430
rect 38780 56306 38836 56364
rect 38780 56254 38782 56306
rect 38834 56254 38836 56306
rect 38780 56242 38836 56254
rect 39116 55524 39172 55534
rect 38892 55410 38948 55422
rect 38892 55358 38894 55410
rect 38946 55358 38948 55410
rect 38892 55300 38948 55358
rect 38892 55234 38948 55244
rect 38780 55074 38836 55086
rect 38780 55022 38782 55074
rect 38834 55022 38836 55074
rect 38780 54628 38836 55022
rect 38780 54514 38836 54572
rect 38780 54462 38782 54514
rect 38834 54462 38836 54514
rect 38780 54450 38836 54462
rect 39116 53170 39172 55468
rect 39116 53118 39118 53170
rect 39170 53118 39172 53170
rect 39116 53106 39172 53118
rect 39228 53172 39284 57708
rect 39452 56308 39508 56318
rect 39452 56214 39508 56252
rect 39788 56082 39844 56094
rect 39788 56030 39790 56082
rect 39842 56030 39844 56082
rect 39788 55972 39844 56030
rect 39788 55906 39844 55916
rect 40124 55468 40180 58268
rect 40348 56642 40404 59200
rect 42812 57988 42868 57998
rect 40348 56590 40350 56642
rect 40402 56590 40404 56642
rect 40348 56578 40404 56590
rect 40684 57316 40740 57326
rect 40236 55972 40292 55982
rect 40236 55878 40292 55916
rect 40124 55412 40292 55468
rect 39340 55298 39396 55310
rect 39340 55246 39342 55298
rect 39394 55246 39396 55298
rect 39340 54740 39396 55246
rect 39564 55300 39620 55310
rect 39396 54684 39508 54740
rect 39340 54674 39396 54684
rect 39340 54516 39396 54526
rect 39340 54422 39396 54460
rect 39452 53954 39508 54684
rect 39452 53902 39454 53954
rect 39506 53902 39508 53954
rect 39452 53890 39508 53902
rect 39564 53954 39620 55244
rect 40012 55300 40068 55310
rect 39564 53902 39566 53954
rect 39618 53902 39620 53954
rect 39564 53890 39620 53902
rect 39788 55074 39844 55086
rect 39788 55022 39790 55074
rect 39842 55022 39844 55074
rect 39788 54404 39844 55022
rect 39900 55076 39956 55086
rect 39900 54982 39956 55020
rect 40012 54516 40068 55244
rect 40124 54516 40180 54526
rect 40012 54514 40180 54516
rect 40012 54462 40126 54514
rect 40178 54462 40180 54514
rect 40012 54460 40180 54462
rect 40124 54450 40180 54460
rect 39900 54404 39956 54414
rect 39788 54402 39956 54404
rect 39788 54350 39902 54402
rect 39954 54350 39956 54402
rect 39788 54348 39956 54350
rect 39788 53844 39844 54348
rect 39900 54338 39956 54348
rect 39788 53750 39844 53788
rect 40124 54292 40180 54302
rect 40012 53732 40068 53742
rect 39900 53620 39956 53630
rect 39900 53526 39956 53564
rect 39564 53172 39620 53182
rect 39228 53170 39620 53172
rect 39228 53118 39566 53170
rect 39618 53118 39620 53170
rect 39228 53116 39620 53118
rect 39564 53106 39620 53116
rect 40012 53170 40068 53676
rect 40012 53118 40014 53170
rect 40066 53118 40068 53170
rect 40012 53106 40068 53118
rect 38668 53004 39060 53060
rect 38668 52836 38724 52846
rect 38668 52742 38724 52780
rect 38444 52052 38500 52062
rect 38444 51958 38500 51996
rect 38556 51940 38612 51950
rect 38556 51846 38612 51884
rect 38780 51940 38836 51950
rect 38780 51938 38948 51940
rect 38780 51886 38782 51938
rect 38834 51886 38948 51938
rect 38780 51884 38948 51886
rect 38780 51874 38836 51884
rect 38892 51490 38948 51884
rect 38892 51438 38894 51490
rect 38946 51438 38948 51490
rect 38892 51426 38948 51438
rect 38108 50866 38164 50876
rect 38220 50876 38388 50932
rect 38780 51378 38836 51390
rect 38780 51326 38782 51378
rect 38834 51326 38836 51378
rect 38108 50706 38164 50718
rect 38108 50654 38110 50706
rect 38162 50654 38164 50706
rect 38108 50596 38164 50654
rect 37884 50540 38164 50596
rect 37324 50530 37380 50540
rect 37212 50372 37380 50428
rect 37100 49074 37156 49084
rect 37324 49698 37380 50372
rect 37884 50036 37940 50046
rect 37884 49942 37940 49980
rect 38220 50036 38276 50876
rect 38332 50484 38388 50494
rect 38332 50390 38388 50428
rect 38780 50260 38836 51326
rect 38780 50194 38836 50204
rect 39004 50036 39060 53004
rect 40012 52276 40068 52286
rect 40124 52276 40180 54236
rect 40012 52274 40180 52276
rect 40012 52222 40014 52274
rect 40066 52222 40180 52274
rect 40012 52220 40180 52222
rect 40012 52210 40068 52220
rect 39228 51938 39284 51950
rect 39564 51940 39620 51950
rect 39228 51886 39230 51938
rect 39282 51886 39284 51938
rect 39228 50260 39284 51886
rect 39228 50194 39284 50204
rect 39452 51938 39620 51940
rect 39452 51886 39566 51938
rect 39618 51886 39620 51938
rect 39452 51884 39620 51886
rect 39116 50036 39172 50046
rect 39004 50034 39172 50036
rect 39004 49982 39118 50034
rect 39170 49982 39172 50034
rect 39004 49980 39172 49982
rect 38220 49970 38276 49980
rect 39116 49970 39172 49980
rect 37324 49646 37326 49698
rect 37378 49646 37380 49698
rect 36988 48916 37044 48926
rect 36876 48802 36932 48814
rect 36876 48750 36878 48802
rect 36930 48750 36932 48802
rect 36876 48580 36932 48750
rect 36876 48514 36932 48524
rect 36652 48300 36932 48356
rect 36428 48242 36596 48244
rect 36428 48190 36430 48242
rect 36482 48190 36596 48242
rect 36428 48188 36596 48190
rect 36428 48178 36484 48188
rect 36204 48018 36260 48030
rect 36204 47966 36206 48018
rect 36258 47966 36260 48018
rect 35756 46722 35812 46732
rect 35980 47236 36036 47246
rect 36092 47236 36148 47246
rect 36036 47234 36148 47236
rect 36036 47182 36094 47234
rect 36146 47182 36148 47234
rect 36036 47180 36148 47182
rect 36204 47236 36260 47966
rect 36540 47572 36596 48188
rect 36876 48242 36932 48300
rect 36988 48354 37044 48860
rect 37324 48468 37380 49646
rect 38220 49700 38276 49710
rect 38220 49606 38276 49644
rect 38668 49700 38724 49710
rect 38668 49698 38836 49700
rect 38668 49646 38670 49698
rect 38722 49646 38836 49698
rect 38668 49644 38836 49646
rect 38668 49634 38724 49644
rect 38668 49476 38724 49486
rect 37772 49028 37828 49038
rect 37772 48934 37828 48972
rect 38108 49028 38164 49038
rect 37548 48914 37604 48926
rect 37548 48862 37550 48914
rect 37602 48862 37604 48914
rect 37548 48468 37604 48862
rect 37884 48802 37940 48814
rect 37884 48750 37886 48802
rect 37938 48750 37940 48802
rect 37884 48692 37940 48750
rect 37884 48626 37940 48636
rect 37996 48802 38052 48814
rect 37996 48750 37998 48802
rect 38050 48750 38052 48802
rect 37996 48468 38052 48750
rect 36988 48302 36990 48354
rect 37042 48302 37044 48354
rect 36988 48290 37044 48302
rect 37100 48412 37604 48468
rect 37772 48412 38052 48468
rect 38108 48468 38164 48972
rect 36876 48190 36878 48242
rect 36930 48190 36932 48242
rect 36876 48178 36932 48190
rect 36988 48132 37044 48142
rect 36428 47236 36484 47246
rect 36204 47234 36484 47236
rect 36204 47182 36430 47234
rect 36482 47182 36484 47234
rect 36204 47180 36484 47182
rect 35756 46564 35812 46574
rect 35756 46562 35924 46564
rect 35756 46510 35758 46562
rect 35810 46510 35924 46562
rect 35756 46508 35924 46510
rect 35756 46498 35812 46508
rect 35756 45332 35812 45342
rect 35756 45106 35812 45276
rect 35756 45054 35758 45106
rect 35810 45054 35812 45106
rect 35756 45042 35812 45054
rect 35644 44594 35700 44604
rect 35644 44436 35700 44446
rect 35644 44342 35700 44380
rect 35868 44324 35924 46508
rect 35980 44882 36036 47180
rect 36092 47170 36148 47180
rect 36316 45444 36372 47180
rect 36428 47170 36484 47180
rect 36540 46898 36596 47516
rect 36652 48018 36708 48030
rect 36652 47966 36654 48018
rect 36706 47966 36708 48018
rect 36652 47460 36708 47966
rect 36652 47394 36708 47404
rect 36764 47908 36820 47918
rect 36540 46846 36542 46898
rect 36594 46846 36596 46898
rect 36540 46834 36596 46846
rect 36652 47124 36708 47134
rect 36428 45892 36484 45902
rect 36428 45798 36484 45836
rect 36540 45668 36596 45678
rect 36652 45668 36708 47068
rect 36764 45890 36820 47852
rect 36988 47124 37044 48076
rect 36988 47058 37044 47068
rect 36764 45838 36766 45890
rect 36818 45838 36820 45890
rect 36764 45826 36820 45838
rect 36876 46788 36932 46798
rect 36652 45612 36820 45668
rect 36540 45574 36596 45612
rect 36652 45444 36708 45454
rect 36316 45388 36596 45444
rect 35980 44830 35982 44882
rect 36034 44830 36036 44882
rect 35980 44660 36036 44830
rect 36092 44884 36148 44894
rect 36092 44790 36148 44828
rect 35980 44604 36260 44660
rect 36204 44324 36260 44604
rect 35868 44268 36148 44324
rect 34412 43586 34468 43596
rect 35532 44210 35588 44222
rect 35532 44158 35534 44210
rect 35586 44158 35588 44210
rect 34300 43486 34302 43538
rect 34354 43486 34356 43538
rect 34188 43428 34244 43438
rect 34188 42756 34244 43372
rect 34300 42868 34356 43486
rect 34524 43538 34580 43550
rect 34524 43486 34526 43538
rect 34578 43486 34580 43538
rect 34524 43428 34580 43486
rect 34636 43540 34692 43550
rect 34636 43446 34692 43484
rect 34972 43540 35028 43550
rect 34524 43362 34580 43372
rect 34860 43316 34916 43326
rect 34300 42812 34692 42868
rect 34636 42756 34692 42812
rect 34860 42866 34916 43260
rect 34860 42814 34862 42866
rect 34914 42814 34916 42866
rect 34860 42802 34916 42814
rect 34188 42700 34468 42756
rect 34412 42644 34468 42700
rect 34636 42690 34692 42700
rect 34412 42512 34468 42588
rect 34972 42642 35028 43484
rect 35084 43540 35140 43550
rect 35532 43540 35588 44158
rect 35756 44212 35812 44222
rect 35756 44210 36036 44212
rect 35756 44158 35758 44210
rect 35810 44158 36036 44210
rect 35756 44156 36036 44158
rect 35756 44146 35812 44156
rect 35980 43988 36036 44156
rect 35868 43932 36036 43988
rect 35644 43540 35700 43550
rect 35084 43538 35700 43540
rect 35084 43486 35086 43538
rect 35138 43486 35646 43538
rect 35698 43486 35700 43538
rect 35084 43484 35700 43486
rect 35084 43474 35140 43484
rect 35644 43474 35700 43484
rect 35868 43316 35924 43932
rect 36092 43540 36148 44268
rect 36204 44322 36372 44324
rect 36204 44270 36206 44322
rect 36258 44270 36372 44322
rect 36204 44268 36372 44270
rect 36204 44258 36260 44268
rect 35868 43222 35924 43260
rect 35980 43484 36148 43540
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34972 42590 34974 42642
rect 35026 42590 35028 42642
rect 34860 42532 34916 42542
rect 34188 42308 34244 42318
rect 34188 42194 34244 42252
rect 34188 42142 34190 42194
rect 34242 42142 34244 42194
rect 34188 42130 34244 42142
rect 34860 42194 34916 42476
rect 34972 42420 35028 42590
rect 34972 42354 35028 42364
rect 35196 42980 35252 42990
rect 35196 42196 35252 42924
rect 35980 42868 36036 43484
rect 36092 43314 36148 43326
rect 36092 43262 36094 43314
rect 36146 43262 36148 43314
rect 36092 43204 36148 43262
rect 36204 43316 36260 43326
rect 36204 43222 36260 43260
rect 36092 43138 36148 43148
rect 36316 42980 36372 44268
rect 36540 43428 36596 45388
rect 36652 45106 36708 45388
rect 36652 45054 36654 45106
rect 36706 45054 36708 45106
rect 36652 45042 36708 45054
rect 36764 44548 36820 45612
rect 36652 44492 36820 44548
rect 36652 43876 36708 44492
rect 36764 44324 36820 44334
rect 36764 44230 36820 44268
rect 36652 43652 36708 43820
rect 36652 43596 36820 43652
rect 36652 43428 36708 43438
rect 36540 43426 36708 43428
rect 36540 43374 36654 43426
rect 36706 43374 36708 43426
rect 36540 43372 36708 43374
rect 36652 43204 36708 43372
rect 36652 43138 36708 43148
rect 36764 42980 36820 43596
rect 36316 42914 36372 42924
rect 36540 42924 36820 42980
rect 35980 42812 36148 42868
rect 34860 42142 34862 42194
rect 34914 42142 34916 42194
rect 34860 42130 34916 42142
rect 34972 42140 35252 42196
rect 35308 42700 35588 42756
rect 34300 42084 34356 42094
rect 34300 41990 34356 42028
rect 34860 40628 34916 40638
rect 34636 40516 34692 40526
rect 33964 40178 34132 40180
rect 33964 40126 33966 40178
rect 34018 40126 34132 40178
rect 33964 40124 34132 40126
rect 34188 40292 34244 40302
rect 33964 40114 34020 40124
rect 33628 39678 33630 39730
rect 33682 39678 33684 39730
rect 33628 39666 33684 39678
rect 33740 39618 33796 39630
rect 33740 39566 33742 39618
rect 33794 39566 33796 39618
rect 33740 38948 33796 39566
rect 33740 38882 33796 38892
rect 34188 39618 34244 40236
rect 34188 39566 34190 39618
rect 34242 39566 34244 39618
rect 34188 38722 34244 39566
rect 34636 38948 34692 40460
rect 34188 38670 34190 38722
rect 34242 38670 34244 38722
rect 33516 38500 33572 38510
rect 33516 38162 33572 38444
rect 34188 38274 34244 38670
rect 34188 38222 34190 38274
rect 34242 38222 34244 38274
rect 34188 38210 34244 38222
rect 34300 38946 34692 38948
rect 34300 38894 34638 38946
rect 34690 38894 34692 38946
rect 34300 38892 34692 38894
rect 33516 38110 33518 38162
rect 33570 38110 33572 38162
rect 33516 38098 33572 38110
rect 33964 38052 34020 38062
rect 33964 37958 34020 37996
rect 33964 37154 34020 37166
rect 33964 37102 33966 37154
rect 34018 37102 34020 37154
rect 33964 36708 34020 37102
rect 33964 36642 34020 36652
rect 33628 36484 33684 36494
rect 33628 36390 33684 36428
rect 33740 36372 33796 36382
rect 33740 36278 33796 36316
rect 33964 36258 34020 36270
rect 33964 36206 33966 36258
rect 34018 36206 34020 36258
rect 33740 36148 33796 36158
rect 33628 35812 33684 35822
rect 33628 35698 33684 35756
rect 33628 35646 33630 35698
rect 33682 35646 33684 35698
rect 33628 35634 33684 35646
rect 33740 34916 33796 36092
rect 33964 36148 34020 36206
rect 33964 36082 34020 36092
rect 34188 35924 34244 35934
rect 34300 35924 34356 38892
rect 34636 38882 34692 38892
rect 34524 38274 34580 38286
rect 34524 38222 34526 38274
rect 34578 38222 34580 38274
rect 34524 38162 34580 38222
rect 34524 38110 34526 38162
rect 34578 38110 34580 38162
rect 34524 38098 34580 38110
rect 34860 38164 34916 40572
rect 34972 40626 35028 42140
rect 35308 42084 35364 42700
rect 35532 42642 35588 42700
rect 35532 42590 35534 42642
rect 35586 42590 35588 42642
rect 35532 42578 35588 42590
rect 35756 42644 35812 42654
rect 35756 42550 35812 42588
rect 35980 42644 36036 42654
rect 35980 42550 36036 42588
rect 34972 40574 34974 40626
rect 35026 40574 35028 40626
rect 34972 40562 35028 40574
rect 35084 42028 35364 42084
rect 35420 42530 35476 42542
rect 35420 42478 35422 42530
rect 35474 42478 35476 42530
rect 35420 42084 35476 42478
rect 35756 42196 35812 42206
rect 35084 41970 35140 42028
rect 35420 42018 35476 42028
rect 35644 42084 35700 42094
rect 35084 41918 35086 41970
rect 35138 41918 35140 41970
rect 35084 40292 35140 41918
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35532 41300 35588 41310
rect 35644 41300 35700 42028
rect 35756 42082 35812 42140
rect 35756 42030 35758 42082
rect 35810 42030 35812 42082
rect 35756 42018 35812 42030
rect 35868 42084 35924 42094
rect 35868 41990 35924 42028
rect 35532 41298 35700 41300
rect 35532 41246 35534 41298
rect 35586 41246 35700 41298
rect 35532 41244 35700 41246
rect 35868 41746 35924 41758
rect 35868 41694 35870 41746
rect 35922 41694 35924 41746
rect 35532 41234 35588 41244
rect 34972 40236 35140 40292
rect 34972 38948 35028 40236
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 34972 38882 35028 38892
rect 35084 39394 35140 39406
rect 35084 39342 35086 39394
rect 35138 39342 35140 39394
rect 35084 38274 35140 39342
rect 35532 38948 35588 38958
rect 35532 38834 35588 38892
rect 35532 38782 35534 38834
rect 35586 38782 35588 38834
rect 35532 38770 35588 38782
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35084 38222 35086 38274
rect 35138 38222 35140 38274
rect 35084 38210 35140 38222
rect 34972 38164 35028 38174
rect 34860 38162 35028 38164
rect 34860 38110 34974 38162
rect 35026 38110 35028 38162
rect 34860 38108 35028 38110
rect 34188 35922 34356 35924
rect 34188 35870 34190 35922
rect 34242 35870 34356 35922
rect 34188 35868 34356 35870
rect 34412 37378 34468 37390
rect 34412 37326 34414 37378
rect 34466 37326 34468 37378
rect 34188 35858 34244 35868
rect 33852 35700 33908 35710
rect 33852 35606 33908 35644
rect 33180 33628 33460 33684
rect 33628 34860 33796 34916
rect 33964 35588 34020 35598
rect 33180 31220 33236 33628
rect 33404 33348 33460 33358
rect 33404 32564 33460 33292
rect 33516 32564 33572 32574
rect 33404 32508 33516 32564
rect 33516 32470 33572 32508
rect 33180 31154 33236 31164
rect 33404 32340 33460 32350
rect 33180 30884 33236 30894
rect 33180 30434 33236 30828
rect 33180 30382 33182 30434
rect 33234 30382 33236 30434
rect 33180 30370 33236 30382
rect 33068 30156 33348 30212
rect 33068 29986 33124 29998
rect 33068 29934 33070 29986
rect 33122 29934 33124 29986
rect 33068 29652 33124 29934
rect 32508 29486 32510 29538
rect 32562 29486 32564 29538
rect 32508 29474 32564 29486
rect 32844 29596 33124 29652
rect 32844 29428 32900 29596
rect 33292 29428 33348 30156
rect 32844 29362 32900 29372
rect 32956 29372 33348 29428
rect 32732 28644 32788 28654
rect 32172 26852 32228 26862
rect 32172 26758 32228 26796
rect 32284 26852 32452 26908
rect 32508 28420 32564 28430
rect 32508 28082 32564 28364
rect 32508 28030 32510 28082
rect 32562 28030 32564 28082
rect 32508 26908 32564 28030
rect 32732 27186 32788 28588
rect 32732 27134 32734 27186
rect 32786 27134 32788 27186
rect 32508 26852 32676 26908
rect 31276 26002 31332 26012
rect 31500 26514 31556 26526
rect 31500 26462 31502 26514
rect 31554 26462 31556 26514
rect 31500 25618 31556 26462
rect 32060 26404 32116 26414
rect 32060 26310 32116 26348
rect 31500 25566 31502 25618
rect 31554 25566 31556 25618
rect 31500 25508 31556 25566
rect 31164 25506 31444 25508
rect 31164 25454 31166 25506
rect 31218 25454 31444 25506
rect 31164 25452 31444 25454
rect 31164 25442 31220 25452
rect 31388 24946 31444 25452
rect 31500 25442 31556 25452
rect 31612 26290 31668 26302
rect 31612 26238 31614 26290
rect 31666 26238 31668 26290
rect 31388 24894 31390 24946
rect 31442 24894 31444 24946
rect 31388 24882 31444 24894
rect 31612 24724 31668 26238
rect 32284 25844 32340 26852
rect 32508 26292 32564 26302
rect 32508 26198 32564 26236
rect 32284 25778 32340 25788
rect 32620 25732 32676 26852
rect 32732 25844 32788 27134
rect 32732 25778 32788 25788
rect 32844 26852 32900 26862
rect 31836 25396 31892 25406
rect 31836 25302 31892 25340
rect 32396 25396 32452 25406
rect 32396 25302 32452 25340
rect 32620 25394 32676 25676
rect 32620 25342 32622 25394
rect 32674 25342 32676 25394
rect 32620 25330 32676 25342
rect 32732 25396 32788 25406
rect 32732 25302 32788 25340
rect 32844 25394 32900 26796
rect 32956 25620 33012 29372
rect 33404 28868 33460 32284
rect 33628 31780 33684 34860
rect 33740 34690 33796 34702
rect 33740 34638 33742 34690
rect 33794 34638 33796 34690
rect 33740 33124 33796 34638
rect 33852 33348 33908 33358
rect 33964 33348 34020 35532
rect 34412 35588 34468 37326
rect 34748 37380 34804 37390
rect 34860 37380 34916 38108
rect 34972 38098 35028 38108
rect 34748 37378 34916 37380
rect 34748 37326 34750 37378
rect 34802 37326 34916 37378
rect 34748 37324 34916 37326
rect 35420 37380 35476 37390
rect 35420 37378 35588 37380
rect 35420 37326 35422 37378
rect 35474 37326 35588 37378
rect 35420 37324 35588 37326
rect 34636 36482 34692 36494
rect 34636 36430 34638 36482
rect 34690 36430 34692 36482
rect 34636 36148 34692 36430
rect 34748 36372 34804 37324
rect 35420 37314 35476 37324
rect 35084 37268 35140 37278
rect 34748 36306 34804 36316
rect 34860 36708 34916 36718
rect 34860 36594 34916 36652
rect 34860 36542 34862 36594
rect 34914 36542 34916 36594
rect 34636 36082 34692 36092
rect 34860 35700 34916 36542
rect 35084 35922 35140 37212
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35084 35870 35086 35922
rect 35138 35870 35140 35922
rect 35084 35858 35140 35870
rect 35420 36484 35476 36494
rect 35420 35924 35476 36428
rect 35532 35924 35588 37324
rect 35644 37268 35700 37278
rect 35644 37174 35700 37212
rect 35868 37268 35924 41694
rect 36092 38668 36148 42812
rect 36316 42084 36372 42094
rect 36316 41298 36372 42028
rect 36540 42084 36596 42924
rect 36876 42308 36932 46732
rect 36988 45892 37044 45902
rect 36988 45106 37044 45836
rect 36988 45054 36990 45106
rect 37042 45054 37044 45106
rect 36988 44436 37044 45054
rect 36988 44370 37044 44380
rect 36540 41952 36596 42028
rect 36652 42252 36932 42308
rect 36316 41246 36318 41298
rect 36370 41246 36372 41298
rect 36316 41234 36372 41246
rect 36540 40628 36596 40638
rect 36652 40628 36708 42252
rect 36876 42084 36932 42094
rect 37100 42084 37156 48412
rect 37772 48356 37828 48412
rect 37436 48354 37828 48356
rect 37436 48302 37774 48354
rect 37826 48302 37828 48354
rect 37436 48300 37828 48302
rect 37436 47682 37492 48300
rect 37772 48290 37828 48300
rect 37884 48242 37940 48254
rect 37884 48190 37886 48242
rect 37938 48190 37940 48242
rect 37548 48132 37604 48142
rect 37548 48038 37604 48076
rect 37884 48020 37940 48190
rect 38108 48242 38164 48412
rect 38108 48190 38110 48242
rect 38162 48190 38164 48242
rect 38108 48178 38164 48190
rect 38220 49026 38276 49038
rect 38220 48974 38222 49026
rect 38274 48974 38276 49026
rect 38220 48020 38276 48974
rect 38668 48802 38724 49420
rect 38668 48750 38670 48802
rect 38722 48750 38724 48802
rect 38556 48356 38612 48366
rect 38556 48262 38612 48300
rect 37884 47964 38276 48020
rect 37884 47796 37940 47964
rect 37436 47630 37438 47682
rect 37490 47630 37492 47682
rect 37436 47618 37492 47630
rect 37660 47740 37940 47796
rect 37212 47460 37268 47470
rect 37212 46674 37268 47404
rect 37212 46622 37214 46674
rect 37266 46622 37268 46674
rect 37212 46610 37268 46622
rect 37436 47012 37492 47022
rect 37436 46674 37492 46956
rect 37660 46786 37716 47740
rect 37884 47572 37940 47582
rect 37940 47516 38052 47572
rect 37884 47478 37940 47516
rect 37884 47124 37940 47134
rect 37660 46734 37662 46786
rect 37714 46734 37716 46786
rect 37660 46722 37716 46734
rect 37772 47012 37828 47022
rect 37436 46622 37438 46674
rect 37490 46622 37492 46674
rect 37436 46610 37492 46622
rect 37548 45668 37604 45678
rect 37212 45218 37268 45230
rect 37212 45166 37214 45218
rect 37266 45166 37268 45218
rect 37212 45108 37268 45166
rect 37212 45052 37492 45108
rect 37436 44996 37492 45052
rect 37548 44996 37604 45612
rect 37660 44996 37716 45006
rect 37436 44994 37716 44996
rect 37436 44942 37662 44994
rect 37714 44942 37716 44994
rect 37436 44940 37716 44942
rect 37324 44882 37380 44894
rect 37324 44830 37326 44882
rect 37378 44830 37380 44882
rect 37324 44324 37380 44830
rect 37324 44258 37380 44268
rect 37212 43764 37268 43774
rect 37212 43670 37268 43708
rect 36876 42082 37156 42084
rect 36876 42030 36878 42082
rect 36930 42030 37156 42082
rect 36876 42028 37156 42030
rect 37436 42308 37492 42318
rect 37436 42082 37492 42252
rect 37436 42030 37438 42082
rect 37490 42030 37492 42082
rect 36876 41860 36932 42028
rect 37436 42018 37492 42030
rect 36876 41794 36932 41804
rect 36596 40572 36708 40628
rect 37100 40964 37156 40974
rect 36540 40496 36596 40572
rect 36876 40404 36932 40414
rect 36876 40310 36932 40348
rect 36876 39844 36932 39854
rect 36876 39730 36932 39788
rect 36876 39678 36878 39730
rect 36930 39678 36932 39730
rect 36876 39060 36932 39678
rect 36876 38994 36932 39004
rect 36988 39172 37044 39182
rect 36988 38946 37044 39116
rect 36988 38894 36990 38946
rect 37042 38894 37044 38946
rect 36204 38836 36260 38846
rect 36876 38836 36932 38846
rect 36204 38834 36932 38836
rect 36204 38782 36206 38834
rect 36258 38782 36878 38834
rect 36930 38782 36932 38834
rect 36204 38780 36932 38782
rect 36204 38770 36260 38780
rect 36876 38770 36932 38780
rect 36092 38612 36260 38668
rect 35868 37266 36036 37268
rect 35868 37214 35870 37266
rect 35922 37214 36036 37266
rect 35868 37212 36036 37214
rect 35868 37202 35924 37212
rect 35756 37154 35812 37166
rect 35756 37102 35758 37154
rect 35810 37102 35812 37154
rect 35756 36596 35812 37102
rect 35756 36530 35812 36540
rect 35980 36482 36036 37212
rect 35980 36430 35982 36482
rect 36034 36430 36036 36482
rect 35980 36418 36036 36430
rect 35756 35924 35812 35934
rect 35532 35922 35812 35924
rect 35532 35870 35758 35922
rect 35810 35870 35812 35922
rect 35532 35868 35812 35870
rect 34412 35522 34468 35532
rect 34524 35698 34916 35700
rect 34524 35646 34862 35698
rect 34914 35646 34916 35698
rect 34524 35644 34916 35646
rect 34524 35026 34580 35644
rect 34860 35476 34916 35644
rect 34972 35698 35028 35710
rect 34972 35646 34974 35698
rect 35026 35646 35028 35698
rect 34972 35588 35028 35646
rect 35420 35698 35476 35868
rect 35756 35858 35812 35868
rect 36092 35924 36148 35934
rect 36092 35830 36148 35868
rect 35420 35646 35422 35698
rect 35474 35646 35476 35698
rect 35420 35634 35476 35646
rect 35868 35810 35924 35822
rect 35868 35758 35870 35810
rect 35922 35758 35924 35810
rect 34972 35522 35028 35532
rect 35868 35588 35924 35758
rect 35868 35522 35924 35532
rect 34860 35410 34916 35420
rect 35644 35476 35700 35486
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 34524 34974 34526 35026
rect 34578 34974 34580 35026
rect 34524 34962 34580 34974
rect 35644 35026 35700 35420
rect 35644 34974 35646 35026
rect 35698 34974 35700 35026
rect 35644 34962 35700 34974
rect 34188 34692 34244 34702
rect 33852 33346 34020 33348
rect 33852 33294 33854 33346
rect 33906 33294 34020 33346
rect 33852 33292 34020 33294
rect 33852 33282 33908 33292
rect 33740 33058 33796 33068
rect 33628 31714 33684 31724
rect 33852 32004 33908 32014
rect 33852 31778 33908 31948
rect 33852 31726 33854 31778
rect 33906 31726 33908 31778
rect 33852 31714 33908 31726
rect 33964 31666 34020 33292
rect 34076 34242 34132 34254
rect 34076 34190 34078 34242
rect 34130 34190 34132 34242
rect 34076 33124 34132 34190
rect 34076 33058 34132 33068
rect 34188 32788 34244 34636
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 36204 32900 36260 38612
rect 36764 38164 36820 38174
rect 36764 38070 36820 38108
rect 36988 36708 37044 38894
rect 36988 36642 37044 36652
rect 36764 36372 36820 36382
rect 36764 36278 36820 36316
rect 37100 35924 37156 40908
rect 37548 40516 37604 44940
rect 37660 44930 37716 44940
rect 37772 44660 37828 46956
rect 37884 46674 37940 47068
rect 37996 46786 38052 47516
rect 38108 47460 38164 47470
rect 38108 47366 38164 47404
rect 38332 47458 38388 47470
rect 38332 47406 38334 47458
rect 38386 47406 38388 47458
rect 37996 46734 37998 46786
rect 38050 46734 38052 46786
rect 37996 46722 38052 46734
rect 38220 47124 38276 47134
rect 37884 46622 37886 46674
rect 37938 46622 37940 46674
rect 37884 46610 37940 46622
rect 38108 46452 38164 46462
rect 38108 45330 38164 46396
rect 38108 45278 38110 45330
rect 38162 45278 38164 45330
rect 38108 45266 38164 45278
rect 37772 44604 38164 44660
rect 37660 43540 37716 43550
rect 37660 43446 37716 43484
rect 37772 43204 37828 44604
rect 38108 44546 38164 44604
rect 38108 44494 38110 44546
rect 38162 44494 38164 44546
rect 38108 44482 38164 44494
rect 37660 43148 37828 43204
rect 37884 44210 37940 44222
rect 37884 44158 37886 44210
rect 37938 44158 37940 44210
rect 37884 43540 37940 44158
rect 37996 43764 38052 43774
rect 37996 43670 38052 43708
rect 37660 42196 37716 43148
rect 37772 42642 37828 42654
rect 37772 42590 37774 42642
rect 37826 42590 37828 42642
rect 37772 42308 37828 42590
rect 37772 42242 37828 42252
rect 37660 42084 37716 42140
rect 37772 42084 37828 42094
rect 37660 42082 37828 42084
rect 37660 42030 37774 42082
rect 37826 42030 37828 42082
rect 37660 42028 37828 42030
rect 37772 42018 37828 42028
rect 37772 41188 37828 41198
rect 37884 41188 37940 43484
rect 38108 42756 38164 42766
rect 38108 42642 38164 42700
rect 38108 42590 38110 42642
rect 38162 42590 38164 42642
rect 38108 42578 38164 42590
rect 38220 41972 38276 47068
rect 38332 47012 38388 47406
rect 38556 47346 38612 47358
rect 38556 47294 38558 47346
rect 38610 47294 38612 47346
rect 38556 47124 38612 47294
rect 38556 47058 38612 47068
rect 38332 46946 38388 46956
rect 38668 46900 38724 48750
rect 38668 46834 38724 46844
rect 38780 46676 38836 49644
rect 39452 49588 39508 51884
rect 39564 51874 39620 51884
rect 39788 51604 39844 51614
rect 40236 51604 40292 55412
rect 40460 55076 40516 55086
rect 40460 55074 40628 55076
rect 40460 55022 40462 55074
rect 40514 55022 40628 55074
rect 40460 55020 40628 55022
rect 40460 55010 40516 55020
rect 40348 54740 40404 54750
rect 40348 54514 40404 54684
rect 40348 54462 40350 54514
rect 40402 54462 40404 54514
rect 40348 54450 40404 54462
rect 40348 53508 40404 53518
rect 40348 53506 40516 53508
rect 40348 53454 40350 53506
rect 40402 53454 40516 53506
rect 40348 53452 40516 53454
rect 40348 53442 40404 53452
rect 40460 52164 40516 53452
rect 40460 52070 40516 52108
rect 40572 51716 40628 55020
rect 40684 52276 40740 57260
rect 41132 56642 41188 56654
rect 41132 56590 41134 56642
rect 41186 56590 41188 56642
rect 41132 56194 41188 56590
rect 41132 56142 41134 56194
rect 41186 56142 41188 56194
rect 41132 56130 41188 56142
rect 42812 56306 42868 57932
rect 42812 56254 42814 56306
rect 42866 56254 42868 56306
rect 42252 56082 42308 56094
rect 42252 56030 42254 56082
rect 42306 56030 42308 56082
rect 41804 55748 41860 55758
rect 41132 55188 41188 55198
rect 40796 55186 41188 55188
rect 40796 55134 41134 55186
rect 41186 55134 41188 55186
rect 40796 55132 41188 55134
rect 40796 54738 40852 55132
rect 41132 55122 41188 55132
rect 40796 54686 40798 54738
rect 40850 54686 40852 54738
rect 40796 54674 40852 54686
rect 41244 55076 41300 55086
rect 41132 54292 41188 54302
rect 41132 53730 41188 54236
rect 41132 53678 41134 53730
rect 41186 53678 41188 53730
rect 41132 53666 41188 53678
rect 40908 53620 40964 53630
rect 41244 53620 41300 55020
rect 41468 55074 41524 55086
rect 41468 55022 41470 55074
rect 41522 55022 41524 55074
rect 41468 54180 41524 55022
rect 41468 54114 41524 54124
rect 41356 53620 41412 53630
rect 41244 53618 41412 53620
rect 41244 53566 41358 53618
rect 41410 53566 41412 53618
rect 41244 53564 41412 53566
rect 40908 53526 40964 53564
rect 41356 53554 41412 53564
rect 41020 53506 41076 53518
rect 41020 53454 41022 53506
rect 41074 53454 41076 53506
rect 41020 53172 41076 53454
rect 41804 53508 41860 55692
rect 41916 55074 41972 55086
rect 41916 55022 41918 55074
rect 41970 55022 41972 55074
rect 41916 54740 41972 55022
rect 42252 54740 42308 56030
rect 41916 54684 42196 54740
rect 42140 54628 42196 54684
rect 42252 54674 42308 54684
rect 42364 55972 42420 55982
rect 42028 54516 42084 54526
rect 42028 54422 42084 54460
rect 42140 54402 42196 54572
rect 42140 54350 42142 54402
rect 42194 54350 42196 54402
rect 42140 53956 42196 54350
rect 42140 53890 42196 53900
rect 42364 53732 42420 55916
rect 42812 55636 42868 56254
rect 43596 56196 43652 56206
rect 43596 56102 43652 56140
rect 46396 56196 46452 59200
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 46396 56130 46452 56140
rect 47292 56196 47348 56206
rect 46620 56082 46676 56094
rect 46620 56030 46622 56082
rect 46674 56030 46676 56082
rect 42812 55570 42868 55580
rect 43148 55970 43204 55982
rect 43148 55918 43150 55970
rect 43202 55918 43204 55970
rect 43148 55468 43204 55918
rect 46172 55972 46228 55982
rect 46620 55972 46676 56030
rect 46172 55970 46676 55972
rect 46172 55918 46174 55970
rect 46226 55918 46676 55970
rect 46172 55916 46676 55918
rect 46172 55906 46228 55916
rect 43484 55860 43540 55870
rect 43148 55412 43316 55468
rect 43148 55300 43204 55310
rect 42924 55244 43148 55300
rect 42476 55188 42532 55198
rect 42476 55094 42532 55132
rect 42924 54628 42980 55244
rect 43148 55206 43204 55244
rect 42812 54626 42980 54628
rect 42812 54574 42926 54626
rect 42978 54574 42980 54626
rect 42812 54572 42980 54574
rect 42700 53956 42756 53966
rect 42812 53956 42868 54572
rect 42924 54562 42980 54572
rect 43036 55076 43092 55086
rect 42700 53954 42868 53956
rect 42700 53902 42702 53954
rect 42754 53902 42868 53954
rect 42700 53900 42868 53902
rect 42924 53956 42980 53966
rect 43036 53956 43092 55020
rect 42924 53954 43092 53956
rect 42924 53902 42926 53954
rect 42978 53902 43092 53954
rect 42924 53900 43092 53902
rect 43148 54180 43204 54190
rect 42700 53890 42756 53900
rect 42924 53890 42980 53900
rect 42028 53676 42420 53732
rect 43148 53730 43204 54124
rect 43148 53678 43150 53730
rect 43202 53678 43204 53730
rect 41916 53508 41972 53518
rect 41804 53506 41972 53508
rect 41804 53454 41918 53506
rect 41970 53454 41972 53506
rect 41804 53452 41972 53454
rect 41020 53116 41860 53172
rect 40796 53060 40852 53070
rect 40852 53004 41300 53060
rect 40796 52966 40852 53004
rect 40908 52276 40964 52286
rect 40684 52274 40964 52276
rect 40684 52222 40910 52274
rect 40962 52222 40964 52274
rect 40684 52220 40964 52222
rect 40908 52210 40964 52220
rect 40572 51650 40628 51660
rect 40348 51604 40404 51614
rect 40236 51602 40404 51604
rect 40236 51550 40350 51602
rect 40402 51550 40404 51602
rect 40236 51548 40404 51550
rect 39788 51510 39844 51548
rect 40348 51538 40404 51548
rect 39676 51380 39732 51390
rect 39676 51286 39732 51324
rect 40796 51268 40852 51278
rect 40684 51266 40852 51268
rect 40684 51214 40798 51266
rect 40850 51214 40852 51266
rect 40684 51212 40852 51214
rect 39564 50594 39620 50606
rect 39564 50542 39566 50594
rect 39618 50542 39620 50594
rect 39564 50260 39620 50542
rect 39564 50194 39620 50204
rect 40236 50482 40292 50494
rect 40236 50430 40238 50482
rect 40290 50430 40292 50482
rect 40236 50148 40292 50430
rect 40236 50092 40628 50148
rect 39564 50036 39620 50046
rect 39564 49942 39620 49980
rect 40572 50034 40628 50092
rect 40572 49982 40574 50034
rect 40626 49982 40628 50034
rect 39452 49522 39508 49532
rect 40124 49810 40180 49822
rect 40124 49758 40126 49810
rect 40178 49758 40180 49810
rect 39788 49028 39844 49038
rect 38892 48468 38948 48478
rect 38892 48374 38948 48412
rect 39788 48356 39844 48972
rect 40124 49028 40180 49758
rect 40348 49810 40404 49822
rect 40348 49758 40350 49810
rect 40402 49758 40404 49810
rect 40236 49700 40292 49710
rect 40236 49606 40292 49644
rect 40124 48962 40180 48972
rect 40236 49028 40292 49038
rect 40348 49028 40404 49758
rect 40572 49252 40628 49982
rect 40684 49476 40740 51212
rect 40796 51202 40852 51212
rect 40796 50372 40852 50382
rect 40796 50370 40964 50372
rect 40796 50318 40798 50370
rect 40850 50318 40964 50370
rect 40796 50316 40964 50318
rect 40796 50306 40852 50316
rect 40908 49924 40964 50316
rect 40908 49858 40964 49868
rect 40684 49410 40740 49420
rect 40684 49252 40740 49262
rect 40572 49250 40740 49252
rect 40572 49198 40686 49250
rect 40738 49198 40740 49250
rect 40572 49196 40740 49198
rect 40684 49186 40740 49196
rect 40236 49026 40404 49028
rect 40236 48974 40238 49026
rect 40290 48974 40404 49026
rect 40236 48972 40404 48974
rect 40460 49028 40516 49038
rect 40236 48916 40292 48972
rect 40460 48934 40516 48972
rect 40236 48850 40292 48860
rect 41132 48916 41188 48926
rect 41132 48822 41188 48860
rect 39788 48262 39844 48300
rect 40012 48692 40068 48702
rect 40012 48242 40068 48636
rect 40012 48190 40014 48242
rect 40066 48190 40068 48242
rect 40012 48178 40068 48190
rect 40348 48132 40404 48142
rect 40348 48038 40404 48076
rect 39228 48020 39284 48030
rect 39004 47572 39060 47582
rect 39004 47478 39060 47516
rect 39228 47124 39284 47964
rect 41020 47796 41076 47806
rect 40460 47516 40740 47572
rect 39676 47348 39732 47358
rect 39676 47254 39732 47292
rect 39228 46900 39284 47068
rect 38780 46610 38836 46620
rect 39004 46898 39284 46900
rect 39004 46846 39230 46898
rect 39282 46846 39284 46898
rect 39004 46844 39284 46846
rect 39004 46002 39060 46844
rect 39228 46834 39284 46844
rect 40124 47124 40180 47134
rect 40012 46674 40068 46686
rect 40012 46622 40014 46674
rect 40066 46622 40068 46674
rect 39004 45950 39006 46002
rect 39058 45950 39060 46002
rect 39004 45938 39060 45950
rect 39676 46004 39732 46014
rect 39676 45910 39732 45948
rect 39452 45890 39508 45902
rect 39452 45838 39454 45890
rect 39506 45838 39508 45890
rect 38332 45666 38388 45678
rect 38332 45614 38334 45666
rect 38386 45614 38388 45666
rect 38332 45332 38388 45614
rect 39452 45556 39508 45838
rect 39900 45778 39956 45790
rect 39900 45726 39902 45778
rect 39954 45726 39956 45778
rect 39452 45490 39508 45500
rect 39788 45556 39844 45566
rect 38332 45266 38388 45276
rect 38892 45332 38948 45342
rect 38892 45238 38948 45276
rect 39228 45108 39284 45118
rect 39004 44996 39060 45006
rect 39004 44902 39060 44940
rect 38332 44884 38388 44894
rect 38332 44548 38388 44828
rect 38668 44884 38724 44894
rect 38668 44882 38948 44884
rect 38668 44830 38670 44882
rect 38722 44830 38948 44882
rect 38668 44828 38948 44830
rect 38668 44818 38724 44828
rect 38332 44546 38500 44548
rect 38332 44494 38334 44546
rect 38386 44494 38500 44546
rect 38332 44492 38500 44494
rect 38332 44482 38388 44492
rect 38444 43708 38500 44492
rect 38556 44436 38612 44446
rect 38556 44322 38612 44380
rect 38556 44270 38558 44322
rect 38610 44270 38612 44322
rect 38556 44212 38612 44270
rect 38556 44146 38612 44156
rect 38444 43652 38724 43708
rect 37772 41186 37940 41188
rect 37772 41134 37774 41186
rect 37826 41134 37940 41186
rect 37772 41132 37940 41134
rect 37772 41122 37828 41132
rect 37772 40516 37828 40526
rect 37548 40514 37828 40516
rect 37548 40462 37774 40514
rect 37826 40462 37828 40514
rect 37548 40460 37828 40462
rect 37436 40404 37492 40414
rect 37436 39844 37492 40348
rect 37548 39844 37604 39854
rect 37436 39842 37604 39844
rect 37436 39790 37550 39842
rect 37602 39790 37604 39842
rect 37436 39788 37604 39790
rect 37548 39778 37604 39788
rect 37660 39844 37716 39854
rect 37660 39730 37716 39788
rect 37660 39678 37662 39730
rect 37714 39678 37716 39730
rect 37660 39666 37716 39678
rect 37772 39172 37828 40460
rect 37884 39844 37940 41132
rect 37996 41916 38220 41972
rect 37996 41074 38052 41916
rect 38220 41906 38276 41916
rect 38444 43540 38500 43550
rect 38444 42532 38500 43484
rect 38668 43538 38724 43652
rect 38668 43486 38670 43538
rect 38722 43486 38724 43538
rect 38668 43474 38724 43486
rect 38892 43314 38948 44828
rect 39004 44548 39060 44558
rect 39004 44454 39060 44492
rect 39228 43764 39284 45052
rect 39564 45106 39620 45118
rect 39564 45054 39566 45106
rect 39618 45054 39620 45106
rect 39564 44884 39620 45054
rect 39788 45106 39844 45500
rect 39900 45220 39956 45726
rect 40012 45668 40068 46622
rect 40124 45892 40180 47068
rect 40460 46898 40516 47516
rect 40460 46846 40462 46898
rect 40514 46846 40516 46898
rect 40460 46834 40516 46846
rect 40572 47348 40628 47358
rect 40348 46674 40404 46686
rect 40348 46622 40350 46674
rect 40402 46622 40404 46674
rect 40348 46004 40404 46622
rect 40572 46676 40628 47292
rect 40684 47236 40740 47516
rect 41020 47458 41076 47740
rect 41020 47406 41022 47458
rect 41074 47406 41076 47458
rect 41020 47236 41076 47406
rect 40684 47180 41076 47236
rect 40572 46674 41076 46676
rect 40572 46622 40574 46674
rect 40626 46622 41076 46674
rect 40572 46620 41076 46622
rect 40572 46610 40628 46620
rect 40348 45938 40404 45948
rect 40124 45890 40292 45892
rect 40124 45838 40126 45890
rect 40178 45838 40292 45890
rect 40124 45836 40292 45838
rect 40124 45826 40180 45836
rect 40012 45612 40180 45668
rect 40124 45330 40180 45612
rect 40124 45278 40126 45330
rect 40178 45278 40180 45330
rect 40124 45266 40180 45278
rect 40012 45220 40068 45230
rect 39900 45218 40068 45220
rect 39900 45166 40014 45218
rect 40066 45166 40068 45218
rect 39900 45164 40068 45166
rect 39788 45054 39790 45106
rect 39842 45054 39844 45106
rect 39788 45042 39844 45054
rect 40012 45108 40068 45164
rect 40012 45042 40068 45052
rect 40236 44884 40292 45836
rect 40460 44996 40516 45006
rect 40460 44994 40628 44996
rect 40460 44942 40462 44994
rect 40514 44942 40628 44994
rect 40460 44940 40628 44942
rect 40460 44930 40516 44940
rect 39564 44828 40292 44884
rect 39228 43538 39284 43708
rect 39452 44436 39508 44446
rect 39452 43652 39508 44380
rect 40124 44436 40180 44446
rect 40236 44436 40292 44828
rect 40124 44434 40292 44436
rect 40124 44382 40126 44434
rect 40178 44382 40292 44434
rect 40124 44380 40292 44382
rect 39676 44324 39732 44334
rect 39676 44230 39732 44268
rect 39900 43652 39956 43662
rect 39452 43650 39956 43652
rect 39452 43598 39454 43650
rect 39506 43598 39902 43650
rect 39954 43598 39956 43650
rect 39452 43596 39956 43598
rect 39452 43586 39508 43596
rect 39900 43586 39956 43596
rect 40124 43652 40180 44380
rect 40124 43586 40180 43596
rect 40460 43764 40516 43774
rect 39228 43486 39230 43538
rect 39282 43486 39284 43538
rect 39228 43474 39284 43486
rect 38892 43262 38894 43314
rect 38946 43262 38948 43314
rect 38892 42756 38948 43262
rect 39340 43428 39396 43438
rect 39340 43314 39396 43372
rect 40348 43426 40404 43438
rect 40348 43374 40350 43426
rect 40402 43374 40404 43426
rect 39340 43262 39342 43314
rect 39394 43262 39396 43314
rect 39340 43250 39396 43262
rect 39676 43314 39732 43326
rect 39676 43262 39678 43314
rect 39730 43262 39732 43314
rect 38892 42690 38948 42700
rect 39116 43204 39172 43214
rect 38444 41298 38500 42476
rect 38444 41246 38446 41298
rect 38498 41246 38500 41298
rect 38444 41234 38500 41246
rect 38556 42530 38612 42542
rect 38556 42478 38558 42530
rect 38610 42478 38612 42530
rect 38556 41300 38612 42478
rect 39004 42532 39060 42542
rect 39004 42438 39060 42476
rect 38892 42196 38948 42206
rect 38668 41972 38724 41982
rect 38668 41878 38724 41916
rect 38892 41970 38948 42140
rect 38892 41918 38894 41970
rect 38946 41918 38948 41970
rect 38892 41906 38948 41918
rect 39116 41970 39172 43148
rect 39564 42756 39620 42766
rect 39116 41918 39118 41970
rect 39170 41918 39172 41970
rect 39116 41906 39172 41918
rect 39228 41972 39284 41982
rect 38668 41300 38724 41310
rect 38556 41244 38668 41300
rect 37996 41022 37998 41074
rect 38050 41022 38052 41074
rect 37996 41010 38052 41022
rect 38668 40626 38724 41244
rect 39004 41300 39060 41310
rect 39004 41206 39060 41244
rect 39228 41186 39284 41916
rect 39340 41746 39396 41758
rect 39340 41694 39342 41746
rect 39394 41694 39396 41746
rect 39340 41300 39396 41694
rect 39564 41410 39620 42700
rect 39564 41358 39566 41410
rect 39618 41358 39620 41410
rect 39564 41346 39620 41358
rect 39676 42754 39732 43262
rect 39676 42702 39678 42754
rect 39730 42702 39732 42754
rect 39340 41234 39396 41244
rect 39676 41300 39732 42702
rect 39900 43316 39956 43326
rect 39900 42978 39956 43260
rect 40348 43314 40404 43374
rect 40348 43262 40350 43314
rect 40402 43262 40404 43314
rect 40348 43250 40404 43262
rect 39900 42926 39902 42978
rect 39954 42926 39956 42978
rect 39788 41748 39844 41758
rect 39788 41654 39844 41692
rect 39788 41412 39844 41422
rect 39900 41412 39956 42926
rect 40348 42980 40404 42990
rect 40460 42980 40516 43708
rect 40572 43540 40628 44940
rect 41020 44322 41076 46620
rect 41020 44270 41022 44322
rect 41074 44270 41076 44322
rect 41020 44258 41076 44270
rect 41132 45780 41188 45790
rect 41132 43708 41188 45724
rect 41244 45332 41300 53004
rect 41580 52948 41636 52958
rect 41580 52854 41636 52892
rect 41804 52946 41860 53116
rect 41804 52894 41806 52946
rect 41858 52894 41860 52946
rect 41804 52882 41860 52894
rect 41580 52724 41636 52734
rect 41580 52274 41636 52668
rect 41580 52222 41582 52274
rect 41634 52222 41636 52274
rect 41244 45266 41300 45276
rect 41356 52164 41412 52174
rect 40796 43652 40852 43662
rect 41132 43652 41300 43708
rect 40796 43558 40852 43596
rect 40572 43474 40628 43484
rect 40348 42978 41076 42980
rect 40348 42926 40350 42978
rect 40402 42926 41076 42978
rect 40348 42924 41076 42926
rect 40348 42914 40404 42924
rect 41020 42866 41076 42924
rect 41020 42814 41022 42866
rect 41074 42814 41076 42866
rect 41020 42802 41076 42814
rect 40124 42756 40180 42766
rect 40124 42662 40180 42700
rect 40236 42530 40292 42542
rect 40236 42478 40238 42530
rect 40290 42478 40292 42530
rect 40236 42082 40292 42478
rect 40236 42030 40238 42082
rect 40290 42030 40292 42082
rect 40236 42018 40292 42030
rect 40684 42084 40740 42094
rect 40684 41990 40740 42028
rect 40460 41972 40516 41982
rect 39788 41410 39956 41412
rect 39788 41358 39790 41410
rect 39842 41358 39956 41410
rect 39788 41356 39956 41358
rect 40348 41916 40460 41972
rect 39788 41346 39844 41356
rect 39676 41234 39732 41244
rect 39228 41134 39230 41186
rect 39282 41134 39284 41186
rect 39228 41122 39284 41134
rect 40012 41076 40068 41086
rect 39900 40964 39956 40974
rect 39900 40870 39956 40908
rect 38668 40574 38670 40626
rect 38722 40574 38724 40626
rect 38668 40562 38724 40574
rect 40012 40628 40068 41020
rect 40348 41076 40404 41916
rect 40460 41840 40516 41916
rect 40796 41970 40852 41982
rect 40796 41918 40798 41970
rect 40850 41918 40852 41970
rect 40572 41748 40628 41758
rect 40348 41010 40404 41020
rect 40460 41074 40516 41086
rect 40460 41022 40462 41074
rect 40514 41022 40516 41074
rect 40460 40964 40516 41022
rect 40572 41074 40628 41692
rect 40796 41300 40852 41918
rect 40572 41022 40574 41074
rect 40626 41022 40628 41074
rect 40572 41010 40628 41022
rect 40684 41244 40852 41300
rect 40460 40898 40516 40908
rect 40684 40964 40740 41244
rect 40684 40898 40740 40908
rect 40796 40964 40852 40974
rect 40796 40962 40964 40964
rect 40796 40910 40798 40962
rect 40850 40910 40964 40962
rect 40796 40908 40964 40910
rect 40796 40898 40852 40908
rect 40796 40628 40852 40638
rect 40012 40496 40068 40572
rect 40684 40572 40796 40628
rect 37884 39778 37940 39788
rect 40684 39730 40740 40572
rect 40796 40534 40852 40572
rect 40908 40292 40964 40908
rect 40908 40226 40964 40236
rect 40684 39678 40686 39730
rect 40738 39678 40740 39730
rect 40684 39666 40740 39678
rect 40796 39844 40852 39854
rect 38892 39618 38948 39630
rect 38892 39566 38894 39618
rect 38946 39566 38948 39618
rect 37772 39106 37828 39116
rect 38108 39394 38164 39406
rect 38108 39342 38110 39394
rect 38162 39342 38164 39394
rect 38108 39172 38164 39342
rect 38108 39106 38164 39116
rect 38892 39058 38948 39566
rect 39340 39620 39396 39630
rect 39340 39526 39396 39564
rect 40572 39620 40628 39630
rect 40572 39526 40628 39564
rect 39228 39396 39284 39406
rect 38892 39006 38894 39058
rect 38946 39006 38948 39058
rect 38892 38994 38948 39006
rect 39004 39394 39284 39396
rect 39004 39342 39230 39394
rect 39282 39342 39284 39394
rect 39004 39340 39284 39342
rect 37212 38948 37268 38958
rect 38332 38948 38388 38958
rect 37212 38946 38388 38948
rect 37212 38894 37214 38946
rect 37266 38894 38334 38946
rect 38386 38894 38388 38946
rect 37212 38892 38388 38894
rect 37212 38882 37268 38892
rect 37660 38722 37716 38734
rect 37660 38670 37662 38722
rect 37714 38670 37716 38722
rect 37660 38668 37716 38670
rect 37548 38612 37716 38668
rect 37772 38724 37828 38734
rect 37548 37604 37604 38612
rect 37548 37490 37604 37548
rect 37548 37438 37550 37490
rect 37602 37438 37604 37490
rect 37548 37426 37604 37438
rect 37212 35924 37268 35934
rect 36988 35922 37604 35924
rect 36988 35870 37214 35922
rect 37266 35870 37604 35922
rect 36988 35868 37604 35870
rect 36316 35698 36372 35710
rect 36316 35646 36318 35698
rect 36370 35646 36372 35698
rect 36316 35476 36372 35646
rect 36316 35410 36372 35420
rect 36988 35252 37044 35868
rect 37212 35858 37268 35868
rect 36876 35196 37044 35252
rect 36764 34690 36820 34702
rect 36764 34638 36766 34690
rect 36818 34638 36820 34690
rect 36764 34468 36820 34638
rect 36764 34402 36820 34412
rect 36316 34018 36372 34030
rect 36316 33966 36318 34018
rect 36370 33966 36372 34018
rect 36316 33348 36372 33966
rect 36316 33282 36372 33292
rect 36764 34020 36820 34030
rect 36316 33124 36372 33134
rect 36316 33122 36484 33124
rect 36316 33070 36318 33122
rect 36370 33070 36484 33122
rect 36316 33068 36484 33070
rect 36316 33058 36372 33068
rect 36204 32844 36372 32900
rect 33964 31614 33966 31666
rect 34018 31614 34020 31666
rect 33964 31602 34020 31614
rect 34076 32732 34244 32788
rect 34076 30434 34132 32732
rect 34188 32562 34244 32574
rect 34188 32510 34190 32562
rect 34242 32510 34244 32562
rect 34188 31778 34244 32510
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 34188 31726 34190 31778
rect 34242 31726 34244 31778
rect 34188 31714 34244 31726
rect 36204 31108 36260 31118
rect 35420 30882 35476 30894
rect 35420 30830 35422 30882
rect 35474 30830 35476 30882
rect 35420 30770 35476 30830
rect 35868 30884 35924 30894
rect 35868 30882 36036 30884
rect 35868 30830 35870 30882
rect 35922 30830 36036 30882
rect 35868 30828 36036 30830
rect 35868 30818 35924 30828
rect 35420 30718 35422 30770
rect 35474 30718 35476 30770
rect 35420 30706 35476 30718
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34076 30382 34078 30434
rect 34130 30382 34132 30434
rect 34076 30370 34132 30382
rect 33740 30324 33796 30334
rect 33740 30230 33796 30268
rect 35308 30324 35364 30334
rect 35084 30098 35140 30110
rect 35084 30046 35086 30098
rect 35138 30046 35140 30098
rect 33964 29986 34020 29998
rect 33964 29934 33966 29986
rect 34018 29934 34020 29986
rect 33516 29428 33572 29438
rect 33516 29334 33572 29372
rect 33964 29428 34020 29934
rect 34524 29986 34580 29998
rect 34524 29934 34526 29986
rect 34578 29934 34580 29986
rect 34524 29876 34580 29934
rect 34524 29810 34580 29820
rect 35084 29876 35140 30046
rect 35084 29810 35140 29820
rect 35196 29986 35252 29998
rect 35196 29934 35198 29986
rect 35250 29934 35252 29986
rect 35196 29652 35252 29934
rect 34972 29596 35252 29652
rect 35308 29650 35364 30268
rect 35420 30100 35476 30110
rect 35868 30100 35924 30110
rect 35420 30098 35924 30100
rect 35420 30046 35422 30098
rect 35474 30046 35870 30098
rect 35922 30046 35924 30098
rect 35420 30044 35924 30046
rect 35420 30034 35476 30044
rect 35868 30034 35924 30044
rect 35980 29876 36036 30828
rect 36092 30770 36148 30782
rect 36092 30718 36094 30770
rect 36146 30718 36148 30770
rect 36092 30100 36148 30718
rect 36204 30324 36260 31052
rect 36204 30258 36260 30268
rect 36092 30098 36260 30100
rect 36092 30046 36094 30098
rect 36146 30046 36260 30098
rect 36092 30044 36260 30046
rect 36092 30034 36148 30044
rect 35980 29810 36036 29820
rect 35308 29598 35310 29650
rect 35362 29598 35364 29650
rect 33964 29362 34020 29372
rect 34860 29428 34916 29438
rect 34972 29428 35028 29596
rect 35308 29586 35364 29598
rect 35532 29764 35588 29774
rect 35532 29540 35588 29708
rect 35532 29538 35700 29540
rect 35532 29486 35534 29538
rect 35586 29486 35700 29538
rect 35532 29484 35700 29486
rect 35532 29474 35588 29484
rect 34860 29426 35028 29428
rect 34860 29374 34862 29426
rect 34914 29374 35028 29426
rect 34860 29372 35028 29374
rect 35084 29426 35140 29438
rect 35084 29374 35086 29426
rect 35138 29374 35140 29426
rect 34076 29314 34132 29326
rect 34076 29262 34078 29314
rect 34130 29262 34132 29314
rect 33292 28812 33460 28868
rect 33516 29092 33572 29102
rect 33292 27076 33348 28812
rect 33404 28644 33460 28654
rect 33404 28530 33460 28588
rect 33404 28478 33406 28530
rect 33458 28478 33460 28530
rect 33404 28466 33460 28478
rect 33292 27010 33348 27020
rect 33516 26908 33572 29036
rect 33628 28420 33684 28430
rect 33628 28082 33684 28364
rect 33628 28030 33630 28082
rect 33682 28030 33684 28082
rect 33628 28018 33684 28030
rect 33740 28418 33796 28430
rect 33740 28366 33742 28418
rect 33794 28366 33796 28418
rect 33740 27972 33796 28366
rect 33740 27906 33796 27916
rect 34076 27972 34132 29262
rect 34636 28868 34692 28878
rect 34636 28644 34692 28812
rect 34076 27906 34132 27916
rect 34524 28642 34692 28644
rect 34524 28590 34638 28642
rect 34690 28590 34692 28642
rect 34524 28588 34692 28590
rect 33964 27858 34020 27870
rect 33964 27806 33966 27858
rect 34018 27806 34020 27858
rect 33964 27748 34020 27806
rect 33964 27682 34020 27692
rect 34076 27636 34132 27646
rect 34076 27074 34132 27580
rect 34524 27188 34580 28588
rect 34636 28578 34692 28588
rect 34636 27634 34692 27646
rect 34636 27582 34638 27634
rect 34690 27582 34692 27634
rect 34636 27300 34692 27582
rect 34748 27636 34804 27646
rect 34860 27636 34916 29372
rect 35084 28756 35140 29374
rect 35420 29428 35476 29438
rect 35420 29204 35476 29372
rect 35420 29202 35588 29204
rect 35420 29150 35422 29202
rect 35474 29150 35588 29202
rect 35420 29148 35588 29150
rect 35420 29138 35476 29148
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35084 28690 35140 28700
rect 35196 28644 35252 28654
rect 35532 28644 35588 29148
rect 35644 28866 35700 29484
rect 35644 28814 35646 28866
rect 35698 28814 35700 28866
rect 35644 28802 35700 28814
rect 35756 28868 35812 28878
rect 35756 28754 35812 28812
rect 35980 28866 36036 28878
rect 35980 28814 35982 28866
rect 36034 28814 36036 28866
rect 35756 28702 35758 28754
rect 35810 28702 35812 28754
rect 35756 28690 35812 28702
rect 35868 28756 35924 28766
rect 35196 28642 35588 28644
rect 35196 28590 35198 28642
rect 35250 28590 35588 28642
rect 35196 28588 35588 28590
rect 35644 28644 35700 28654
rect 35196 28578 35252 28588
rect 35084 28532 35140 28542
rect 35644 28532 35700 28588
rect 35084 28438 35140 28476
rect 35532 28476 35700 28532
rect 34972 28420 35028 28430
rect 34972 27860 35028 28364
rect 35084 27860 35140 27870
rect 34972 27858 35140 27860
rect 34972 27806 35086 27858
rect 35138 27806 35140 27858
rect 34972 27804 35140 27806
rect 35084 27794 35140 27804
rect 35196 27748 35252 27758
rect 34804 27580 34916 27636
rect 34972 27636 35028 27646
rect 35196 27636 35252 27692
rect 34972 27634 35252 27636
rect 34972 27582 34974 27634
rect 35026 27582 35252 27634
rect 34972 27580 35252 27582
rect 34748 27542 34804 27580
rect 34972 27570 35028 27580
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 34636 27244 35140 27300
rect 34524 27132 34804 27188
rect 34076 27022 34078 27074
rect 34130 27022 34132 27074
rect 34076 27010 34132 27022
rect 33180 26852 33572 26908
rect 33180 26292 33236 26852
rect 33516 26514 33572 26852
rect 33516 26462 33518 26514
rect 33570 26462 33572 26514
rect 33516 26450 33572 26462
rect 33964 26962 34020 26974
rect 33964 26910 33966 26962
rect 34018 26910 34020 26962
rect 33180 26226 33236 26236
rect 33516 26180 33572 26190
rect 32956 25554 33012 25564
rect 33292 25844 33348 25854
rect 32844 25342 32846 25394
rect 32898 25342 32900 25394
rect 32508 25282 32564 25294
rect 32508 25230 32510 25282
rect 32562 25230 32564 25282
rect 31948 24724 32004 24734
rect 31612 24722 32004 24724
rect 31612 24670 31950 24722
rect 32002 24670 32004 24722
rect 31612 24668 32004 24670
rect 30828 24612 30884 24622
rect 30828 24610 30996 24612
rect 30828 24558 30830 24610
rect 30882 24558 30996 24610
rect 30828 24556 30996 24558
rect 30828 24546 30884 24556
rect 30940 23716 30996 24556
rect 31052 23716 31108 23726
rect 30940 23660 31052 23716
rect 30716 22866 30772 22876
rect 30828 23604 30884 23614
rect 30716 22146 30772 22158
rect 30716 22094 30718 22146
rect 30770 22094 30772 22146
rect 30716 22036 30772 22094
rect 30716 21970 30772 21980
rect 30716 21812 30772 21822
rect 30828 21812 30884 23548
rect 31052 23378 31108 23660
rect 31612 23604 31668 24668
rect 31948 24658 32004 24668
rect 31836 24498 31892 24510
rect 31836 24446 31838 24498
rect 31890 24446 31892 24498
rect 31612 23538 31668 23548
rect 31724 23938 31780 23950
rect 31724 23886 31726 23938
rect 31778 23886 31780 23938
rect 31052 23326 31054 23378
rect 31106 23326 31108 23378
rect 31052 23314 31108 23326
rect 31724 23268 31780 23886
rect 31836 23716 31892 24446
rect 32396 24498 32452 24510
rect 32396 24446 32398 24498
rect 32450 24446 32452 24498
rect 32172 24052 32228 24062
rect 32172 23958 32228 23996
rect 31836 23650 31892 23660
rect 31724 23202 31780 23212
rect 31388 23154 31444 23166
rect 31388 23102 31390 23154
rect 31442 23102 31444 23154
rect 31388 23044 31444 23102
rect 31836 23044 31892 23054
rect 31388 23042 31892 23044
rect 31388 22990 31838 23042
rect 31890 22990 31892 23042
rect 31388 22988 31892 22990
rect 31724 22820 31780 22830
rect 31612 22708 31668 22718
rect 30716 21810 30884 21812
rect 30716 21758 30718 21810
rect 30770 21758 30884 21810
rect 30716 21756 30884 21758
rect 30716 21746 30772 21756
rect 30604 21646 30606 21698
rect 30658 21646 30660 21698
rect 30604 21252 30660 21646
rect 30604 21186 30660 21196
rect 30828 21140 30884 21756
rect 31388 22258 31444 22270
rect 31388 22206 31390 22258
rect 31442 22206 31444 22258
rect 31388 22148 31444 22206
rect 30940 21700 30996 21710
rect 30940 21606 30996 21644
rect 31388 21586 31444 22092
rect 31388 21534 31390 21586
rect 31442 21534 31444 21586
rect 31388 21522 31444 21534
rect 31612 21588 31668 22652
rect 31724 22258 31780 22764
rect 31724 22206 31726 22258
rect 31778 22206 31780 22258
rect 31724 22036 31780 22206
rect 31724 21970 31780 21980
rect 31724 21588 31780 21598
rect 31612 21586 31780 21588
rect 31612 21534 31726 21586
rect 31778 21534 31780 21586
rect 31612 21532 31780 21534
rect 31724 21522 31780 21532
rect 30828 21084 31220 21140
rect 30492 20972 30996 21028
rect 30716 20804 30772 20814
rect 30604 20244 30660 20254
rect 30716 20244 30772 20748
rect 30604 20242 30772 20244
rect 30604 20190 30606 20242
rect 30658 20190 30772 20242
rect 30604 20188 30772 20190
rect 30604 20178 30660 20188
rect 30716 20020 30772 20030
rect 30716 19926 30772 19964
rect 30828 20018 30884 20030
rect 30828 19966 30830 20018
rect 30882 19966 30884 20018
rect 30380 19740 30772 19796
rect 30380 19684 30436 19740
rect 30380 19618 30436 19628
rect 30156 19058 30212 19068
rect 30604 19124 30660 19134
rect 29148 15250 29204 15260
rect 29596 15540 29652 15550
rect 29148 15090 29204 15102
rect 29148 15038 29150 15090
rect 29202 15038 29204 15090
rect 29148 13634 29204 15038
rect 29596 15092 29652 15484
rect 30044 15538 30100 15596
rect 30380 18338 30436 18350
rect 30380 18286 30382 18338
rect 30434 18286 30436 18338
rect 30380 17556 30436 18286
rect 30380 15652 30436 17500
rect 30492 18116 30548 18126
rect 30492 17442 30548 18060
rect 30492 17390 30494 17442
rect 30546 17390 30548 17442
rect 30492 17378 30548 17390
rect 30604 17890 30660 19068
rect 30716 18450 30772 19740
rect 30828 19458 30884 19966
rect 30828 19406 30830 19458
rect 30882 19406 30884 19458
rect 30828 19394 30884 19406
rect 30828 19124 30884 19134
rect 30828 19030 30884 19068
rect 30716 18398 30718 18450
rect 30770 18398 30772 18450
rect 30716 18226 30772 18398
rect 30716 18174 30718 18226
rect 30770 18174 30772 18226
rect 30716 18162 30772 18174
rect 30604 17838 30606 17890
rect 30658 17838 30660 17890
rect 30492 17108 30548 17118
rect 30604 17108 30660 17838
rect 30828 17892 30884 17902
rect 30828 17798 30884 17836
rect 30492 17106 30660 17108
rect 30492 17054 30494 17106
rect 30546 17054 30660 17106
rect 30492 17052 30660 17054
rect 30828 17332 30884 17342
rect 30492 17042 30548 17052
rect 30828 16884 30884 17276
rect 30828 16790 30884 16828
rect 30380 15586 30436 15596
rect 30044 15486 30046 15538
rect 30098 15486 30100 15538
rect 30044 15474 30100 15486
rect 29596 15026 29652 15036
rect 30380 15316 30436 15326
rect 29484 14532 29540 14542
rect 29484 14438 29540 14476
rect 29820 14418 29876 14430
rect 29820 14366 29822 14418
rect 29874 14366 29876 14418
rect 29708 14306 29764 14318
rect 29708 14254 29710 14306
rect 29762 14254 29764 14306
rect 29148 13582 29150 13634
rect 29202 13582 29204 13634
rect 29148 13570 29204 13582
rect 29260 13746 29316 13758
rect 29260 13694 29262 13746
rect 29314 13694 29316 13746
rect 29260 13636 29316 13694
rect 29260 13570 29316 13580
rect 29708 13524 29764 14254
rect 29596 13076 29652 13086
rect 29596 12982 29652 13020
rect 29708 12964 29764 13468
rect 29820 14308 29876 14366
rect 29820 13188 29876 14252
rect 30268 14308 30324 14318
rect 30268 14214 30324 14252
rect 30268 13748 30324 13758
rect 30268 13654 30324 13692
rect 29932 13188 29988 13198
rect 29820 13186 29988 13188
rect 29820 13134 29934 13186
rect 29986 13134 29988 13186
rect 29820 13132 29988 13134
rect 29932 13122 29988 13132
rect 29708 12898 29764 12908
rect 29260 12740 29316 12750
rect 29260 12402 29316 12684
rect 29708 12740 29764 12750
rect 29708 12646 29764 12684
rect 29260 12350 29262 12402
rect 29314 12350 29316 12402
rect 29260 12338 29316 12350
rect 30380 12402 30436 15260
rect 30940 14868 30996 20972
rect 31052 20916 31108 20926
rect 31052 20822 31108 20860
rect 31164 20580 31220 21084
rect 31276 20916 31332 20926
rect 31276 20822 31332 20860
rect 31836 20804 31892 22988
rect 32396 23042 32452 24446
rect 32508 24276 32564 25230
rect 32732 24946 32788 24958
rect 32732 24894 32734 24946
rect 32786 24894 32788 24946
rect 32732 24724 32788 24894
rect 32732 24658 32788 24668
rect 32844 24612 32900 25342
rect 32956 24612 33012 24622
rect 32844 24556 32956 24612
rect 32956 24546 33012 24556
rect 32620 24500 32676 24510
rect 32620 24498 32900 24500
rect 32620 24446 32622 24498
rect 32674 24446 32900 24498
rect 32620 24444 32900 24446
rect 32620 24434 32676 24444
rect 32508 24220 32788 24276
rect 32732 23938 32788 24220
rect 32732 23886 32734 23938
rect 32786 23886 32788 23938
rect 32732 23874 32788 23886
rect 32396 22990 32398 23042
rect 32450 22990 32452 23042
rect 32172 22932 32228 22942
rect 32172 22482 32228 22876
rect 32396 22594 32452 22990
rect 32396 22542 32398 22594
rect 32450 22542 32452 22594
rect 32396 22530 32452 22542
rect 32844 23042 32900 24444
rect 32844 22990 32846 23042
rect 32898 22990 32900 23042
rect 32172 22430 32174 22482
rect 32226 22430 32228 22482
rect 32172 22372 32228 22430
rect 32172 22306 32228 22316
rect 32732 22148 32788 22158
rect 32508 22146 32788 22148
rect 32508 22094 32734 22146
rect 32786 22094 32788 22146
rect 32508 22092 32788 22094
rect 31948 21700 32004 21710
rect 31948 21606 32004 21644
rect 32172 21588 32228 21598
rect 32508 21588 32564 22092
rect 32732 22082 32788 22092
rect 32844 21924 32900 22990
rect 32060 21586 32564 21588
rect 32060 21534 32174 21586
rect 32226 21534 32564 21586
rect 32060 21532 32564 21534
rect 32732 21868 32900 21924
rect 32956 24050 33012 24062
rect 32956 23998 32958 24050
rect 33010 23998 33012 24050
rect 31164 20514 31220 20524
rect 31724 20748 31892 20804
rect 31948 21474 32004 21486
rect 31948 21422 31950 21474
rect 32002 21422 32004 21474
rect 30940 14802 30996 14812
rect 31052 20130 31108 20142
rect 31052 20078 31054 20130
rect 31106 20078 31108 20130
rect 31052 19348 31108 20078
rect 31724 20020 31780 20748
rect 31836 20580 31892 20590
rect 31836 20242 31892 20524
rect 31836 20190 31838 20242
rect 31890 20190 31892 20242
rect 31836 20178 31892 20190
rect 31724 19964 31892 20020
rect 31724 19794 31780 19806
rect 31724 19742 31726 19794
rect 31778 19742 31780 19794
rect 31052 14644 31108 19292
rect 31164 19458 31220 19470
rect 31612 19460 31668 19470
rect 31724 19460 31780 19742
rect 31164 19406 31166 19458
rect 31218 19406 31220 19458
rect 31164 17892 31220 19406
rect 31500 19458 31780 19460
rect 31500 19406 31614 19458
rect 31666 19406 31780 19458
rect 31500 19404 31780 19406
rect 31164 17826 31220 17836
rect 31276 19236 31332 19246
rect 31164 17554 31220 17566
rect 31164 17502 31166 17554
rect 31218 17502 31220 17554
rect 31164 17220 31220 17502
rect 31276 17332 31332 19180
rect 31388 19124 31444 19134
rect 31388 19030 31444 19068
rect 31388 18676 31444 18686
rect 31500 18676 31556 19404
rect 31612 19394 31668 19404
rect 31836 19348 31892 19964
rect 31836 19282 31892 19292
rect 31948 19236 32004 21422
rect 31948 19170 32004 19180
rect 32060 19794 32116 21532
rect 32172 21522 32228 21532
rect 32620 21474 32676 21486
rect 32620 21422 32622 21474
rect 32674 21422 32676 21474
rect 32620 21252 32676 21422
rect 32620 21186 32676 21196
rect 32172 21028 32228 21038
rect 32172 20802 32228 20972
rect 32620 21028 32676 21038
rect 32620 20914 32676 20972
rect 32620 20862 32622 20914
rect 32674 20862 32676 20914
rect 32620 20850 32676 20862
rect 32172 20750 32174 20802
rect 32226 20750 32228 20802
rect 32172 20738 32228 20750
rect 32060 19742 32062 19794
rect 32114 19742 32116 19794
rect 31388 18674 31556 18676
rect 31388 18622 31390 18674
rect 31442 18622 31556 18674
rect 31388 18620 31556 18622
rect 31724 19012 31780 19022
rect 31388 18610 31444 18620
rect 31612 18564 31668 18574
rect 31612 18470 31668 18508
rect 31500 18338 31556 18350
rect 31500 18286 31502 18338
rect 31554 18286 31556 18338
rect 31500 17780 31556 18286
rect 31500 17714 31556 17724
rect 31388 17556 31444 17566
rect 31724 17556 31780 18956
rect 31948 19010 32004 19022
rect 31948 18958 31950 19010
rect 32002 18958 32004 19010
rect 31948 18452 32004 18958
rect 32060 18676 32116 19742
rect 32508 19906 32564 19918
rect 32508 19854 32510 19906
rect 32562 19854 32564 19906
rect 32396 19348 32452 19358
rect 32396 19254 32452 19292
rect 32060 18620 32340 18676
rect 31948 18386 32004 18396
rect 32060 18452 32116 18462
rect 32060 18450 32228 18452
rect 32060 18398 32062 18450
rect 32114 18398 32228 18450
rect 32060 18396 32228 18398
rect 32060 18386 32116 18396
rect 31388 17554 31780 17556
rect 31388 17502 31390 17554
rect 31442 17502 31780 17554
rect 31388 17500 31780 17502
rect 31836 18340 31892 18350
rect 31388 17490 31444 17500
rect 31276 17276 31444 17332
rect 31164 17154 31220 17164
rect 31276 17108 31332 17118
rect 31276 17014 31332 17052
rect 31388 16098 31444 17276
rect 31612 17108 31668 17500
rect 31612 17042 31668 17052
rect 31836 16884 31892 18284
rect 32172 18226 32228 18396
rect 32284 18340 32340 18620
rect 32396 18340 32452 18350
rect 32284 18284 32396 18340
rect 32396 18246 32452 18284
rect 32172 18174 32174 18226
rect 32226 18174 32228 18226
rect 32172 18162 32228 18174
rect 32508 17892 32564 19854
rect 32732 19348 32788 21868
rect 32732 19282 32788 19292
rect 32844 21028 32900 21038
rect 32844 19346 32900 20972
rect 32844 19294 32846 19346
rect 32898 19294 32900 19346
rect 32844 19282 32900 19294
rect 32956 18564 33012 23998
rect 33180 23826 33236 23838
rect 33180 23774 33182 23826
rect 33234 23774 33236 23826
rect 32732 18508 33012 18564
rect 33068 23268 33124 23278
rect 33068 22148 33124 23212
rect 33180 22484 33236 23774
rect 33180 22418 33236 22428
rect 33292 22260 33348 25788
rect 33516 25396 33572 26124
rect 33852 25732 33908 25742
rect 33404 24612 33460 24622
rect 33404 22820 33460 24556
rect 33404 22754 33460 22764
rect 33516 23042 33572 25340
rect 33740 25394 33796 25406
rect 33740 25342 33742 25394
rect 33794 25342 33796 25394
rect 33740 25060 33796 25342
rect 33740 24994 33796 25004
rect 33628 24724 33684 24734
rect 33628 24630 33684 24668
rect 33852 23380 33908 25676
rect 33964 25508 34020 26910
rect 34636 26964 34692 27002
rect 34636 26898 34692 26908
rect 34300 26850 34356 26862
rect 34300 26798 34302 26850
rect 34354 26798 34356 26850
rect 34300 25620 34356 26798
rect 34524 26628 34580 26638
rect 34524 26290 34580 26572
rect 34748 26514 34804 27132
rect 34860 27076 34916 27114
rect 34860 27010 34916 27020
rect 34972 26964 35028 26974
rect 34748 26462 34750 26514
rect 34802 26462 34804 26514
rect 34748 26450 34804 26462
rect 34860 26852 35028 26908
rect 34524 26238 34526 26290
rect 34578 26238 34580 26290
rect 34300 25564 34468 25620
rect 33964 25442 34020 25452
rect 34300 25396 34356 25406
rect 34300 25302 34356 25340
rect 33964 25282 34020 25294
rect 33964 25230 33966 25282
rect 34018 25230 34020 25282
rect 33964 24948 34020 25230
rect 34300 24948 34356 24958
rect 33964 24946 34356 24948
rect 33964 24894 34302 24946
rect 34354 24894 34356 24946
rect 33964 24892 34356 24894
rect 34300 24882 34356 24892
rect 33964 24722 34020 24734
rect 33964 24670 33966 24722
rect 34018 24670 34020 24722
rect 33964 24164 34020 24670
rect 34076 24722 34132 24734
rect 34076 24670 34078 24722
rect 34130 24670 34132 24722
rect 34076 24612 34132 24670
rect 34076 24546 34132 24556
rect 34188 24610 34244 24622
rect 34188 24558 34190 24610
rect 34242 24558 34244 24610
rect 34188 24388 34244 24558
rect 34188 24322 34244 24332
rect 34300 24500 34356 24510
rect 34300 24164 34356 24444
rect 33964 24098 34020 24108
rect 34188 24108 34356 24164
rect 34188 24050 34244 24108
rect 34188 23998 34190 24050
rect 34242 23998 34244 24050
rect 34188 23986 34244 23998
rect 34076 23940 34132 23950
rect 33964 23938 34132 23940
rect 33964 23886 34078 23938
rect 34130 23886 34132 23938
rect 33964 23884 34132 23886
rect 33964 23828 34020 23884
rect 34076 23874 34132 23884
rect 33964 23548 34020 23772
rect 34188 23604 34244 23614
rect 33964 23492 34132 23548
rect 33964 23380 34020 23390
rect 33516 22990 33518 23042
rect 33570 22990 33572 23042
rect 33292 22194 33348 22204
rect 33404 22594 33460 22606
rect 33404 22542 33406 22594
rect 33458 22542 33460 22594
rect 33180 22148 33236 22158
rect 33068 22146 33236 22148
rect 33068 22094 33182 22146
rect 33234 22094 33236 22146
rect 33068 22092 33236 22094
rect 33068 18564 33124 22092
rect 33180 22082 33236 22092
rect 33180 21252 33236 21262
rect 33180 20914 33236 21196
rect 33180 20862 33182 20914
rect 33234 20862 33236 20914
rect 33180 20850 33236 20862
rect 33292 21026 33348 21038
rect 33292 20974 33294 21026
rect 33346 20974 33348 21026
rect 33292 19796 33348 20974
rect 32508 17826 32564 17836
rect 32620 18452 32676 18462
rect 32396 17668 32452 17678
rect 32396 17574 32452 17612
rect 32620 17666 32676 18396
rect 32620 17614 32622 17666
rect 32674 17614 32676 17666
rect 31948 17554 32004 17566
rect 31948 17502 31950 17554
rect 32002 17502 32004 17554
rect 31948 17332 32004 17502
rect 32172 17444 32228 17454
rect 31948 17266 32004 17276
rect 32060 17442 32228 17444
rect 32060 17390 32174 17442
rect 32226 17390 32228 17442
rect 32060 17388 32228 17390
rect 31948 17108 32004 17118
rect 32060 17108 32116 17388
rect 32172 17378 32228 17388
rect 32284 17442 32340 17454
rect 32284 17390 32286 17442
rect 32338 17390 32340 17442
rect 31948 17106 32116 17108
rect 31948 17054 31950 17106
rect 32002 17054 32116 17106
rect 31948 17052 32116 17054
rect 31948 17042 32004 17052
rect 32060 16884 32116 16894
rect 31836 16882 32004 16884
rect 31836 16830 31838 16882
rect 31890 16830 32004 16882
rect 31836 16828 32004 16830
rect 31836 16818 31892 16828
rect 31388 16046 31390 16098
rect 31442 16046 31444 16098
rect 31388 16034 31444 16046
rect 31948 16100 32004 16828
rect 32060 16790 32116 16828
rect 32284 16324 32340 17390
rect 31948 16034 32004 16044
rect 32172 16268 32340 16324
rect 32396 17108 32452 17118
rect 31836 15874 31892 15886
rect 31836 15822 31838 15874
rect 31890 15822 31892 15874
rect 31836 15204 31892 15822
rect 31948 15874 32004 15886
rect 31948 15822 31950 15874
rect 32002 15822 32004 15874
rect 31948 15316 32004 15822
rect 31948 15250 32004 15260
rect 32060 15874 32116 15886
rect 32060 15822 32062 15874
rect 32114 15822 32116 15874
rect 31836 15138 31892 15148
rect 30828 14588 31108 14644
rect 31388 14642 31444 14654
rect 31388 14590 31390 14642
rect 31442 14590 31444 14642
rect 30492 14308 30548 14318
rect 30492 13074 30548 14252
rect 30492 13022 30494 13074
rect 30546 13022 30548 13074
rect 30492 13010 30548 13022
rect 30380 12350 30382 12402
rect 30434 12350 30436 12402
rect 30380 12180 30436 12350
rect 30380 12114 30436 12124
rect 29932 12068 29988 12078
rect 29932 11974 29988 12012
rect 30492 12068 30548 12078
rect 29036 11618 29652 11620
rect 29036 11566 29038 11618
rect 29090 11566 29652 11618
rect 29036 11564 29652 11566
rect 29036 11554 29092 11564
rect 29596 11394 29652 11564
rect 29596 11342 29598 11394
rect 29650 11342 29652 11394
rect 29596 11330 29652 11342
rect 29932 11282 29988 11294
rect 29932 11230 29934 11282
rect 29986 11230 29988 11282
rect 29820 11170 29876 11182
rect 29820 11118 29822 11170
rect 29874 11118 29876 11170
rect 28924 10446 28926 10498
rect 28978 10446 28980 10498
rect 28924 10434 28980 10446
rect 29148 10610 29204 10622
rect 29148 10558 29150 10610
rect 29202 10558 29204 10610
rect 28812 9886 28814 9938
rect 28866 9886 28868 9938
rect 27804 9436 28196 9492
rect 28028 9156 28084 9166
rect 27692 9100 27972 9156
rect 27468 8876 27636 8932
rect 27468 8260 27524 8876
rect 27356 8148 27412 8158
rect 27468 8148 27524 8204
rect 27692 8148 27748 8158
rect 27468 8146 27748 8148
rect 27468 8094 27694 8146
rect 27746 8094 27748 8146
rect 27468 8092 27748 8094
rect 27356 6356 27412 8092
rect 27692 8082 27748 8092
rect 27804 8148 27860 8158
rect 27804 8054 27860 8092
rect 27468 7364 27524 7374
rect 27468 7270 27524 7308
rect 27468 6692 27524 6702
rect 27468 6598 27524 6636
rect 27356 6300 27636 6356
rect 27244 6188 27412 6244
rect 27244 6020 27300 6030
rect 27132 6018 27300 6020
rect 27132 5966 27246 6018
rect 27298 5966 27300 6018
rect 27132 5964 27300 5966
rect 27244 5954 27300 5964
rect 26348 4452 26404 4462
rect 26348 4358 26404 4396
rect 26684 4340 26740 4350
rect 26684 4246 26740 4284
rect 25564 4162 25620 4172
rect 26796 3556 26852 3566
rect 26796 3462 26852 3500
rect 27356 3556 27412 6188
rect 27580 6130 27636 6300
rect 27580 6078 27582 6130
rect 27634 6078 27636 6130
rect 27580 6066 27636 6078
rect 27356 3490 27412 3500
rect 27580 3666 27636 3678
rect 27580 3614 27582 3666
rect 27634 3614 27636 3666
rect 23884 2706 23940 2716
rect 27580 800 27636 3614
rect 27916 3108 27972 9100
rect 28028 8258 28084 9100
rect 28028 8206 28030 8258
rect 28082 8206 28084 8258
rect 28028 8194 28084 8206
rect 28140 7812 28196 9436
rect 28812 9268 28868 9886
rect 29148 9716 29204 10558
rect 29372 10610 29428 10622
rect 29372 10558 29374 10610
rect 29426 10558 29428 10610
rect 29372 10500 29428 10558
rect 29820 10500 29876 11118
rect 29932 10724 29988 11230
rect 29932 10658 29988 10668
rect 30380 11284 30436 11294
rect 29372 10444 30100 10500
rect 29484 9828 29540 9838
rect 29820 9828 29876 9838
rect 29484 9734 29540 9772
rect 29708 9826 29876 9828
rect 29708 9774 29822 9826
rect 29874 9774 29876 9826
rect 29708 9772 29876 9774
rect 29148 9650 29204 9660
rect 29036 9268 29092 9278
rect 29708 9268 29764 9772
rect 29820 9762 29876 9772
rect 30044 9826 30100 10444
rect 30044 9774 30046 9826
rect 30098 9774 30100 9826
rect 30044 9762 30100 9774
rect 29820 9602 29876 9614
rect 29820 9550 29822 9602
rect 29874 9550 29876 9602
rect 29820 9492 29876 9550
rect 29820 9436 30100 9492
rect 28812 9266 29876 9268
rect 28812 9214 29038 9266
rect 29090 9214 29876 9266
rect 28812 9212 29876 9214
rect 29036 9202 29092 9212
rect 29820 9154 29876 9212
rect 29820 9102 29822 9154
rect 29874 9102 29876 9154
rect 29820 9090 29876 9102
rect 29820 8484 29876 8494
rect 28028 7756 28196 7812
rect 28476 8148 28532 8158
rect 28476 8034 28532 8092
rect 28476 7982 28478 8034
rect 28530 7982 28532 8034
rect 28476 7812 28532 7982
rect 28028 6692 28084 7756
rect 28476 7746 28532 7756
rect 29596 8146 29652 8158
rect 29596 8094 29598 8146
rect 29650 8094 29652 8146
rect 28476 7588 28532 7598
rect 28476 7494 28532 7532
rect 29372 7588 29428 7598
rect 29596 7588 29652 8094
rect 29372 7586 29652 7588
rect 29372 7534 29374 7586
rect 29426 7534 29652 7586
rect 29372 7532 29652 7534
rect 29372 7522 29428 7532
rect 28140 7476 28196 7486
rect 28140 7382 28196 7420
rect 28700 7476 28756 7486
rect 28028 6560 28084 6636
rect 28252 7362 28308 7374
rect 28252 7310 28254 7362
rect 28306 7310 28308 7362
rect 28140 6578 28196 6590
rect 28140 6526 28142 6578
rect 28194 6526 28196 6578
rect 28140 6356 28196 6526
rect 28140 6290 28196 6300
rect 28252 6244 28308 7310
rect 28252 6178 28308 6188
rect 28364 7364 28420 7374
rect 28364 6020 28420 7308
rect 28700 6802 28756 7420
rect 29036 7476 29092 7514
rect 29036 7410 29092 7420
rect 29820 7476 29876 8428
rect 30044 8258 30100 9436
rect 30156 9044 30212 9054
rect 30156 8950 30212 8988
rect 30044 8206 30046 8258
rect 30098 8206 30100 8258
rect 30044 7588 30100 8206
rect 30044 7522 30100 7532
rect 29820 7362 29876 7420
rect 29820 7310 29822 7362
rect 29874 7310 29876 7362
rect 29036 7250 29092 7262
rect 29036 7198 29038 7250
rect 29090 7198 29092 7250
rect 29036 7140 29092 7198
rect 29036 7074 29092 7084
rect 28700 6750 28702 6802
rect 28754 6750 28756 6802
rect 28700 6738 28756 6750
rect 29484 6466 29540 6478
rect 29484 6414 29486 6466
rect 29538 6414 29540 6466
rect 29484 6356 29540 6414
rect 29484 6290 29540 6300
rect 29820 6244 29876 7310
rect 29820 6178 29876 6188
rect 28028 5964 28420 6020
rect 28028 5234 28084 5964
rect 28364 5906 28420 5964
rect 28364 5854 28366 5906
rect 28418 5854 28420 5906
rect 28364 5842 28420 5854
rect 28028 5182 28030 5234
rect 28082 5182 28084 5234
rect 28028 5170 28084 5182
rect 28140 5794 28196 5806
rect 28140 5742 28142 5794
rect 28194 5742 28196 5794
rect 28140 5236 28196 5742
rect 28700 5684 28756 5694
rect 28476 5682 28756 5684
rect 28476 5630 28702 5682
rect 28754 5630 28756 5682
rect 28476 5628 28756 5630
rect 28364 5236 28420 5246
rect 28140 5180 28364 5236
rect 28364 5122 28420 5180
rect 28364 5070 28366 5122
rect 28418 5070 28420 5122
rect 28364 5058 28420 5070
rect 28476 4338 28532 5628
rect 28700 5618 28756 5628
rect 28476 4286 28478 4338
rect 28530 4286 28532 4338
rect 28476 4274 28532 4286
rect 28812 5010 28868 5022
rect 28812 4958 28814 5010
rect 28866 4958 28868 5010
rect 28588 4228 28644 4238
rect 28812 4228 28868 4958
rect 29372 4564 29428 4574
rect 29372 4338 29428 4508
rect 29372 4286 29374 4338
rect 29426 4286 29428 4338
rect 29372 4274 29428 4286
rect 29820 4564 29876 4574
rect 28924 4228 28980 4238
rect 28812 4226 28980 4228
rect 28812 4174 28926 4226
rect 28978 4174 28980 4226
rect 28812 4172 28980 4174
rect 28588 4134 28644 4172
rect 28924 4116 28980 4172
rect 28924 4060 29428 4116
rect 29372 3666 29428 4060
rect 29372 3614 29374 3666
rect 29426 3614 29428 3666
rect 29372 3602 29428 3614
rect 27916 3042 27972 3052
rect 28476 3556 28532 3566
rect 28476 1652 28532 3500
rect 29820 3554 29876 4508
rect 30268 4338 30324 4350
rect 30268 4286 30270 4338
rect 30322 4286 30324 4338
rect 30268 3666 30324 4286
rect 30268 3614 30270 3666
rect 30322 3614 30324 3666
rect 30268 3602 30324 3614
rect 29820 3502 29822 3554
rect 29874 3502 29876 3554
rect 29820 3490 29876 3502
rect 30380 3556 30436 11228
rect 30492 11172 30548 12012
rect 30828 11788 30884 14588
rect 31052 14420 31108 14430
rect 31052 14326 31108 14364
rect 31388 13970 31444 14590
rect 32060 14644 32116 15822
rect 32060 14578 32116 14588
rect 31948 14532 32004 14542
rect 31948 14438 32004 14476
rect 31388 13918 31390 13970
rect 31442 13918 31444 13970
rect 31388 13906 31444 13918
rect 31276 13858 31332 13870
rect 31276 13806 31278 13858
rect 31330 13806 31332 13858
rect 30940 12740 30996 12750
rect 30940 11956 30996 12684
rect 31164 12516 31220 12526
rect 31164 12402 31220 12460
rect 31164 12350 31166 12402
rect 31218 12350 31220 12402
rect 31164 12338 31220 12350
rect 31276 12404 31332 13806
rect 31500 13524 31556 13534
rect 31500 13076 31556 13468
rect 31836 13412 31892 13422
rect 31612 13076 31668 13086
rect 31836 13076 31892 13356
rect 31500 13074 31668 13076
rect 31500 13022 31614 13074
rect 31666 13022 31668 13074
rect 31500 13020 31668 13022
rect 31612 13010 31668 13020
rect 31724 13020 32004 13076
rect 31500 12852 31556 12862
rect 31276 12348 31444 12404
rect 31052 12178 31108 12190
rect 31052 12126 31054 12178
rect 31106 12126 31108 12178
rect 31052 12068 31108 12126
rect 31276 12180 31332 12190
rect 31276 12086 31332 12124
rect 31052 12002 31108 12012
rect 30940 11890 30996 11900
rect 30716 11732 30884 11788
rect 30604 11396 30660 11406
rect 30604 11302 30660 11340
rect 30492 11106 30548 11116
rect 30492 10724 30548 10734
rect 30492 10630 30548 10668
rect 30604 9716 30660 9726
rect 30604 9602 30660 9660
rect 30604 9550 30606 9602
rect 30658 9550 30660 9602
rect 30604 8484 30660 9550
rect 30604 8418 30660 8428
rect 30492 8372 30548 8382
rect 30492 8278 30548 8316
rect 30716 8148 30772 11732
rect 31388 11618 31444 12348
rect 31500 12178 31556 12796
rect 31500 12126 31502 12178
rect 31554 12126 31556 12178
rect 31500 12114 31556 12126
rect 31388 11566 31390 11618
rect 31442 11566 31444 11618
rect 31052 11396 31108 11406
rect 31052 11302 31108 11340
rect 31276 11172 31332 11182
rect 31276 11078 31332 11116
rect 31164 10612 31220 10622
rect 31164 10518 31220 10556
rect 31388 10610 31444 11566
rect 31724 11172 31780 13020
rect 31948 12962 32004 13020
rect 31948 12910 31950 12962
rect 32002 12910 32004 12962
rect 31948 12898 32004 12910
rect 31836 12850 31892 12862
rect 31836 12798 31838 12850
rect 31890 12798 31892 12850
rect 31836 12404 31892 12798
rect 32172 12516 32228 16268
rect 32396 16100 32452 17052
rect 32620 16996 32676 17614
rect 32620 16930 32676 16940
rect 32508 16882 32564 16894
rect 32508 16830 32510 16882
rect 32562 16830 32564 16882
rect 32508 16660 32564 16830
rect 32508 16594 32564 16604
rect 32508 16100 32564 16110
rect 32732 16100 32788 18508
rect 33068 18498 33124 18508
rect 33180 19740 33348 19796
rect 32844 18340 32900 18350
rect 32844 18338 33124 18340
rect 32844 18286 32846 18338
rect 32898 18286 33124 18338
rect 32844 18284 33124 18286
rect 32844 18226 32900 18284
rect 32844 18174 32846 18226
rect 32898 18174 32900 18226
rect 32844 18162 32900 18174
rect 32956 17892 33012 17902
rect 32956 17106 33012 17836
rect 32956 17054 32958 17106
rect 33010 17054 33012 17106
rect 32956 17042 33012 17054
rect 32396 16098 32564 16100
rect 32396 16046 32510 16098
rect 32562 16046 32564 16098
rect 32396 16044 32564 16046
rect 32508 16034 32564 16044
rect 32620 16044 32788 16100
rect 32620 15540 32676 16044
rect 32844 15986 32900 15998
rect 32844 15934 32846 15986
rect 32898 15934 32900 15986
rect 32732 15876 32788 15886
rect 32732 15782 32788 15820
rect 32620 15474 32676 15484
rect 32284 15204 32340 15242
rect 32284 15138 32340 15148
rect 32732 15202 32788 15214
rect 32732 15150 32734 15202
rect 32786 15150 32788 15202
rect 32732 14644 32788 15150
rect 32844 15204 32900 15934
rect 32844 15138 32900 15148
rect 32732 14578 32788 14588
rect 32732 14308 32788 14318
rect 32396 13634 32452 13646
rect 32396 13582 32398 13634
rect 32450 13582 32452 13634
rect 32396 13412 32452 13582
rect 32396 13346 32452 13356
rect 32620 12852 32676 12862
rect 32620 12758 32676 12796
rect 32172 12460 32340 12516
rect 31836 12348 32004 12404
rect 31948 12292 32004 12348
rect 31948 12236 32228 12292
rect 31836 12180 31892 12190
rect 31836 12086 31892 12124
rect 31724 11106 31780 11116
rect 31836 11732 31892 11742
rect 31388 10558 31390 10610
rect 31442 10558 31444 10610
rect 31388 9154 31444 10558
rect 31388 9102 31390 9154
rect 31442 9102 31444 9154
rect 31388 9090 31444 9102
rect 31612 9266 31668 9278
rect 31612 9214 31614 9266
rect 31666 9214 31668 9266
rect 31164 8372 31220 8382
rect 31164 8278 31220 8316
rect 30604 8092 30772 8148
rect 30492 6466 30548 6478
rect 30492 6414 30494 6466
rect 30546 6414 30548 6466
rect 30492 5796 30548 6414
rect 30604 6020 30660 8092
rect 30940 7812 30996 7822
rect 30940 7364 30996 7756
rect 30940 7270 30996 7308
rect 31612 7698 31668 9214
rect 31836 8820 31892 11676
rect 32060 11620 32116 11630
rect 32060 11506 32116 11564
rect 32060 11454 32062 11506
rect 32114 11454 32116 11506
rect 32060 11442 32116 11454
rect 31948 11396 32004 11406
rect 31948 11302 32004 11340
rect 32172 11284 32228 12236
rect 32060 11228 32172 11284
rect 32060 10722 32116 11228
rect 32172 11152 32228 11228
rect 32060 10670 32062 10722
rect 32114 10670 32116 10722
rect 32060 10612 32116 10670
rect 32060 10546 32116 10556
rect 31836 8754 31892 8764
rect 32172 10050 32228 10062
rect 32172 9998 32174 10050
rect 32226 9998 32228 10050
rect 32172 9044 32228 9998
rect 32172 8930 32228 8988
rect 32172 8878 32174 8930
rect 32226 8878 32228 8930
rect 32172 7812 32228 8878
rect 32284 8372 32340 12460
rect 32620 12290 32676 12302
rect 32620 12238 32622 12290
rect 32674 12238 32676 12290
rect 32508 12180 32564 12190
rect 32508 12086 32564 12124
rect 32396 11954 32452 11966
rect 32396 11902 32398 11954
rect 32450 11902 32452 11954
rect 32396 11284 32452 11902
rect 32620 11956 32676 12238
rect 32508 11844 32564 11854
rect 32508 11618 32564 11788
rect 32508 11566 32510 11618
rect 32562 11566 32564 11618
rect 32508 11554 32564 11566
rect 32620 11394 32676 11900
rect 32620 11342 32622 11394
rect 32674 11342 32676 11394
rect 32620 11330 32676 11342
rect 32396 11218 32452 11228
rect 32396 10610 32452 10622
rect 32396 10558 32398 10610
rect 32450 10558 32452 10610
rect 32396 10050 32452 10558
rect 32396 9998 32398 10050
rect 32450 9998 32452 10050
rect 32396 9986 32452 9998
rect 32508 9602 32564 9614
rect 32508 9550 32510 9602
rect 32562 9550 32564 9602
rect 32508 9268 32564 9550
rect 32508 9202 32564 9212
rect 32284 8306 32340 8316
rect 32172 7746 32228 7756
rect 31612 7646 31614 7698
rect 31666 7646 31668 7698
rect 31276 7252 31332 7262
rect 30828 6692 30884 6702
rect 30828 6598 30884 6636
rect 30716 6580 30772 6590
rect 30716 6486 30772 6524
rect 31164 6132 31220 6142
rect 30604 5964 30884 6020
rect 30716 5796 30772 5806
rect 30492 5794 30772 5796
rect 30492 5742 30718 5794
rect 30770 5742 30772 5794
rect 30492 5740 30772 5742
rect 30716 5730 30772 5740
rect 30604 4452 30660 4462
rect 30604 4358 30660 4396
rect 30380 3490 30436 3500
rect 30828 3388 30884 5964
rect 31164 6018 31220 6076
rect 31164 5966 31166 6018
rect 31218 5966 31220 6018
rect 31164 5954 31220 5966
rect 31164 5236 31220 5246
rect 31164 5142 31220 5180
rect 31276 5010 31332 7196
rect 31388 6690 31444 6702
rect 31388 6638 31390 6690
rect 31442 6638 31444 6690
rect 31388 6580 31444 6638
rect 31612 6692 31668 7646
rect 31724 7474 31780 7486
rect 31724 7422 31726 7474
rect 31778 7422 31780 7474
rect 31724 7364 31780 7422
rect 31948 7474 32004 7486
rect 31948 7422 31950 7474
rect 32002 7422 32004 7474
rect 31724 7298 31780 7308
rect 31836 7362 31892 7374
rect 31836 7310 31838 7362
rect 31890 7310 31892 7362
rect 31612 6560 31668 6636
rect 31836 6692 31892 7310
rect 31836 6626 31892 6636
rect 31724 6578 31780 6590
rect 31388 6514 31444 6524
rect 31724 6526 31726 6578
rect 31778 6526 31780 6578
rect 31724 6468 31780 6526
rect 31948 6468 32004 7422
rect 31724 6412 32004 6468
rect 32172 7474 32228 7486
rect 32172 7422 32174 7474
rect 32226 7422 32228 7474
rect 32172 6690 32228 7422
rect 32172 6638 32174 6690
rect 32226 6638 32228 6690
rect 31724 5796 31780 6412
rect 32172 5908 32228 6638
rect 32172 5842 32228 5852
rect 32396 6468 32452 6478
rect 31724 5730 31780 5740
rect 31500 5348 31556 5358
rect 31500 5254 31556 5292
rect 32396 5348 32452 6412
rect 32396 5282 32452 5292
rect 32508 6130 32564 6142
rect 32508 6078 32510 6130
rect 32562 6078 32564 6130
rect 32508 5122 32564 6078
rect 32620 6020 32676 6030
rect 32620 5926 32676 5964
rect 32508 5070 32510 5122
rect 32562 5070 32564 5122
rect 31276 4958 31278 5010
rect 31330 4958 31332 5010
rect 31276 4946 31332 4958
rect 32396 5010 32452 5022
rect 32396 4958 32398 5010
rect 32450 4958 32452 5010
rect 32396 4676 32452 4958
rect 31836 4340 31892 4350
rect 31836 4246 31892 4284
rect 32396 4338 32452 4620
rect 32396 4286 32398 4338
rect 32450 4286 32452 4338
rect 32396 4274 32452 4286
rect 32508 4228 32564 5070
rect 32620 4228 32676 4238
rect 32508 4226 32676 4228
rect 32508 4174 32622 4226
rect 32674 4174 32676 4226
rect 32508 4172 32676 4174
rect 32620 4162 32676 4172
rect 30828 3332 30996 3388
rect 30940 2996 30996 3332
rect 30940 2930 30996 2940
rect 32732 2884 32788 14252
rect 32956 12964 33012 12974
rect 32956 12870 33012 12908
rect 32844 10498 32900 10510
rect 32844 10446 32846 10498
rect 32898 10446 32900 10498
rect 32844 10050 32900 10446
rect 32844 9998 32846 10050
rect 32898 9998 32900 10050
rect 32844 9986 32900 9998
rect 33068 9828 33124 18284
rect 33180 16884 33236 19740
rect 33292 19010 33348 19022
rect 33292 18958 33294 19010
rect 33346 18958 33348 19010
rect 33292 17332 33348 18958
rect 33404 18676 33460 22542
rect 33516 22372 33572 22990
rect 33516 22306 33572 22316
rect 33628 23378 34020 23380
rect 33628 23326 33966 23378
rect 34018 23326 34020 23378
rect 33628 23324 34020 23326
rect 33516 22148 33572 22158
rect 33516 21026 33572 22092
rect 33628 21364 33684 23324
rect 33964 23314 34020 23324
rect 33740 23044 33796 23054
rect 33740 22370 33796 22988
rect 34076 22484 34132 23492
rect 33740 22318 33742 22370
rect 33794 22318 33796 22370
rect 33740 22306 33796 22318
rect 33964 22428 34132 22484
rect 33852 22146 33908 22158
rect 33852 22094 33854 22146
rect 33906 22094 33908 22146
rect 33740 21812 33796 21822
rect 33740 21586 33796 21756
rect 33740 21534 33742 21586
rect 33794 21534 33796 21586
rect 33740 21522 33796 21534
rect 33684 21308 33796 21364
rect 33628 21298 33684 21308
rect 33516 20974 33518 21026
rect 33570 20974 33572 21026
rect 33516 20914 33572 20974
rect 33516 20862 33518 20914
rect 33570 20862 33572 20914
rect 33516 20850 33572 20862
rect 33404 18610 33460 18620
rect 33516 19908 33572 19918
rect 33516 19124 33572 19852
rect 33628 19236 33684 19246
rect 33628 19142 33684 19180
rect 33516 18674 33572 19068
rect 33516 18622 33518 18674
rect 33570 18622 33572 18674
rect 33516 18610 33572 18622
rect 33740 18228 33796 21308
rect 33516 18172 33796 18228
rect 33516 17666 33572 18172
rect 33516 17614 33518 17666
rect 33570 17614 33572 17666
rect 33292 17266 33348 17276
rect 33404 17442 33460 17454
rect 33404 17390 33406 17442
rect 33458 17390 33460 17442
rect 33404 17108 33460 17390
rect 33404 17042 33460 17052
rect 33180 16212 33236 16828
rect 33516 16322 33572 17614
rect 33852 17666 33908 22094
rect 33964 21588 34020 22428
rect 34076 22260 34132 22270
rect 34076 22166 34132 22204
rect 34076 21810 34132 21822
rect 34076 21758 34078 21810
rect 34130 21758 34132 21810
rect 34076 21700 34132 21758
rect 34188 21812 34244 23548
rect 34412 22596 34468 25564
rect 34524 25172 34580 26238
rect 34524 25106 34580 25116
rect 34412 22530 34468 22540
rect 34524 24164 34580 24174
rect 34300 22258 34356 22270
rect 34300 22206 34302 22258
rect 34354 22206 34356 22258
rect 34300 21924 34356 22206
rect 34412 22260 34468 22270
rect 34412 22036 34468 22204
rect 34524 22148 34580 24108
rect 34860 23940 34916 26852
rect 35084 25732 35140 27244
rect 35420 26516 35476 26526
rect 35532 26516 35588 28476
rect 35756 27970 35812 27982
rect 35756 27918 35758 27970
rect 35810 27918 35812 27970
rect 35756 27636 35812 27918
rect 35756 27570 35812 27580
rect 35756 27300 35812 27310
rect 35644 27188 35700 27198
rect 35644 26852 35700 27132
rect 35756 27074 35812 27244
rect 35756 27022 35758 27074
rect 35810 27022 35812 27074
rect 35756 27010 35812 27022
rect 35644 26786 35700 26796
rect 35868 26516 35924 28700
rect 35980 28532 36036 28814
rect 36092 28756 36148 28766
rect 36092 28662 36148 28700
rect 35980 28476 36148 28532
rect 35980 27860 36036 27870
rect 35980 27188 36036 27804
rect 35980 27122 36036 27132
rect 35532 26460 35812 26516
rect 35420 26422 35476 26460
rect 35532 26292 35588 26302
rect 35644 26292 35700 26302
rect 35532 26290 35644 26292
rect 35532 26238 35534 26290
rect 35586 26238 35644 26290
rect 35532 26236 35644 26238
rect 35532 26226 35588 26236
rect 35420 26180 35476 26190
rect 35420 26066 35476 26124
rect 35420 26014 35422 26066
rect 35474 26014 35476 26066
rect 35420 26002 35476 26014
rect 35532 26068 35588 26078
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35084 25666 35140 25676
rect 35420 25508 35476 25518
rect 35420 25414 35476 25452
rect 34972 25282 35028 25294
rect 34972 25230 34974 25282
rect 35026 25230 35028 25282
rect 34972 24500 35028 25230
rect 34972 24434 35028 24444
rect 35084 25282 35140 25294
rect 35084 25230 35086 25282
rect 35138 25230 35140 25282
rect 34748 23884 34916 23940
rect 34972 24050 35028 24062
rect 34972 23998 34974 24050
rect 35026 23998 35028 24050
rect 34972 23940 35028 23998
rect 35084 23940 35140 25230
rect 35196 25284 35252 25294
rect 35196 24722 35252 25228
rect 35196 24670 35198 24722
rect 35250 24670 35252 24722
rect 35196 24658 35252 24670
rect 35420 24500 35476 24538
rect 35420 24434 35476 24444
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 23940 35252 23950
rect 35084 23938 35252 23940
rect 35084 23886 35198 23938
rect 35250 23886 35252 23938
rect 35084 23884 35252 23886
rect 34748 23268 34804 23884
rect 34972 23874 35028 23884
rect 35196 23874 35252 23884
rect 35420 23826 35476 23838
rect 35420 23774 35422 23826
rect 35474 23774 35476 23826
rect 34860 23716 34916 23726
rect 34860 23622 34916 23660
rect 34972 23716 35028 23726
rect 34972 23714 35252 23716
rect 34972 23662 34974 23714
rect 35026 23662 35252 23714
rect 34972 23660 35252 23662
rect 34972 23650 35028 23660
rect 34748 23212 34916 23268
rect 34636 23154 34692 23166
rect 34636 23102 34638 23154
rect 34690 23102 34692 23154
rect 34636 23044 34692 23102
rect 34636 22978 34692 22988
rect 34748 23042 34804 23054
rect 34748 22990 34750 23042
rect 34802 22990 34804 23042
rect 34748 22708 34804 22990
rect 34748 22642 34804 22652
rect 34860 22372 34916 23212
rect 34972 23154 35028 23166
rect 34972 23102 34974 23154
rect 35026 23102 35028 23154
rect 34972 22594 35028 23102
rect 34972 22542 34974 22594
rect 35026 22542 35028 22594
rect 34972 22530 35028 22542
rect 35084 23154 35140 23166
rect 35084 23102 35086 23154
rect 35138 23102 35140 23154
rect 35084 22596 35140 23102
rect 35196 22932 35252 23660
rect 35420 23604 35476 23774
rect 35420 23538 35476 23548
rect 35532 23492 35588 26012
rect 35644 25730 35700 26236
rect 35644 25678 35646 25730
rect 35698 25678 35700 25730
rect 35644 25620 35700 25678
rect 35644 24722 35700 25564
rect 35644 24670 35646 24722
rect 35698 24670 35700 24722
rect 35644 24658 35700 24670
rect 35532 23426 35588 23436
rect 35756 23268 35812 26460
rect 35868 26180 35924 26460
rect 35980 26404 36036 26414
rect 35980 26310 36036 26348
rect 35868 26124 36036 26180
rect 35868 25732 35924 25742
rect 35868 25638 35924 25676
rect 35868 25508 35924 25518
rect 35868 24722 35924 25452
rect 35868 24670 35870 24722
rect 35922 24670 35924 24722
rect 35868 24658 35924 24670
rect 35980 24724 36036 26124
rect 35980 24658 36036 24668
rect 35980 24498 36036 24510
rect 35980 24446 35982 24498
rect 36034 24446 36036 24498
rect 35980 24388 36036 24446
rect 35980 24322 36036 24332
rect 35980 23828 36036 23838
rect 35980 23734 36036 23772
rect 35644 23212 35812 23268
rect 35868 23266 35924 23278
rect 35868 23214 35870 23266
rect 35922 23214 35924 23266
rect 35196 22876 35588 22932
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35532 22596 35588 22876
rect 35084 22530 35140 22540
rect 35196 22540 35588 22596
rect 35196 22482 35252 22540
rect 35196 22430 35198 22482
rect 35250 22430 35252 22482
rect 34860 22316 35028 22372
rect 34860 22148 34916 22158
rect 34524 22146 34916 22148
rect 34524 22094 34862 22146
rect 34914 22094 34916 22146
rect 34524 22092 34916 22094
rect 34860 22082 34916 22092
rect 34412 21980 34804 22036
rect 34300 21868 34692 21924
rect 34188 21756 34356 21812
rect 34076 21644 34244 21700
rect 33964 21532 34132 21588
rect 34076 21474 34132 21532
rect 34076 21422 34078 21474
rect 34130 21422 34132 21474
rect 33964 21364 34020 21374
rect 33964 21270 34020 21308
rect 33964 20244 34020 20254
rect 33964 19012 34020 20188
rect 34076 19236 34132 21422
rect 34188 19572 34244 21644
rect 34300 20356 34356 21756
rect 34636 21810 34692 21868
rect 34636 21758 34638 21810
rect 34690 21758 34692 21810
rect 34300 20290 34356 20300
rect 34412 20802 34468 20814
rect 34412 20750 34414 20802
rect 34466 20750 34468 20802
rect 34188 19506 34244 19516
rect 34300 20018 34356 20030
rect 34300 19966 34302 20018
rect 34354 19966 34356 20018
rect 34300 19460 34356 19966
rect 34300 19394 34356 19404
rect 34412 19236 34468 20750
rect 34524 20578 34580 20590
rect 34524 20526 34526 20578
rect 34578 20526 34580 20578
rect 34524 20356 34580 20526
rect 34636 20468 34692 21758
rect 34748 20802 34804 21980
rect 34972 21588 35028 22316
rect 34860 21532 35028 21588
rect 34860 21364 34916 21532
rect 35196 21364 35252 22430
rect 35420 22372 35476 22382
rect 35420 21588 35476 22316
rect 35644 22260 35700 23212
rect 35868 23156 35924 23214
rect 36092 23156 36148 28476
rect 36204 24836 36260 30044
rect 36316 29204 36372 32844
rect 36428 32674 36484 33068
rect 36428 32622 36430 32674
rect 36482 32622 36484 32674
rect 36428 31892 36484 32622
rect 36428 31666 36484 31836
rect 36764 31778 36820 33964
rect 36876 33570 36932 35196
rect 37548 35138 37604 35868
rect 37548 35086 37550 35138
rect 37602 35086 37604 35138
rect 37548 35074 37604 35086
rect 37772 35026 37828 38668
rect 37996 38162 38052 38174
rect 37996 38110 37998 38162
rect 38050 38110 38052 38162
rect 37996 37604 38052 38110
rect 37996 37538 38052 37548
rect 38220 37938 38276 38892
rect 38332 38882 38388 38892
rect 38220 37886 38222 37938
rect 38274 37886 38276 37938
rect 38108 37268 38164 37278
rect 38220 37268 38276 37886
rect 38556 38612 38612 38622
rect 38108 37266 38276 37268
rect 38108 37214 38110 37266
rect 38162 37214 38276 37266
rect 38108 37212 38276 37214
rect 38332 37604 38388 37614
rect 38556 37604 38612 38556
rect 39004 38164 39060 39340
rect 39228 39330 39284 39340
rect 39452 39394 39508 39406
rect 39452 39342 39454 39394
rect 39506 39342 39508 39394
rect 39452 39058 39508 39342
rect 39452 39006 39454 39058
rect 39506 39006 39508 39058
rect 39452 38994 39508 39006
rect 40012 38836 40068 38846
rect 40012 38742 40068 38780
rect 39564 38724 39620 38734
rect 39452 38668 39564 38724
rect 38388 37548 38612 37604
rect 38668 38108 39060 38164
rect 39340 38388 39396 38398
rect 38332 37266 38388 37548
rect 38668 37490 38724 38108
rect 38668 37438 38670 37490
rect 38722 37438 38724 37490
rect 38668 37426 38724 37438
rect 38332 37214 38334 37266
rect 38386 37214 38388 37266
rect 38108 37202 38164 37212
rect 38332 37202 38388 37214
rect 38668 36596 38724 36606
rect 38444 36260 38500 36270
rect 38444 36036 38500 36204
rect 38668 36260 38724 36540
rect 38668 36194 38724 36204
rect 39116 36370 39172 36382
rect 39116 36318 39118 36370
rect 39170 36318 39172 36370
rect 38444 35922 38500 35980
rect 38444 35870 38446 35922
rect 38498 35870 38500 35922
rect 38444 35858 38500 35870
rect 39004 36036 39060 36046
rect 39004 35922 39060 35980
rect 39004 35870 39006 35922
rect 39058 35870 39060 35922
rect 39004 35858 39060 35870
rect 39116 35922 39172 36318
rect 39116 35870 39118 35922
rect 39170 35870 39172 35922
rect 39116 35858 39172 35870
rect 39228 36372 39284 36382
rect 39228 35810 39284 36316
rect 39228 35758 39230 35810
rect 39282 35758 39284 35810
rect 39228 35746 39284 35758
rect 37772 34974 37774 35026
rect 37826 34974 37828 35026
rect 37772 34962 37828 34974
rect 37772 34690 37828 34702
rect 37772 34638 37774 34690
rect 37826 34638 37828 34690
rect 37100 34468 37156 34478
rect 37100 34242 37156 34412
rect 37100 34190 37102 34242
rect 37154 34190 37156 34242
rect 37100 34178 37156 34190
rect 37212 34356 37268 34366
rect 36876 33518 36878 33570
rect 36930 33518 36932 33570
rect 36876 33506 36932 33518
rect 37212 32786 37268 34300
rect 37772 34356 37828 34638
rect 39004 34692 39060 34702
rect 39004 34598 39060 34636
rect 37772 34290 37828 34300
rect 39340 34244 39396 38332
rect 39452 38276 39508 38668
rect 39564 38592 39620 38668
rect 40460 38724 40516 38734
rect 40460 38630 40516 38668
rect 39452 38050 39508 38220
rect 39452 37998 39454 38050
rect 39506 37998 39508 38050
rect 39452 37986 39508 37998
rect 40124 37938 40180 37950
rect 40124 37886 40126 37938
rect 40178 37886 40180 37938
rect 40124 36484 40180 37886
rect 40796 36594 40852 39788
rect 40796 36542 40798 36594
rect 40850 36542 40852 36594
rect 40796 36530 40852 36542
rect 41132 37826 41188 37838
rect 41132 37774 41134 37826
rect 41186 37774 41188 37826
rect 41132 36932 41188 37774
rect 40124 36352 40180 36428
rect 41132 36036 41188 36876
rect 41132 35970 41188 35980
rect 39900 34914 39956 34926
rect 39900 34862 39902 34914
rect 39954 34862 39956 34914
rect 39340 34178 39396 34188
rect 39452 34692 39508 34702
rect 39900 34692 39956 34862
rect 39452 34690 39956 34692
rect 39452 34638 39454 34690
rect 39506 34638 39956 34690
rect 39452 34636 39956 34638
rect 40460 34914 40516 34926
rect 40460 34862 40462 34914
rect 40514 34862 40516 34914
rect 40460 34692 40516 34862
rect 38220 34020 38276 34030
rect 38220 33926 38276 33964
rect 37212 32734 37214 32786
rect 37266 32734 37268 32786
rect 37212 32722 37268 32734
rect 37436 33348 37492 33358
rect 37436 32788 37492 33292
rect 37660 33348 37716 33358
rect 37996 33348 38052 33358
rect 37548 32788 37604 32798
rect 37436 32786 37604 32788
rect 37436 32734 37550 32786
rect 37602 32734 37604 32786
rect 37436 32732 37604 32734
rect 37548 32676 37604 32732
rect 37548 32610 37604 32620
rect 36764 31726 36766 31778
rect 36818 31726 36820 31778
rect 36764 31714 36820 31726
rect 36428 31614 36430 31666
rect 36482 31614 36484 31666
rect 36428 31602 36484 31614
rect 36764 31332 36820 31342
rect 36428 30322 36484 30334
rect 36428 30270 36430 30322
rect 36482 30270 36484 30322
rect 36428 29764 36484 30270
rect 36428 29698 36484 29708
rect 36652 30322 36708 30334
rect 36652 30270 36654 30322
rect 36706 30270 36708 30322
rect 36652 29876 36708 30270
rect 36764 29986 36820 31276
rect 37436 31108 37492 31118
rect 37436 30996 37492 31052
rect 37660 30996 37716 33292
rect 37884 33346 38052 33348
rect 37884 33294 37998 33346
rect 38050 33294 38052 33346
rect 37884 33292 38052 33294
rect 37884 31332 37940 33292
rect 37996 33282 38052 33292
rect 39452 33348 39508 34636
rect 40460 34626 40516 34636
rect 39452 33282 39508 33292
rect 41020 33348 41076 33358
rect 40348 33122 40404 33134
rect 40348 33070 40350 33122
rect 40402 33070 40404 33122
rect 40348 32900 40404 33070
rect 40236 32844 40404 32900
rect 37996 32676 38052 32686
rect 37996 32582 38052 32620
rect 38668 32452 38724 32462
rect 39116 32452 39172 32462
rect 38668 32450 39172 32452
rect 38668 32398 38670 32450
rect 38722 32398 39118 32450
rect 39170 32398 39172 32450
rect 38668 32396 39172 32398
rect 38444 31668 38500 31678
rect 38444 31574 38500 31612
rect 38668 31668 38724 32396
rect 39116 32386 39172 32396
rect 40236 31948 40292 32844
rect 40348 32674 40404 32686
rect 40348 32622 40350 32674
rect 40402 32622 40404 32674
rect 40348 32340 40404 32622
rect 40348 32284 40516 32340
rect 40460 31948 40516 32284
rect 39452 31890 39508 31902
rect 40236 31892 40404 31948
rect 40460 31892 40628 31948
rect 39452 31838 39454 31890
rect 39506 31838 39508 31890
rect 39452 31780 39508 31838
rect 40124 31780 40180 31790
rect 39452 31778 40292 31780
rect 39452 31726 40126 31778
rect 40178 31726 40292 31778
rect 39452 31724 40292 31726
rect 40124 31714 40180 31724
rect 38668 31602 38724 31612
rect 37884 31266 37940 31276
rect 40124 31556 40180 31566
rect 37436 30994 37716 30996
rect 37436 30942 37438 30994
rect 37490 30942 37716 30994
rect 37436 30940 37716 30942
rect 37436 30930 37492 30940
rect 37660 30436 37716 30940
rect 37660 30370 37716 30380
rect 37772 30994 37828 31006
rect 37772 30942 37774 30994
rect 37826 30942 37828 30994
rect 36764 29934 36766 29986
rect 36818 29934 36820 29986
rect 36764 29922 36820 29934
rect 37436 29986 37492 29998
rect 37436 29934 37438 29986
rect 37490 29934 37492 29986
rect 36540 29540 36596 29550
rect 36540 29446 36596 29484
rect 36428 29428 36484 29438
rect 36428 29334 36484 29372
rect 36652 29428 36708 29820
rect 37436 29764 37492 29934
rect 37436 29698 37492 29708
rect 37660 29652 37716 29662
rect 37772 29652 37828 30942
rect 38108 30436 38164 30446
rect 38108 30342 38164 30380
rect 37660 29650 37828 29652
rect 37660 29598 37662 29650
rect 37714 29598 37828 29650
rect 37660 29596 37828 29598
rect 37660 29586 37716 29596
rect 37884 29540 37940 29550
rect 36652 29362 36708 29372
rect 36764 29428 36820 29438
rect 37100 29428 37156 29438
rect 36764 29426 37156 29428
rect 36764 29374 36766 29426
rect 36818 29374 37102 29426
rect 37154 29374 37156 29426
rect 36764 29372 37156 29374
rect 36764 29362 36820 29372
rect 37100 29362 37156 29372
rect 37324 29428 37380 29438
rect 36316 29148 36484 29204
rect 36316 26852 36372 26862
rect 36316 26758 36372 26796
rect 36428 26068 36484 29148
rect 36540 28866 36596 28878
rect 36540 28814 36542 28866
rect 36594 28814 36596 28866
rect 36540 28754 36596 28814
rect 36540 28702 36542 28754
rect 36594 28702 36596 28754
rect 36540 28690 36596 28702
rect 37324 28084 37380 29372
rect 37548 29426 37604 29438
rect 37548 29374 37550 29426
rect 37602 29374 37604 29426
rect 37548 28644 37604 29374
rect 37772 29428 37828 29438
rect 37772 29334 37828 29372
rect 37548 28578 37604 28588
rect 37772 28644 37828 28654
rect 37884 28644 37940 29484
rect 38332 29540 38388 29550
rect 38332 29446 38388 29484
rect 38668 29540 38724 29550
rect 38668 29446 38724 29484
rect 39116 29540 39172 29550
rect 39116 29446 39172 29484
rect 37772 28642 37940 28644
rect 37772 28590 37774 28642
rect 37826 28590 37940 28642
rect 37772 28588 37940 28590
rect 37772 28578 37828 28588
rect 37436 28420 37492 28430
rect 37436 28326 37492 28364
rect 37660 28418 37716 28430
rect 37660 28366 37662 28418
rect 37714 28366 37716 28418
rect 37548 28084 37604 28094
rect 37324 28082 37604 28084
rect 37324 28030 37550 28082
rect 37602 28030 37604 28082
rect 37324 28028 37604 28030
rect 37548 28018 37604 28028
rect 36540 27748 36596 27758
rect 36988 27748 37044 27758
rect 36596 27746 37044 27748
rect 36596 27694 36990 27746
rect 37042 27694 37044 27746
rect 36596 27692 37044 27694
rect 36540 27616 36596 27692
rect 36764 27524 36820 27534
rect 36764 26404 36820 27468
rect 36876 26962 36932 26974
rect 36876 26910 36878 26962
rect 36930 26910 36932 26962
rect 36876 26516 36932 26910
rect 36988 26964 37044 27692
rect 37548 27636 37604 27646
rect 36988 26898 37044 26908
rect 37100 27412 37156 27422
rect 36876 26450 36932 26460
rect 37100 26514 37156 27356
rect 37100 26462 37102 26514
rect 37154 26462 37156 26514
rect 37100 26450 37156 26462
rect 36764 26338 36820 26348
rect 36428 26002 36484 26012
rect 36540 26290 36596 26302
rect 36540 26238 36542 26290
rect 36594 26238 36596 26290
rect 36540 25844 36596 26238
rect 36540 25732 36596 25788
rect 36316 25676 36596 25732
rect 36876 26290 36932 26302
rect 36876 26238 36878 26290
rect 36930 26238 36932 26290
rect 36316 25284 36372 25676
rect 36876 25620 36932 26238
rect 37548 26180 37604 27580
rect 37660 27074 37716 28366
rect 37772 28196 37828 28206
rect 37772 27636 37828 28140
rect 37772 27570 37828 27580
rect 37884 27412 37940 28588
rect 38220 29204 38276 29214
rect 38220 28644 38276 29148
rect 38220 28550 38276 28588
rect 38780 28756 38836 28766
rect 38444 27972 38500 27982
rect 38500 27916 38612 27972
rect 37884 27346 37940 27356
rect 38108 27858 38164 27870
rect 38108 27806 38110 27858
rect 38162 27806 38164 27858
rect 38444 27840 38500 27916
rect 37660 27022 37662 27074
rect 37714 27022 37716 27074
rect 37660 26964 37716 27022
rect 37996 27076 38052 27086
rect 37996 26982 38052 27020
rect 37660 26514 37716 26908
rect 37660 26462 37662 26514
rect 37714 26462 37716 26514
rect 37660 26450 37716 26462
rect 37772 26962 37828 26974
rect 37772 26910 37774 26962
rect 37826 26910 37828 26962
rect 37548 26124 37716 26180
rect 37212 26066 37268 26078
rect 37212 26014 37214 26066
rect 37266 26014 37268 26066
rect 37100 25956 37156 25966
rect 37212 25956 37268 26014
rect 37212 25900 37380 25956
rect 37100 25844 37156 25900
rect 37100 25788 37268 25844
rect 36428 25564 36932 25620
rect 36428 25394 36484 25564
rect 36876 25508 36932 25564
rect 36876 25442 36932 25452
rect 36988 25732 37044 25742
rect 36428 25342 36430 25394
rect 36482 25342 36484 25394
rect 36428 25330 36484 25342
rect 36764 25394 36820 25406
rect 36764 25342 36766 25394
rect 36818 25342 36820 25394
rect 36316 25218 36372 25228
rect 36764 25284 36820 25342
rect 36988 25284 37044 25676
rect 36764 25218 36820 25228
rect 36876 25228 37044 25284
rect 37100 25620 37156 25630
rect 36764 24836 36820 24912
rect 36204 24770 36260 24780
rect 36428 24780 36764 24836
rect 36316 24500 36372 24510
rect 36428 24500 36484 24780
rect 36764 24770 36820 24780
rect 36652 24610 36708 24622
rect 36652 24558 36654 24610
rect 36706 24558 36708 24610
rect 36372 24444 36484 24500
rect 36540 24498 36596 24510
rect 36540 24446 36542 24498
rect 36594 24446 36596 24498
rect 36316 24434 36372 24444
rect 36540 24388 36596 24446
rect 36540 24322 36596 24332
rect 36540 23940 36596 23950
rect 36316 23828 36372 23838
rect 36316 23734 36372 23772
rect 36540 23716 36596 23884
rect 36540 23378 36596 23660
rect 36652 23604 36708 24558
rect 36652 23538 36708 23548
rect 36764 24612 36820 24622
rect 36764 23714 36820 24556
rect 36764 23662 36766 23714
rect 36818 23662 36820 23714
rect 36540 23326 36542 23378
rect 36594 23326 36596 23378
rect 36540 23314 36596 23326
rect 36764 23268 36820 23662
rect 36764 23202 36820 23212
rect 35868 23090 35924 23100
rect 35980 23100 36148 23156
rect 36540 23156 36596 23166
rect 35756 23044 35812 23054
rect 35756 22950 35812 22988
rect 35756 22596 35812 22606
rect 35756 22482 35812 22540
rect 35756 22430 35758 22482
rect 35810 22430 35812 22482
rect 35756 22418 35812 22430
rect 35980 22260 36036 23100
rect 36092 22932 36148 22942
rect 36316 22932 36372 22942
rect 36092 22930 36372 22932
rect 36092 22878 36094 22930
rect 36146 22878 36318 22930
rect 36370 22878 36372 22930
rect 36092 22876 36372 22878
rect 36092 22866 36148 22876
rect 36316 22866 36372 22876
rect 36092 22708 36148 22718
rect 36092 22594 36148 22652
rect 36092 22542 36094 22594
rect 36146 22542 36148 22594
rect 36092 22482 36148 22542
rect 36092 22430 36094 22482
rect 36146 22430 36148 22482
rect 36092 22418 36148 22430
rect 36428 22708 36484 22718
rect 36428 22260 36484 22652
rect 36540 22482 36596 23100
rect 36540 22430 36542 22482
rect 36594 22430 36596 22482
rect 36540 22418 36596 22430
rect 36652 22930 36708 22942
rect 36652 22878 36654 22930
rect 36706 22878 36708 22930
rect 35644 22204 35924 22260
rect 35980 22204 36148 22260
rect 36428 22204 36596 22260
rect 35420 21586 35700 21588
rect 35420 21534 35422 21586
rect 35474 21534 35700 21586
rect 35420 21532 35700 21534
rect 35420 21522 35476 21532
rect 34860 21308 35028 21364
rect 34748 20750 34750 20802
rect 34802 20750 34804 20802
rect 34748 20738 34804 20750
rect 34860 21026 34916 21038
rect 34860 20974 34862 21026
rect 34914 20974 34916 21026
rect 34636 20402 34692 20412
rect 34524 20290 34580 20300
rect 34860 20130 34916 20974
rect 34972 20802 35028 21308
rect 34972 20750 34974 20802
rect 35026 20750 35028 20802
rect 34972 20244 35028 20750
rect 35084 21308 35252 21364
rect 35532 21362 35588 21374
rect 35532 21310 35534 21362
rect 35586 21310 35588 21362
rect 35084 20244 35140 21308
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35532 20916 35588 21310
rect 35644 21364 35700 21532
rect 35756 21364 35812 21374
rect 35644 21362 35812 21364
rect 35644 21310 35758 21362
rect 35810 21310 35812 21362
rect 35644 21308 35812 21310
rect 35756 21298 35812 21308
rect 35532 20850 35588 20860
rect 35532 20578 35588 20590
rect 35532 20526 35534 20578
rect 35586 20526 35588 20578
rect 35420 20244 35476 20254
rect 35084 20188 35252 20244
rect 34972 20178 35028 20188
rect 34860 20078 34862 20130
rect 34914 20078 34916 20130
rect 34860 20066 34916 20078
rect 35084 20018 35140 20030
rect 35084 19966 35086 20018
rect 35138 19966 35140 20018
rect 34972 19908 35028 19918
rect 34636 19906 35028 19908
rect 34636 19854 34974 19906
rect 35026 19854 35028 19906
rect 34636 19852 35028 19854
rect 34524 19236 34580 19246
rect 34412 19234 34580 19236
rect 34412 19182 34526 19234
rect 34578 19182 34580 19234
rect 34412 19180 34580 19182
rect 34076 19170 34132 19180
rect 34188 19012 34244 19022
rect 33964 19010 34244 19012
rect 33964 18958 34190 19010
rect 34242 18958 34244 19010
rect 33964 18956 34244 18958
rect 34188 18946 34244 18956
rect 33964 18340 34020 18350
rect 33964 18246 34020 18284
rect 33852 17614 33854 17666
rect 33906 17614 33908 17666
rect 33852 17602 33908 17614
rect 34412 17668 34468 17678
rect 34412 17574 34468 17612
rect 33740 17556 33796 17566
rect 33628 17444 33684 17454
rect 33628 17350 33684 17388
rect 33628 16884 33684 16922
rect 33628 16818 33684 16828
rect 33740 16772 33796 17500
rect 33852 17444 33908 17454
rect 33852 16996 33908 17388
rect 34524 17444 34580 19180
rect 33964 16996 34020 17006
rect 33852 16994 34020 16996
rect 33852 16942 33966 16994
rect 34018 16942 34020 16994
rect 33852 16940 34020 16942
rect 33964 16930 34020 16940
rect 34524 16994 34580 17388
rect 34524 16942 34526 16994
rect 34578 16942 34580 16994
rect 34524 16930 34580 16942
rect 33740 16716 34244 16772
rect 33516 16270 33518 16322
rect 33570 16270 33572 16322
rect 33516 16258 33572 16270
rect 33628 16658 33684 16670
rect 33628 16606 33630 16658
rect 33682 16606 33684 16658
rect 33404 16212 33460 16222
rect 33180 16210 33460 16212
rect 33180 16158 33406 16210
rect 33458 16158 33460 16210
rect 33180 16156 33460 16158
rect 33404 16146 33460 16156
rect 33628 15314 33684 16606
rect 34188 16210 34244 16716
rect 34188 16158 34190 16210
rect 34242 16158 34244 16210
rect 34188 16146 34244 16158
rect 34300 16548 34356 16558
rect 33740 15988 33796 15998
rect 33740 15894 33796 15932
rect 33628 15262 33630 15314
rect 33682 15262 33684 15314
rect 33292 15204 33348 15214
rect 33180 14868 33236 14878
rect 33180 13188 33236 14812
rect 33292 14308 33348 15148
rect 33292 14214 33348 14252
rect 33180 13132 33348 13188
rect 33180 12962 33236 12974
rect 33180 12910 33182 12962
rect 33234 12910 33236 12962
rect 33180 12852 33236 12910
rect 33180 12786 33236 12796
rect 33180 11172 33236 11182
rect 33180 10724 33236 11116
rect 33180 10658 33236 10668
rect 33180 10052 33236 10062
rect 33180 9958 33236 9996
rect 32956 9772 33124 9828
rect 32844 9268 32900 9278
rect 32844 9174 32900 9212
rect 32956 7812 33012 9772
rect 33068 9604 33124 9614
rect 33068 9510 33124 9548
rect 33292 9044 33348 13132
rect 33628 12964 33684 15262
rect 33740 15652 33796 15662
rect 33740 15316 33796 15596
rect 33964 15316 34020 15326
rect 33740 15314 34132 15316
rect 33740 15262 33966 15314
rect 34018 15262 34132 15314
rect 33740 15260 34132 15262
rect 33740 14642 33796 15260
rect 33964 15250 34020 15260
rect 33740 14590 33742 14642
rect 33794 14590 33796 14642
rect 33740 14578 33796 14590
rect 33964 12964 34020 12974
rect 33628 12908 33796 12964
rect 33628 12738 33684 12750
rect 33628 12686 33630 12738
rect 33682 12686 33684 12738
rect 33516 12068 33572 12078
rect 33516 11974 33572 12012
rect 33628 11844 33684 12686
rect 33628 11778 33684 11788
rect 33628 11396 33684 11406
rect 33628 11302 33684 11340
rect 33740 10724 33796 12908
rect 33964 12870 34020 12908
rect 33852 12852 33908 12862
rect 33852 12758 33908 12796
rect 33964 12066 34020 12078
rect 33964 12014 33966 12066
rect 34018 12014 34020 12066
rect 33964 11956 34020 12014
rect 33964 11890 34020 11900
rect 34076 11172 34132 15260
rect 34188 11956 34244 11966
rect 34188 11506 34244 11900
rect 34188 11454 34190 11506
rect 34242 11454 34244 11506
rect 34188 11442 34244 11454
rect 33628 10668 33796 10724
rect 33852 11116 34132 11172
rect 33404 10052 33460 10062
rect 33628 10052 33684 10668
rect 33404 10050 33684 10052
rect 33404 9998 33406 10050
rect 33458 9998 33684 10050
rect 33404 9996 33684 9998
rect 33404 9986 33460 9996
rect 33628 9044 33684 9996
rect 33740 10500 33796 10510
rect 33740 10052 33796 10444
rect 33740 9986 33796 9996
rect 33852 9826 33908 11116
rect 34300 10948 34356 16492
rect 34188 10892 34356 10948
rect 34524 15988 34580 15998
rect 34188 10612 34244 10892
rect 34188 10546 34244 10556
rect 34300 10610 34356 10622
rect 34300 10558 34302 10610
rect 34354 10558 34356 10610
rect 33964 10052 34020 10062
rect 33964 9958 34020 9996
rect 33852 9774 33854 9826
rect 33906 9774 33908 9826
rect 33852 9268 33908 9774
rect 33292 8988 33572 9044
rect 33292 8484 33348 8494
rect 33292 8370 33348 8428
rect 33292 8318 33294 8370
rect 33346 8318 33348 8370
rect 33292 8306 33348 8318
rect 33068 8148 33124 8158
rect 33068 8054 33124 8092
rect 33180 8036 33236 8046
rect 33180 7942 33236 7980
rect 32956 7756 33236 7812
rect 32844 6692 32900 6702
rect 32844 6598 32900 6636
rect 33068 6690 33124 6702
rect 33068 6638 33070 6690
rect 33122 6638 33124 6690
rect 32956 6466 33012 6478
rect 32956 6414 32958 6466
rect 33010 6414 33012 6466
rect 32956 5122 33012 6414
rect 33068 6468 33124 6638
rect 33180 6468 33236 7756
rect 33292 6802 33348 6814
rect 33292 6750 33294 6802
rect 33346 6750 33348 6802
rect 33292 6692 33348 6750
rect 33292 6626 33348 6636
rect 33180 6412 33348 6468
rect 33068 6402 33124 6412
rect 32956 5070 32958 5122
rect 33010 5070 33012 5122
rect 32956 5058 33012 5070
rect 32956 4898 33012 4910
rect 32956 4846 32958 4898
rect 33010 4846 33012 4898
rect 32956 4564 33012 4846
rect 32956 4498 33012 4508
rect 33180 4676 33236 4686
rect 33180 3666 33236 4620
rect 33180 3614 33182 3666
rect 33234 3614 33236 3666
rect 33180 3602 33236 3614
rect 32732 2818 32788 2828
rect 28476 1586 28532 1596
rect 33292 1540 33348 6412
rect 33516 5012 33572 8988
rect 33628 8978 33684 8988
rect 33740 9044 33796 9054
rect 33852 9044 33908 9212
rect 34076 9716 34132 9726
rect 33740 9042 33908 9044
rect 33740 8990 33742 9042
rect 33794 8990 33908 9042
rect 33740 8988 33908 8990
rect 33964 9044 34020 9054
rect 34076 9044 34132 9660
rect 34300 9156 34356 10558
rect 34412 10498 34468 10510
rect 34412 10446 34414 10498
rect 34466 10446 34468 10498
rect 34412 10164 34468 10446
rect 34412 10098 34468 10108
rect 34300 9090 34356 9100
rect 34412 9940 34468 9950
rect 33964 9042 34132 9044
rect 33964 8990 33966 9042
rect 34018 8990 34132 9042
rect 33964 8988 34132 8990
rect 34188 9044 34244 9054
rect 33740 8978 33796 8988
rect 33964 8978 34020 8988
rect 34188 8950 34244 8988
rect 34412 9042 34468 9884
rect 34412 8990 34414 9042
rect 34466 8990 34468 9042
rect 34412 8932 34468 8990
rect 34412 8866 34468 8876
rect 33628 8818 33684 8830
rect 33628 8766 33630 8818
rect 33682 8766 33684 8818
rect 33628 8484 33684 8766
rect 33628 8418 33684 8428
rect 34188 8258 34244 8270
rect 34188 8206 34190 8258
rect 34242 8206 34244 8258
rect 34188 8148 34244 8206
rect 34188 8082 34244 8092
rect 34524 7476 34580 15932
rect 34636 10836 34692 19852
rect 34972 19842 35028 19852
rect 34972 19460 35028 19470
rect 35084 19460 35140 19966
rect 35196 19908 35252 20188
rect 35420 20130 35476 20188
rect 35420 20078 35422 20130
rect 35474 20078 35476 20130
rect 35420 20066 35476 20078
rect 35532 20132 35588 20526
rect 35532 20066 35588 20076
rect 35868 20356 35924 22204
rect 35980 21812 36036 21822
rect 35980 21718 36036 21756
rect 36092 21028 36148 22204
rect 36428 21474 36484 21486
rect 36428 21422 36430 21474
rect 36482 21422 36484 21474
rect 36428 21364 36484 21422
rect 36428 21298 36484 21308
rect 36092 20972 36484 21028
rect 35868 20130 35924 20300
rect 35868 20078 35870 20130
rect 35922 20078 35924 20130
rect 35868 20066 35924 20078
rect 35980 20690 36036 20702
rect 35980 20638 35982 20690
rect 36034 20638 36036 20690
rect 35196 19842 35252 19852
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35084 19404 35364 19460
rect 34860 19236 34916 19246
rect 34860 19142 34916 19180
rect 34748 19124 34804 19134
rect 34748 19030 34804 19068
rect 34860 18564 34916 18574
rect 34748 18338 34804 18350
rect 34748 18286 34750 18338
rect 34802 18286 34804 18338
rect 34748 17892 34804 18286
rect 34748 17826 34804 17836
rect 34748 17108 34804 17118
rect 34748 17014 34804 17052
rect 34860 16660 34916 18508
rect 34972 18450 35028 19404
rect 35308 19234 35364 19404
rect 35308 19182 35310 19234
rect 35362 19182 35364 19234
rect 35308 19170 35364 19182
rect 35644 19122 35700 19134
rect 35644 19070 35646 19122
rect 35698 19070 35700 19122
rect 35532 19012 35588 19022
rect 35532 18918 35588 18956
rect 35308 18564 35364 18574
rect 35644 18564 35700 19070
rect 35980 18788 36036 20638
rect 36092 20690 36148 20702
rect 36092 20638 36094 20690
rect 36146 20638 36148 20690
rect 36092 19908 36148 20638
rect 36204 20692 36260 20702
rect 36204 20598 36260 20636
rect 36092 19842 36148 19852
rect 36204 20244 36260 20254
rect 36204 19346 36260 20188
rect 36204 19294 36206 19346
rect 36258 19294 36260 19346
rect 36204 19282 36260 19294
rect 36316 19906 36372 19918
rect 36316 19854 36318 19906
rect 36370 19854 36372 19906
rect 36316 19460 36372 19854
rect 35364 18508 35700 18564
rect 35756 18732 36036 18788
rect 34972 18398 34974 18450
rect 35026 18398 35028 18450
rect 34972 17108 35028 18398
rect 35084 18452 35140 18462
rect 35308 18432 35364 18508
rect 35756 18452 35812 18732
rect 35084 17666 35140 18396
rect 35756 18320 35812 18396
rect 35980 18562 36036 18574
rect 35980 18510 35982 18562
rect 36034 18510 36036 18562
rect 35980 18340 36036 18510
rect 36092 18564 36148 18574
rect 36092 18470 36148 18508
rect 36316 18452 36372 19404
rect 36316 18386 36372 18396
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35980 17892 36036 18284
rect 35980 17826 36036 17836
rect 35084 17614 35086 17666
rect 35138 17614 35140 17666
rect 35084 17602 35140 17614
rect 35308 17668 35364 17678
rect 36204 17668 36260 17678
rect 35308 17666 36260 17668
rect 35308 17614 35310 17666
rect 35362 17614 36206 17666
rect 36258 17614 36260 17666
rect 35308 17612 36260 17614
rect 35308 17602 35364 17612
rect 36204 17602 36260 17612
rect 35196 17554 35252 17566
rect 35196 17502 35198 17554
rect 35250 17502 35252 17554
rect 34972 17042 35028 17052
rect 35084 17332 35140 17342
rect 34972 16884 35028 16894
rect 34972 16790 35028 16828
rect 34748 16322 34804 16334
rect 34748 16270 34750 16322
rect 34802 16270 34804 16322
rect 34748 16210 34804 16270
rect 34748 16158 34750 16210
rect 34802 16158 34804 16210
rect 34748 16146 34804 16158
rect 34860 15426 34916 16604
rect 34860 15374 34862 15426
rect 34914 15374 34916 15426
rect 34860 15362 34916 15374
rect 35084 15314 35140 17276
rect 35196 17106 35252 17502
rect 35756 17442 35812 17454
rect 35756 17390 35758 17442
rect 35810 17390 35812 17442
rect 35196 17054 35198 17106
rect 35250 17054 35252 17106
rect 35196 17042 35252 17054
rect 35308 17108 35364 17118
rect 35196 16884 35252 16894
rect 35308 16884 35364 17052
rect 35196 16882 35364 16884
rect 35196 16830 35198 16882
rect 35250 16830 35364 16882
rect 35196 16828 35364 16830
rect 35532 16884 35588 16894
rect 35196 16818 35252 16828
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35084 15262 35086 15314
rect 35138 15262 35140 15314
rect 35084 15250 35140 15262
rect 35196 15876 35252 15886
rect 34972 15202 35028 15214
rect 34972 15150 34974 15202
rect 35026 15150 35028 15202
rect 34860 13860 34916 13870
rect 34860 13074 34916 13804
rect 34860 13022 34862 13074
rect 34914 13022 34916 13074
rect 34860 13010 34916 13022
rect 34748 12852 34804 12862
rect 34748 12850 34916 12852
rect 34748 12798 34750 12850
rect 34802 12798 34916 12850
rect 34748 12796 34916 12798
rect 34748 12786 34804 12796
rect 34748 12404 34804 12414
rect 34748 12310 34804 12348
rect 34860 11284 34916 12796
rect 34860 11218 34916 11228
rect 34636 10780 34804 10836
rect 34636 10610 34692 10622
rect 34636 10558 34638 10610
rect 34690 10558 34692 10610
rect 34636 9268 34692 10558
rect 34748 10610 34804 10780
rect 34748 10558 34750 10610
rect 34802 10558 34804 10610
rect 34748 9938 34804 10558
rect 34748 9886 34750 9938
rect 34802 9886 34804 9938
rect 34748 9828 34804 9886
rect 34860 9940 34916 9950
rect 34860 9846 34916 9884
rect 34972 9828 35028 15150
rect 35196 15092 35252 15820
rect 35196 15026 35252 15036
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35308 14642 35364 14654
rect 35308 14590 35310 14642
rect 35362 14590 35364 14642
rect 35308 14532 35364 14590
rect 35308 14466 35364 14476
rect 35420 14420 35476 14430
rect 35532 14420 35588 16828
rect 35644 16772 35700 16782
rect 35644 16210 35700 16716
rect 35644 16158 35646 16210
rect 35698 16158 35700 16210
rect 35644 16146 35700 16158
rect 35756 15652 35812 17390
rect 36092 17444 36148 17454
rect 35980 17332 36036 17342
rect 35980 16884 36036 17276
rect 35980 16818 36036 16828
rect 36092 16770 36148 17388
rect 36316 17442 36372 17454
rect 36316 17390 36318 17442
rect 36370 17390 36372 17442
rect 36316 17332 36372 17390
rect 36316 17266 36372 17276
rect 36316 16884 36372 16894
rect 36316 16790 36372 16828
rect 36092 16718 36094 16770
rect 36146 16718 36148 16770
rect 36092 16706 36148 16718
rect 35868 16660 35924 16670
rect 36428 16660 36484 20972
rect 36540 19346 36596 22204
rect 36652 21028 36708 22878
rect 36652 20962 36708 20972
rect 36764 21362 36820 21374
rect 36764 21310 36766 21362
rect 36818 21310 36820 21362
rect 36764 20914 36820 21310
rect 36764 20862 36766 20914
rect 36818 20862 36820 20914
rect 36764 20850 36820 20862
rect 36540 19294 36542 19346
rect 36594 19294 36596 19346
rect 36540 19124 36596 19294
rect 36540 19058 36596 19068
rect 36652 20468 36708 20478
rect 36540 18452 36596 18462
rect 36540 18358 36596 18396
rect 36540 17668 36596 17678
rect 36652 17668 36708 20412
rect 36876 20130 36932 25228
rect 37100 23378 37156 25564
rect 37100 23326 37102 23378
rect 37154 23326 37156 23378
rect 37100 23314 37156 23326
rect 37100 21700 37156 21710
rect 37100 21606 37156 21644
rect 36988 21586 37044 21598
rect 36988 21534 36990 21586
rect 37042 21534 37044 21586
rect 36988 21476 37044 21534
rect 37212 21476 37268 25788
rect 37324 25732 37380 25900
rect 37548 25732 37604 25742
rect 37324 25730 37604 25732
rect 37324 25678 37550 25730
rect 37602 25678 37604 25730
rect 37324 25676 37604 25678
rect 37660 25732 37716 26124
rect 37772 26068 37828 26910
rect 38108 26964 38164 27806
rect 38444 27300 38500 27310
rect 38220 27188 38276 27198
rect 38220 27074 38276 27132
rect 38220 27022 38222 27074
rect 38274 27022 38276 27074
rect 38220 27010 38276 27022
rect 38444 27076 38500 27244
rect 38108 26898 38164 26908
rect 38444 26514 38500 27020
rect 38444 26462 38446 26514
rect 38498 26462 38500 26514
rect 38444 26450 38500 26462
rect 37772 26002 37828 26012
rect 37996 26404 38052 26414
rect 37660 25676 37828 25732
rect 37548 25666 37604 25676
rect 37660 25508 37716 25518
rect 37660 25414 37716 25452
rect 37772 25284 37828 25676
rect 37884 25396 37940 25406
rect 37884 25302 37940 25340
rect 37436 25228 37828 25284
rect 37324 24836 37380 24846
rect 37324 24742 37380 24780
rect 37436 24052 37492 25228
rect 37772 25060 37828 25070
rect 37772 24946 37828 25004
rect 37772 24894 37774 24946
rect 37826 24894 37828 24946
rect 37324 23996 37492 24052
rect 37548 24498 37604 24510
rect 37548 24446 37550 24498
rect 37602 24446 37604 24498
rect 37324 22372 37380 23996
rect 37436 23828 37492 23838
rect 37436 23604 37492 23772
rect 37436 23378 37492 23548
rect 37436 23326 37438 23378
rect 37490 23326 37492 23378
rect 37436 23314 37492 23326
rect 37548 23826 37604 24446
rect 37548 23774 37550 23826
rect 37602 23774 37604 23826
rect 37548 22708 37604 23774
rect 37548 22642 37604 22652
rect 37772 22708 37828 24894
rect 37996 24498 38052 26348
rect 38220 26292 38276 26302
rect 38108 25732 38164 25742
rect 38108 25638 38164 25676
rect 38220 24946 38276 26236
rect 38444 26068 38500 26078
rect 38332 25844 38388 25854
rect 38332 25730 38388 25788
rect 38332 25678 38334 25730
rect 38386 25678 38388 25730
rect 38332 25396 38388 25678
rect 38332 25330 38388 25340
rect 38220 24894 38222 24946
rect 38274 24894 38276 24946
rect 38220 24882 38276 24894
rect 38332 25172 38388 25182
rect 38444 25172 38500 26012
rect 38388 25116 38500 25172
rect 37996 24446 37998 24498
rect 38050 24446 38052 24498
rect 37996 24434 38052 24446
rect 37884 23828 37940 23838
rect 37884 23826 38052 23828
rect 37884 23774 37886 23826
rect 37938 23774 38052 23826
rect 37884 23772 38052 23774
rect 37884 23762 37940 23772
rect 37884 23042 37940 23054
rect 37884 22990 37886 23042
rect 37938 22990 37940 23042
rect 37884 22930 37940 22990
rect 37996 23044 38052 23772
rect 38332 23716 38388 25116
rect 38444 23940 38500 23950
rect 38556 23940 38612 27916
rect 38668 26964 38724 26974
rect 38668 26870 38724 26908
rect 38668 24836 38724 24846
rect 38668 24742 38724 24780
rect 38780 24164 38836 28700
rect 39676 27972 39732 27982
rect 39452 27970 39732 27972
rect 39452 27918 39678 27970
rect 39730 27918 39732 27970
rect 39452 27916 39732 27918
rect 39004 27748 39060 27758
rect 39004 27746 39172 27748
rect 39004 27694 39006 27746
rect 39058 27694 39172 27746
rect 39004 27692 39172 27694
rect 39004 27682 39060 27692
rect 38892 27300 38948 27310
rect 38892 27074 38948 27244
rect 38892 27022 38894 27074
rect 38946 27022 38948 27074
rect 38892 27010 38948 27022
rect 38892 26852 38948 26862
rect 38892 26514 38948 26796
rect 38892 26462 38894 26514
rect 38946 26462 38948 26514
rect 38892 26450 38948 26462
rect 39004 26850 39060 26862
rect 39004 26798 39006 26850
rect 39058 26798 39060 26850
rect 38892 25956 38948 25966
rect 38892 25506 38948 25900
rect 39004 25844 39060 26798
rect 39116 26068 39172 27692
rect 39228 26962 39284 26974
rect 39228 26910 39230 26962
rect 39282 26910 39284 26962
rect 39228 26852 39284 26910
rect 39228 26786 39284 26796
rect 39340 26292 39396 26302
rect 39340 26198 39396 26236
rect 39116 26002 39172 26012
rect 39004 25778 39060 25788
rect 39228 25844 39284 25854
rect 38892 25454 38894 25506
rect 38946 25454 38948 25506
rect 38892 25442 38948 25454
rect 39116 25508 39172 25518
rect 39116 25414 39172 25452
rect 38892 24164 38948 24174
rect 38780 24162 38948 24164
rect 38780 24110 38894 24162
rect 38946 24110 38948 24162
rect 38780 24108 38948 24110
rect 38444 23938 38612 23940
rect 38444 23886 38446 23938
rect 38498 23886 38612 23938
rect 38444 23884 38612 23886
rect 38444 23874 38500 23884
rect 38332 23660 38500 23716
rect 38332 23044 38388 23054
rect 37996 23042 38388 23044
rect 37996 22990 38334 23042
rect 38386 22990 38388 23042
rect 37996 22988 38388 22990
rect 37884 22878 37886 22930
rect 37938 22878 37940 22930
rect 37884 22866 37940 22878
rect 37772 22642 37828 22652
rect 37996 22484 38052 22494
rect 37996 22390 38052 22428
rect 37660 22372 37716 22382
rect 37324 22316 37492 22372
rect 37324 22146 37380 22158
rect 37324 22094 37326 22146
rect 37378 22094 37380 22146
rect 37324 21810 37380 22094
rect 37324 21758 37326 21810
rect 37378 21758 37380 21810
rect 37324 21746 37380 21758
rect 36988 21420 37268 21476
rect 36876 20078 36878 20130
rect 36930 20078 36932 20130
rect 36876 20066 36932 20078
rect 36988 20692 37044 20702
rect 36988 20130 37044 20636
rect 36988 20078 36990 20130
rect 37042 20078 37044 20130
rect 36988 20066 37044 20078
rect 37212 20132 37268 21420
rect 37324 20244 37380 20254
rect 37324 20150 37380 20188
rect 37212 20066 37268 20076
rect 37100 20018 37156 20030
rect 37100 19966 37102 20018
rect 37154 19966 37156 20018
rect 37100 19796 37156 19966
rect 37100 19730 37156 19740
rect 37436 19236 37492 22316
rect 37548 22370 37716 22372
rect 37548 22318 37662 22370
rect 37714 22318 37716 22370
rect 37548 22316 37716 22318
rect 37548 22146 37604 22316
rect 37660 22260 37716 22316
rect 37660 22204 37940 22260
rect 37548 22094 37550 22146
rect 37602 22094 37604 22146
rect 37548 22082 37604 22094
rect 37884 21588 37940 22204
rect 37996 22148 38052 22158
rect 37996 22054 38052 22092
rect 37996 21588 38052 21598
rect 37884 21586 38052 21588
rect 37884 21534 37998 21586
rect 38050 21534 38052 21586
rect 37884 21532 38052 21534
rect 37996 21522 38052 21532
rect 38108 21588 38164 22988
rect 38332 22978 38388 22988
rect 38444 22930 38500 23660
rect 38556 23268 38612 23884
rect 38668 23938 38724 23950
rect 38668 23886 38670 23938
rect 38722 23886 38724 23938
rect 38668 23492 38724 23886
rect 38668 23426 38724 23436
rect 38780 23378 38836 24108
rect 38892 24098 38948 24108
rect 39116 23940 39172 23950
rect 39228 23940 39284 25788
rect 39340 25508 39396 25518
rect 39340 25284 39396 25452
rect 39340 25218 39396 25228
rect 39452 24948 39508 27916
rect 39676 27906 39732 27916
rect 40012 27860 40068 27870
rect 40012 27766 40068 27804
rect 39676 27188 39732 27198
rect 39676 27094 39732 27132
rect 40124 27076 40180 31500
rect 40236 30098 40292 31724
rect 40348 31218 40404 31836
rect 40348 31166 40350 31218
rect 40402 31166 40404 31218
rect 40348 31154 40404 31166
rect 40460 31778 40516 31790
rect 40460 31726 40462 31778
rect 40514 31726 40516 31778
rect 40460 30884 40516 31726
rect 40572 31444 40628 31892
rect 40572 31378 40628 31388
rect 40460 30818 40516 30828
rect 40908 30770 40964 30782
rect 40908 30718 40910 30770
rect 40962 30718 40964 30770
rect 40908 30660 40964 30718
rect 40908 30594 40964 30604
rect 41020 30212 41076 33292
rect 41132 33236 41188 33246
rect 41244 33236 41300 43652
rect 41356 39732 41412 52108
rect 41580 51604 41636 52222
rect 41916 52052 41972 53452
rect 41916 51986 41972 51996
rect 41692 51604 41748 51614
rect 41580 51602 41748 51604
rect 41580 51550 41694 51602
rect 41746 51550 41748 51602
rect 41580 51548 41748 51550
rect 41692 51538 41748 51548
rect 41580 51156 41636 51166
rect 41580 50596 41636 51100
rect 41580 50594 41972 50596
rect 41580 50542 41582 50594
rect 41634 50542 41972 50594
rect 41580 50540 41972 50542
rect 41580 50530 41636 50540
rect 41916 50034 41972 50540
rect 41916 49982 41918 50034
rect 41970 49982 41972 50034
rect 41916 49970 41972 49982
rect 41804 49924 41860 49934
rect 41804 49830 41860 49868
rect 41692 48914 41748 48926
rect 41692 48862 41694 48914
rect 41746 48862 41748 48914
rect 41580 48802 41636 48814
rect 41580 48750 41582 48802
rect 41634 48750 41636 48802
rect 41580 48242 41636 48750
rect 41580 48190 41582 48242
rect 41634 48190 41636 48242
rect 41580 48178 41636 48190
rect 41692 48132 41748 48862
rect 41468 47460 41524 47470
rect 41692 47460 41748 48076
rect 41804 48018 41860 48030
rect 41804 47966 41806 48018
rect 41858 47966 41860 48018
rect 41804 47796 41860 47966
rect 41804 47730 41860 47740
rect 41468 47458 41748 47460
rect 41468 47406 41470 47458
rect 41522 47406 41748 47458
rect 41468 47404 41748 47406
rect 41468 47394 41524 47404
rect 41916 47346 41972 47358
rect 41916 47294 41918 47346
rect 41970 47294 41972 47346
rect 41916 47124 41972 47294
rect 41916 47058 41972 47068
rect 41804 44324 41860 44334
rect 41804 44230 41860 44268
rect 41804 43540 41860 43550
rect 41804 43446 41860 43484
rect 41468 41972 41524 41982
rect 41468 41878 41524 41916
rect 41692 40516 41748 40526
rect 41356 39666 41412 39676
rect 41580 40402 41636 40414
rect 41580 40350 41582 40402
rect 41634 40350 41636 40402
rect 41580 38946 41636 40350
rect 41692 39844 41748 40460
rect 41804 40402 41860 40414
rect 41804 40350 41806 40402
rect 41858 40350 41860 40402
rect 41804 40292 41860 40350
rect 41860 40236 41972 40292
rect 41804 40226 41860 40236
rect 41692 39788 41860 39844
rect 41692 39620 41748 39630
rect 41692 39058 41748 39564
rect 41692 39006 41694 39058
rect 41746 39006 41748 39058
rect 41692 38994 41748 39006
rect 41804 39060 41860 39788
rect 41916 39620 41972 40236
rect 42028 39844 42084 53676
rect 43148 53666 43204 53678
rect 42588 53620 42644 53630
rect 42140 53618 42644 53620
rect 42140 53566 42590 53618
rect 42642 53566 42644 53618
rect 42140 53564 42644 53566
rect 42140 52946 42196 53564
rect 42588 53554 42644 53564
rect 43036 53284 43092 53294
rect 43036 53170 43092 53228
rect 43036 53118 43038 53170
rect 43090 53118 43092 53170
rect 43036 53106 43092 53118
rect 42476 53060 42532 53070
rect 42476 52966 42532 53004
rect 42140 52894 42142 52946
rect 42194 52894 42196 52946
rect 42140 52882 42196 52894
rect 42252 52946 42308 52958
rect 42252 52894 42254 52946
rect 42306 52894 42308 52946
rect 42252 52276 42308 52894
rect 42364 52836 42420 52846
rect 42364 52742 42420 52780
rect 42252 52210 42308 52220
rect 42476 52724 42532 52734
rect 42476 52276 42532 52668
rect 43260 52276 43316 55412
rect 43372 55298 43428 55310
rect 43372 55246 43374 55298
rect 43426 55246 43428 55298
rect 43372 55076 43428 55246
rect 43372 55010 43428 55020
rect 43484 53732 43540 55804
rect 43932 55636 43988 55646
rect 43596 54626 43652 54638
rect 43596 54574 43598 54626
rect 43650 54574 43652 54626
rect 43596 54516 43652 54574
rect 43708 54628 43764 54638
rect 43708 54534 43764 54572
rect 43596 54450 43652 54460
rect 43596 54292 43652 54302
rect 43596 54198 43652 54236
rect 43596 53732 43652 53742
rect 43484 53730 43652 53732
rect 43484 53678 43598 53730
rect 43650 53678 43652 53730
rect 43484 53676 43652 53678
rect 43596 53666 43652 53676
rect 43596 53284 43652 53294
rect 43596 53058 43652 53228
rect 43932 53172 43988 55580
rect 46620 55468 46676 55916
rect 47292 55970 47348 56140
rect 47292 55918 47294 55970
rect 47346 55918 47348 55970
rect 47292 55906 47348 55918
rect 47516 56084 47572 56094
rect 44604 55412 44660 55422
rect 44604 55318 44660 55356
rect 45836 55412 45892 55422
rect 46620 55412 46788 55468
rect 45836 55318 45892 55356
rect 44044 55298 44100 55310
rect 44044 55246 44046 55298
rect 44098 55246 44100 55298
rect 44044 54292 44100 55246
rect 44492 55300 44548 55310
rect 44492 55206 44548 55244
rect 45724 55298 45780 55310
rect 45724 55246 45726 55298
rect 45778 55246 45780 55298
rect 44716 55076 44772 55086
rect 44772 55020 44996 55076
rect 44716 54944 44772 55020
rect 44156 54628 44212 54638
rect 44156 54534 44212 54572
rect 44044 54226 44100 54236
rect 44044 53508 44100 53518
rect 44044 53414 44100 53452
rect 44492 53508 44548 53518
rect 43932 53116 44100 53172
rect 43596 53006 43598 53058
rect 43650 53006 43652 53058
rect 43596 52994 43652 53006
rect 43708 53058 43764 53070
rect 43708 53006 43710 53058
rect 43762 53006 43764 53058
rect 42476 52274 42756 52276
rect 42476 52222 42478 52274
rect 42530 52222 42756 52274
rect 42476 52220 42756 52222
rect 42476 52210 42532 52220
rect 42364 52052 42420 52062
rect 42140 51378 42196 51390
rect 42140 51326 42142 51378
rect 42194 51326 42196 51378
rect 42140 50034 42196 51326
rect 42140 49982 42142 50034
rect 42194 49982 42196 50034
rect 42140 49970 42196 49982
rect 42252 50594 42308 50606
rect 42252 50542 42254 50594
rect 42306 50542 42308 50594
rect 42252 49924 42308 50542
rect 42252 49858 42308 49868
rect 42140 48804 42196 48814
rect 42140 48466 42196 48748
rect 42140 48414 42142 48466
rect 42194 48414 42196 48466
rect 42140 48402 42196 48414
rect 42364 46452 42420 51996
rect 42700 51268 42756 52220
rect 43148 52220 43316 52276
rect 42812 52164 42868 52174
rect 42812 52162 42980 52164
rect 42812 52110 42814 52162
rect 42866 52110 42980 52162
rect 42812 52108 42980 52110
rect 42812 52098 42868 52108
rect 42924 51378 42980 52108
rect 42924 51326 42926 51378
rect 42978 51326 42980 51378
rect 42812 51268 42868 51278
rect 42700 51266 42868 51268
rect 42700 51214 42814 51266
rect 42866 51214 42868 51266
rect 42700 51212 42868 51214
rect 42812 51202 42868 51212
rect 42476 50596 42532 50606
rect 42924 50596 42980 51326
rect 42476 50594 42980 50596
rect 42476 50542 42478 50594
rect 42530 50542 42980 50594
rect 42476 50540 42980 50542
rect 42476 50530 42532 50540
rect 42476 49924 42532 49934
rect 43148 49924 43204 52220
rect 43260 52050 43316 52062
rect 43260 51998 43262 52050
rect 43314 51998 43316 52050
rect 43260 51940 43316 51998
rect 43260 51874 43316 51884
rect 43596 51492 43652 51502
rect 43708 51492 43764 53006
rect 43932 52946 43988 52958
rect 43932 52894 43934 52946
rect 43986 52894 43988 52946
rect 43932 52164 43988 52894
rect 43932 52098 43988 52108
rect 43596 51490 43764 51492
rect 43596 51438 43598 51490
rect 43650 51438 43764 51490
rect 43596 51436 43764 51438
rect 43596 51380 43652 51436
rect 43596 51314 43652 51324
rect 42476 49830 42532 49868
rect 42588 49868 43204 49924
rect 42588 49476 42644 49868
rect 42364 46386 42420 46396
rect 42476 49420 42644 49476
rect 42812 49700 42868 49710
rect 42364 44660 42420 44670
rect 42364 44434 42420 44604
rect 42364 44382 42366 44434
rect 42418 44382 42420 44434
rect 42364 43764 42420 44382
rect 42364 43540 42420 43708
rect 42364 43446 42420 43484
rect 42140 40628 42196 40638
rect 42140 40402 42196 40572
rect 42140 40350 42142 40402
rect 42194 40350 42196 40402
rect 42140 40338 42196 40350
rect 42028 39778 42084 39788
rect 42476 39732 42532 49420
rect 42700 48916 42756 48926
rect 42700 48822 42756 48860
rect 42812 48914 42868 49644
rect 43484 49700 43540 49710
rect 43484 49606 43540 49644
rect 43596 49588 43652 49598
rect 43596 49586 43988 49588
rect 43596 49534 43598 49586
rect 43650 49534 43988 49586
rect 43596 49532 43988 49534
rect 43596 49522 43652 49532
rect 43708 49028 43764 49038
rect 43596 49026 43764 49028
rect 43596 48974 43710 49026
rect 43762 48974 43764 49026
rect 43596 48972 43764 48974
rect 42812 48862 42814 48914
rect 42866 48862 42868 48914
rect 42812 48850 42868 48862
rect 43484 48916 43540 48926
rect 43484 48822 43540 48860
rect 43036 48802 43092 48814
rect 43036 48750 43038 48802
rect 43090 48750 43092 48802
rect 43036 48356 43092 48750
rect 43036 48290 43092 48300
rect 43372 48804 43428 48814
rect 43372 48692 43428 48748
rect 43596 48692 43652 48972
rect 43708 48962 43764 48972
rect 43932 49026 43988 49532
rect 43932 48974 43934 49026
rect 43986 48974 43988 49026
rect 43932 48962 43988 48974
rect 43708 48804 43764 48814
rect 43708 48710 43764 48748
rect 43372 48636 43652 48692
rect 43372 48242 43428 48636
rect 43372 48190 43374 48242
rect 43426 48190 43428 48242
rect 43372 48178 43428 48190
rect 43932 48356 43988 48366
rect 43484 48130 43540 48142
rect 43484 48078 43486 48130
rect 43538 48078 43540 48130
rect 43484 47458 43540 48078
rect 43708 48132 43764 48142
rect 43708 48038 43764 48076
rect 43484 47406 43486 47458
rect 43538 47406 43540 47458
rect 43484 47394 43540 47406
rect 43932 47458 43988 48300
rect 43932 47406 43934 47458
rect 43986 47406 43988 47458
rect 43932 47394 43988 47406
rect 43372 47348 43428 47358
rect 43372 47254 43428 47292
rect 44044 47236 44100 53116
rect 44492 52834 44548 53452
rect 44492 52782 44494 52834
rect 44546 52782 44548 52834
rect 44380 52162 44436 52174
rect 44380 52110 44382 52162
rect 44434 52110 44436 52162
rect 44380 52052 44436 52110
rect 44380 51604 44436 51996
rect 44380 51538 44436 51548
rect 44492 51380 44548 52782
rect 44828 52946 44884 52958
rect 44828 52894 44830 52946
rect 44882 52894 44884 52946
rect 44716 52388 44772 52398
rect 44716 52294 44772 52332
rect 44604 51940 44660 51950
rect 44604 51846 44660 51884
rect 44156 51378 44548 51380
rect 44156 51326 44494 51378
rect 44546 51326 44548 51378
rect 44156 51324 44548 51326
rect 44156 50706 44212 51324
rect 44492 51314 44548 51324
rect 44828 51380 44884 52894
rect 44940 51490 44996 55020
rect 45724 54068 45780 55246
rect 46620 55188 46676 55198
rect 46620 55094 46676 55132
rect 45836 54740 45892 54750
rect 45836 54646 45892 54684
rect 45724 54002 45780 54012
rect 46172 54514 46228 54526
rect 46172 54462 46174 54514
rect 46226 54462 46228 54514
rect 45836 53620 45892 53630
rect 45724 53618 45892 53620
rect 45724 53566 45838 53618
rect 45890 53566 45892 53618
rect 45724 53564 45892 53566
rect 45388 52164 45444 52174
rect 45388 52070 45444 52108
rect 44940 51438 44942 51490
rect 44994 51438 44996 51490
rect 44940 51426 44996 51438
rect 44828 51314 44884 51324
rect 44156 50654 44158 50706
rect 44210 50654 44212 50706
rect 44156 50642 44212 50654
rect 45052 51268 45108 51278
rect 45052 50034 45108 51212
rect 45724 51268 45780 53564
rect 45836 53554 45892 53564
rect 45948 53506 46004 53518
rect 45948 53454 45950 53506
rect 46002 53454 46004 53506
rect 45948 52946 46004 53454
rect 45948 52894 45950 52946
rect 46002 52894 46004 52946
rect 45948 52882 46004 52894
rect 46060 53506 46116 53518
rect 46060 53454 46062 53506
rect 46114 53454 46116 53506
rect 46060 52388 46116 53454
rect 46172 52722 46228 54462
rect 46172 52670 46174 52722
rect 46226 52670 46228 52722
rect 46172 52658 46228 52670
rect 46060 52322 46116 52332
rect 46060 52052 46116 52062
rect 45724 51136 45780 51212
rect 45836 51940 45892 51950
rect 45836 50594 45892 51884
rect 45948 51938 46004 51950
rect 45948 51886 45950 51938
rect 46002 51886 46004 51938
rect 45948 51378 46004 51886
rect 45948 51326 45950 51378
rect 46002 51326 46004 51378
rect 45948 51314 46004 51326
rect 46060 51938 46116 51996
rect 46060 51886 46062 51938
rect 46114 51886 46116 51938
rect 46060 50706 46116 51886
rect 46060 50654 46062 50706
rect 46114 50654 46116 50706
rect 46060 50642 46116 50654
rect 46508 50706 46564 50718
rect 46508 50654 46510 50706
rect 46562 50654 46564 50706
rect 45836 50542 45838 50594
rect 45890 50542 45892 50594
rect 45836 50530 45892 50542
rect 45052 49982 45054 50034
rect 45106 49982 45108 50034
rect 45052 49970 45108 49982
rect 44716 49810 44772 49822
rect 44716 49758 44718 49810
rect 44770 49758 44772 49810
rect 44716 48804 44772 49758
rect 45164 49810 45220 49822
rect 45164 49758 45166 49810
rect 45218 49758 45220 49810
rect 45164 48916 45220 49758
rect 45388 49812 45444 49822
rect 46508 49812 46564 50654
rect 45388 49810 46564 49812
rect 45388 49758 45390 49810
rect 45442 49758 46564 49810
rect 45388 49756 46564 49758
rect 45388 49746 45444 49756
rect 46508 49026 46564 49756
rect 46508 48974 46510 49026
rect 46562 48974 46564 49026
rect 46508 48962 46564 48974
rect 46620 49138 46676 49150
rect 46620 49086 46622 49138
rect 46674 49086 46676 49138
rect 45164 48850 45220 48860
rect 45500 48914 45556 48926
rect 45500 48862 45502 48914
rect 45554 48862 45556 48914
rect 44716 48738 44772 48748
rect 45500 48804 45556 48862
rect 45500 48738 45556 48748
rect 45612 48916 45668 48926
rect 44268 48356 44324 48366
rect 44268 48262 44324 48300
rect 44492 48356 44548 48366
rect 43708 47180 44100 47236
rect 44156 47236 44212 47246
rect 43708 46786 43764 47180
rect 44156 46900 44212 47180
rect 43708 46734 43710 46786
rect 43762 46734 43764 46786
rect 43708 46722 43764 46734
rect 44044 46844 44212 46900
rect 44492 47124 44548 48300
rect 45388 48356 45444 48366
rect 45388 48262 45444 48300
rect 45276 48132 45332 48142
rect 45276 48038 45332 48076
rect 44604 48018 44660 48030
rect 45164 48020 45220 48030
rect 44604 47966 44606 48018
rect 44658 47966 44660 48018
rect 44604 47460 44660 47966
rect 44604 47394 44660 47404
rect 44716 48018 45220 48020
rect 44716 47966 45166 48018
rect 45218 47966 45220 48018
rect 44716 47964 45220 47966
rect 44044 45890 44100 46844
rect 44492 46788 44548 47068
rect 44156 46732 44548 46788
rect 44156 46674 44212 46732
rect 44604 46676 44660 46686
rect 44716 46676 44772 47964
rect 45164 47954 45220 47964
rect 45612 47570 45668 48860
rect 45836 48804 45892 48814
rect 46620 48804 46676 49086
rect 45836 48802 46676 48804
rect 45836 48750 45838 48802
rect 45890 48750 46676 48802
rect 45836 48748 46676 48750
rect 45836 48738 45892 48748
rect 45612 47518 45614 47570
rect 45666 47518 45668 47570
rect 45612 47506 45668 47518
rect 46060 47460 46116 47470
rect 46060 47366 46116 47404
rect 44156 46622 44158 46674
rect 44210 46622 44212 46674
rect 44156 46610 44212 46622
rect 44268 46674 44772 46676
rect 44268 46622 44606 46674
rect 44658 46622 44772 46674
rect 44268 46620 44772 46622
rect 44940 47236 44996 47246
rect 44268 46002 44324 46620
rect 44604 46610 44660 46620
rect 44268 45950 44270 46002
rect 44322 45950 44324 46002
rect 44268 45938 44324 45950
rect 44044 45838 44046 45890
rect 44098 45838 44100 45890
rect 44044 45826 44100 45838
rect 44380 45780 44436 45790
rect 44380 45686 44436 45724
rect 43036 45218 43092 45230
rect 44492 45220 44548 45230
rect 43036 45166 43038 45218
rect 43090 45166 43092 45218
rect 42700 45106 42756 45118
rect 42700 45054 42702 45106
rect 42754 45054 42756 45106
rect 42700 44548 42756 45054
rect 42588 44492 42700 44548
rect 42588 43650 42644 44492
rect 42700 44482 42756 44492
rect 42812 44322 42868 44334
rect 42812 44270 42814 44322
rect 42866 44270 42868 44322
rect 42812 43708 42868 44270
rect 43036 44324 43092 45166
rect 44268 45218 44548 45220
rect 44268 45166 44494 45218
rect 44546 45166 44548 45218
rect 44268 45164 44548 45166
rect 43932 45106 43988 45118
rect 44156 45108 44212 45118
rect 43932 45054 43934 45106
rect 43986 45054 43988 45106
rect 43484 44436 43540 44446
rect 43484 44342 43540 44380
rect 43148 44324 43204 44334
rect 43036 44322 43204 44324
rect 43036 44270 43150 44322
rect 43202 44270 43204 44322
rect 43036 44268 43204 44270
rect 43148 44212 43204 44268
rect 43932 44324 43988 45054
rect 43932 44258 43988 44268
rect 44044 45106 44212 45108
rect 44044 45054 44158 45106
rect 44210 45054 44212 45106
rect 44044 45052 44212 45054
rect 44044 44322 44100 45052
rect 44156 45042 44212 45052
rect 44268 44548 44324 45164
rect 44492 45154 44548 45164
rect 44044 44270 44046 44322
rect 44098 44270 44100 44322
rect 43148 44146 43204 44156
rect 44044 44212 44100 44270
rect 44156 44492 44324 44548
rect 44380 44994 44436 45006
rect 44380 44942 44382 44994
rect 44434 44942 44436 44994
rect 44156 44436 44212 44492
rect 44156 44322 44212 44380
rect 44156 44270 44158 44322
rect 44210 44270 44212 44322
rect 44156 44258 44212 44270
rect 44268 44324 44324 44334
rect 44268 44230 44324 44268
rect 43372 44098 43428 44110
rect 43372 44046 43374 44098
rect 43426 44046 43428 44098
rect 43372 43764 43428 44046
rect 42588 43598 42590 43650
rect 42642 43598 42644 43650
rect 42588 43586 42644 43598
rect 42700 43652 42868 43708
rect 42700 43538 42756 43652
rect 42812 43586 42868 43596
rect 43260 43652 43428 43708
rect 43932 43762 43988 43774
rect 43932 43710 43934 43762
rect 43986 43710 43988 43762
rect 43708 43652 43764 43662
rect 42700 43486 42702 43538
rect 42754 43486 42756 43538
rect 42700 43428 42756 43486
rect 42700 43362 42756 43372
rect 43260 43540 43316 43652
rect 43708 43558 43764 43596
rect 43148 43316 43204 43326
rect 43148 43222 43204 43260
rect 43260 42866 43316 43484
rect 43932 42980 43988 43710
rect 44044 43650 44100 44156
rect 44044 43598 44046 43650
rect 44098 43598 44100 43650
rect 44044 43586 44100 43598
rect 44156 43540 44212 43550
rect 44156 43446 44212 43484
rect 44380 43540 44436 44942
rect 44716 44324 44772 44334
rect 44716 44230 44772 44268
rect 44380 43474 44436 43484
rect 44828 43540 44884 43550
rect 44828 43446 44884 43484
rect 44156 43316 44212 43326
rect 44156 42980 44212 43260
rect 43932 42978 44100 42980
rect 43932 42926 43934 42978
rect 43986 42926 44100 42978
rect 43932 42924 44100 42926
rect 43932 42914 43988 42924
rect 43260 42814 43262 42866
rect 43314 42814 43316 42866
rect 43260 42802 43316 42814
rect 43708 42754 43764 42766
rect 43708 42702 43710 42754
rect 43762 42702 43764 42754
rect 43708 42084 43764 42702
rect 44044 42308 44100 42924
rect 44156 42978 44436 42980
rect 44156 42926 44158 42978
rect 44210 42926 44436 42978
rect 44156 42924 44436 42926
rect 44156 42914 44212 42924
rect 44268 42756 44324 42766
rect 44268 42662 44324 42700
rect 43708 42018 43764 42028
rect 43820 42252 44100 42308
rect 43820 41860 43876 42252
rect 43708 41804 43876 41860
rect 43932 42084 43988 42094
rect 43484 41748 43540 41758
rect 43036 41746 43540 41748
rect 43036 41694 43486 41746
rect 43538 41694 43540 41746
rect 43036 41692 43540 41694
rect 42924 41188 42980 41198
rect 42924 41094 42980 41132
rect 43036 41074 43092 41692
rect 43484 41682 43540 41692
rect 43708 41186 43764 41804
rect 43932 41748 43988 42028
rect 44044 41972 44100 42252
rect 44156 41972 44212 41982
rect 44044 41970 44212 41972
rect 44044 41918 44158 41970
rect 44210 41918 44212 41970
rect 44044 41916 44212 41918
rect 44156 41906 44212 41916
rect 44380 41970 44436 42924
rect 44380 41918 44382 41970
rect 44434 41918 44436 41970
rect 43932 41746 44100 41748
rect 43932 41694 43934 41746
rect 43986 41694 44100 41746
rect 43932 41692 44100 41694
rect 43932 41682 43988 41692
rect 43708 41134 43710 41186
rect 43762 41134 43764 41186
rect 43708 41122 43764 41134
rect 43820 41188 43876 41198
rect 43820 41094 43876 41132
rect 43036 41022 43038 41074
rect 43090 41022 43092 41074
rect 43036 41010 43092 41022
rect 44044 41076 44100 41692
rect 44156 41076 44212 41086
rect 44044 41074 44212 41076
rect 44044 41022 44158 41074
rect 44210 41022 44212 41074
rect 44044 41020 44212 41022
rect 44156 41010 44212 41020
rect 43260 40964 43316 40974
rect 43260 40870 43316 40908
rect 43820 40964 43876 40974
rect 43708 40516 43764 40526
rect 43708 40422 43764 40460
rect 42364 39676 42532 39732
rect 42812 40404 42868 40414
rect 42028 39620 42084 39630
rect 41916 39618 42084 39620
rect 41916 39566 42030 39618
rect 42082 39566 42084 39618
rect 41916 39564 42084 39566
rect 42028 39554 42084 39564
rect 41916 39060 41972 39070
rect 41804 39058 41972 39060
rect 41804 39006 41918 39058
rect 41970 39006 41972 39058
rect 41804 39004 41972 39006
rect 41916 38994 41972 39004
rect 41580 38894 41582 38946
rect 41634 38894 41636 38946
rect 41580 38882 41636 38894
rect 42364 38388 42420 39676
rect 42364 38322 42420 38332
rect 42476 39506 42532 39518
rect 42476 39454 42478 39506
rect 42530 39454 42532 39506
rect 42476 38946 42532 39454
rect 42812 39058 42868 40348
rect 43596 40404 43652 40414
rect 43596 40310 43652 40348
rect 42812 39006 42814 39058
rect 42866 39006 42868 39058
rect 42812 38994 42868 39006
rect 43708 39730 43764 39742
rect 43708 39678 43710 39730
rect 43762 39678 43764 39730
rect 42476 38894 42478 38946
rect 42530 38894 42532 38946
rect 41916 38164 41972 38174
rect 41916 38070 41972 38108
rect 41692 38052 41748 38062
rect 41580 37938 41636 37950
rect 41580 37886 41582 37938
rect 41634 37886 41636 37938
rect 41468 36708 41524 36718
rect 41580 36708 41636 37886
rect 41468 36706 41636 36708
rect 41468 36654 41470 36706
rect 41522 36654 41636 36706
rect 41468 36652 41636 36654
rect 41468 36642 41524 36652
rect 41356 36484 41412 36494
rect 41412 36428 41636 36484
rect 41356 36390 41412 36428
rect 41468 36260 41524 36270
rect 41468 36166 41524 36204
rect 41580 35810 41636 36428
rect 41692 35922 41748 37996
rect 42140 38050 42196 38062
rect 42140 37998 42142 38050
rect 42194 37998 42196 38050
rect 41804 37938 41860 37950
rect 41804 37886 41806 37938
rect 41858 37886 41860 37938
rect 41804 37154 41860 37886
rect 41804 37102 41806 37154
rect 41858 37102 41860 37154
rect 41804 36932 41860 37102
rect 41804 36866 41860 36876
rect 42140 36372 42196 37998
rect 42364 38052 42420 38062
rect 42364 37958 42420 37996
rect 42476 37266 42532 38894
rect 42588 38946 42644 38958
rect 42588 38894 42590 38946
rect 42642 38894 42644 38946
rect 42588 38164 42644 38894
rect 42644 38108 42868 38164
rect 42588 38098 42644 38108
rect 42476 37214 42478 37266
rect 42530 37214 42532 37266
rect 42476 37202 42532 37214
rect 42812 37266 42868 38108
rect 42812 37214 42814 37266
rect 42866 37214 42868 37266
rect 42812 37202 42868 37214
rect 42364 37156 42420 37166
rect 42140 36306 42196 36316
rect 42252 37154 42420 37156
rect 42252 37102 42366 37154
rect 42418 37102 42420 37154
rect 42252 37100 42420 37102
rect 41692 35870 41694 35922
rect 41746 35870 41748 35922
rect 41692 35858 41748 35870
rect 41804 36260 41860 36270
rect 41804 35922 41860 36204
rect 41804 35870 41806 35922
rect 41858 35870 41860 35922
rect 41804 35858 41860 35870
rect 41580 35758 41582 35810
rect 41634 35758 41636 35810
rect 41580 35746 41636 35758
rect 41468 33348 41524 33358
rect 41468 33254 41524 33292
rect 41188 33180 41300 33236
rect 41132 33122 41188 33180
rect 41132 33070 41134 33122
rect 41186 33070 41188 33122
rect 41132 32340 41188 33070
rect 41132 32274 41188 32284
rect 41468 32450 41524 32462
rect 41468 32398 41470 32450
rect 41522 32398 41524 32450
rect 41468 31444 41524 32398
rect 41524 31388 41636 31444
rect 41468 31378 41524 31388
rect 41580 30882 41636 31388
rect 42252 31332 42308 37100
rect 42364 37090 42420 37100
rect 43036 37044 43092 37054
rect 42476 36932 42532 36942
rect 42364 36594 42420 36606
rect 42364 36542 42366 36594
rect 42418 36542 42420 36594
rect 42364 36372 42420 36542
rect 42476 36482 42532 36876
rect 42476 36430 42478 36482
rect 42530 36430 42532 36482
rect 42476 36418 42532 36430
rect 42364 36306 42420 36316
rect 43036 34916 43092 36988
rect 43148 36596 43204 36606
rect 43148 36502 43204 36540
rect 42924 34860 43092 34916
rect 42364 34020 42420 34030
rect 42364 33234 42420 33964
rect 42364 33182 42366 33234
rect 42418 33182 42420 33234
rect 42364 33170 42420 33182
rect 42252 31266 42308 31276
rect 42924 31108 42980 34860
rect 43036 34690 43092 34702
rect 43036 34638 43038 34690
rect 43090 34638 43092 34690
rect 43036 33460 43092 34638
rect 43596 34690 43652 34702
rect 43596 34638 43598 34690
rect 43650 34638 43652 34690
rect 43596 34580 43652 34638
rect 43596 34514 43652 34524
rect 43708 33572 43764 39678
rect 43820 39508 43876 40908
rect 43932 40962 43988 40974
rect 43932 40910 43934 40962
rect 43986 40910 43988 40962
rect 43932 40852 43988 40910
rect 44380 40852 44436 41918
rect 43932 40796 44436 40852
rect 43932 40628 43988 40638
rect 43932 39730 43988 40572
rect 44940 40626 44996 47180
rect 45500 47234 45556 47246
rect 45500 47182 45502 47234
rect 45554 47182 45556 47234
rect 45500 45780 45556 47182
rect 45724 47236 45780 47246
rect 45724 47142 45780 47180
rect 45500 44546 45556 45724
rect 45500 44494 45502 44546
rect 45554 44494 45556 44546
rect 45500 44482 45556 44494
rect 45052 44324 45108 44334
rect 45052 43538 45108 44268
rect 45500 44324 45556 44334
rect 45500 44230 45556 44268
rect 45836 44212 45892 44222
rect 45836 44210 46116 44212
rect 45836 44158 45838 44210
rect 45890 44158 46116 44210
rect 45836 44156 46116 44158
rect 45836 44146 45892 44156
rect 46060 43762 46116 44156
rect 46060 43710 46062 43762
rect 46114 43710 46116 43762
rect 46060 43698 46116 43710
rect 46172 43650 46228 43662
rect 46172 43598 46174 43650
rect 46226 43598 46228 43650
rect 45052 43486 45054 43538
rect 45106 43486 45108 43538
rect 45052 43474 45108 43486
rect 45948 43540 46004 43550
rect 45948 43446 46004 43484
rect 45388 43314 45444 43326
rect 45388 43262 45390 43314
rect 45442 43262 45444 43314
rect 44940 40574 44942 40626
rect 44994 40574 44996 40626
rect 44940 40562 44996 40574
rect 45164 40964 45220 40974
rect 44492 40516 44548 40526
rect 44492 40422 44548 40460
rect 44380 40404 44436 40414
rect 44380 40310 44436 40348
rect 45164 40290 45220 40908
rect 45164 40238 45166 40290
rect 45218 40238 45220 40290
rect 45388 40404 45444 43262
rect 46172 42756 46228 43598
rect 45724 41188 45780 41226
rect 45724 41122 45780 41132
rect 46060 41188 46116 41198
rect 46172 41188 46228 42700
rect 46060 41186 46228 41188
rect 46060 41134 46062 41186
rect 46114 41134 46228 41186
rect 46060 41132 46228 41134
rect 46060 41122 46116 41132
rect 45500 41074 45556 41086
rect 45500 41022 45502 41074
rect 45554 41022 45556 41074
rect 45500 40628 45556 41022
rect 45500 40562 45556 40572
rect 45724 40962 45780 40974
rect 45724 40910 45726 40962
rect 45778 40910 45780 40962
rect 45388 40272 45444 40348
rect 45612 40516 45668 40526
rect 45164 40226 45220 40238
rect 43932 39678 43934 39730
rect 43986 39678 43988 39730
rect 43932 39666 43988 39678
rect 44044 39618 44100 39630
rect 44044 39566 44046 39618
rect 44098 39566 44100 39618
rect 44044 39508 44100 39566
rect 43820 39452 44100 39508
rect 45612 36596 45668 40460
rect 45724 40404 45780 40910
rect 46620 40404 46676 40414
rect 45724 40402 46676 40404
rect 45724 40350 46622 40402
rect 46674 40350 46676 40402
rect 45724 40348 46676 40350
rect 46620 40338 46676 40348
rect 45612 36530 45668 36540
rect 43708 33506 43764 33516
rect 46284 33684 46340 33694
rect 43036 31554 43092 33404
rect 44492 33460 44548 33470
rect 44492 33366 44548 33404
rect 46172 32452 46228 32462
rect 46172 32358 46228 32396
rect 45724 31890 45780 31902
rect 45724 31838 45726 31890
rect 45778 31838 45780 31890
rect 43036 31502 43038 31554
rect 43090 31502 43092 31554
rect 43036 31490 43092 31502
rect 43596 31556 43652 31566
rect 43596 31462 43652 31500
rect 45724 31220 45780 31838
rect 46060 31778 46116 31790
rect 46060 31726 46062 31778
rect 46114 31726 46116 31778
rect 45836 31220 45892 31230
rect 45724 31218 45892 31220
rect 45724 31166 45838 31218
rect 45890 31166 45892 31218
rect 45724 31164 45892 31166
rect 45836 31154 45892 31164
rect 46060 31220 46116 31726
rect 46060 31154 46116 31164
rect 44268 31108 44324 31118
rect 42924 31106 43316 31108
rect 42924 31054 42926 31106
rect 42978 31054 43316 31106
rect 42924 31052 43316 31054
rect 42924 31042 42980 31052
rect 41580 30830 41582 30882
rect 41634 30830 41636 30882
rect 41580 30818 41636 30830
rect 42252 30884 42308 30894
rect 41132 30212 41188 30222
rect 41020 30210 41188 30212
rect 41020 30158 41134 30210
rect 41186 30158 41188 30210
rect 41020 30156 41188 30158
rect 41132 30146 41188 30156
rect 41692 30100 41748 30110
rect 40236 30046 40238 30098
rect 40290 30046 40292 30098
rect 40236 30034 40292 30046
rect 41468 30044 41692 30100
rect 41356 29652 41412 29662
rect 40684 29540 40740 29550
rect 40348 28756 40404 28766
rect 40348 28662 40404 28700
rect 40684 27970 40740 29484
rect 40908 28868 40964 28878
rect 40796 28644 40852 28654
rect 40796 28550 40852 28588
rect 40684 27918 40686 27970
rect 40738 27918 40740 27970
rect 40460 27860 40516 27870
rect 40460 27858 40628 27860
rect 40460 27806 40462 27858
rect 40514 27806 40628 27858
rect 40460 27804 40628 27806
rect 40460 27794 40516 27804
rect 40572 27076 40628 27804
rect 40124 27020 40292 27076
rect 40236 26908 40292 27020
rect 40572 26908 40628 27020
rect 40124 26852 40180 26862
rect 40236 26852 40404 26908
rect 39788 26404 39844 26414
rect 39788 26310 39844 26348
rect 40124 25956 40180 26796
rect 40124 25890 40180 25900
rect 40348 26178 40404 26852
rect 40348 26126 40350 26178
rect 40402 26126 40404 26178
rect 40348 25732 40404 26126
rect 40348 25666 40404 25676
rect 40460 26852 40628 26908
rect 40684 26908 40740 27918
rect 40796 27972 40852 27982
rect 40908 27972 40964 28812
rect 41356 28644 41412 29596
rect 41356 28530 41412 28588
rect 41468 28756 41524 30044
rect 41692 30006 41748 30044
rect 42028 29986 42084 29998
rect 42028 29934 42030 29986
rect 42082 29934 42084 29986
rect 42028 29764 42084 29934
rect 41916 29652 41972 29662
rect 41916 29558 41972 29596
rect 41580 29540 41636 29550
rect 41580 29446 41636 29484
rect 41468 28642 41524 28700
rect 41468 28590 41470 28642
rect 41522 28590 41524 28642
rect 41468 28578 41524 28590
rect 41580 28868 41636 28878
rect 41356 28478 41358 28530
rect 41410 28478 41412 28530
rect 41356 28466 41412 28478
rect 40796 27970 40964 27972
rect 40796 27918 40798 27970
rect 40850 27918 40964 27970
rect 40796 27916 40964 27918
rect 41132 28418 41188 28430
rect 41132 28366 41134 28418
rect 41186 28366 41188 28418
rect 40796 27906 40852 27916
rect 41132 27860 41188 28366
rect 41580 28196 41636 28812
rect 41132 27076 41188 27804
rect 41132 27010 41188 27020
rect 41468 28140 41636 28196
rect 41356 26962 41412 26974
rect 41356 26910 41358 26962
rect 41410 26910 41412 26962
rect 40684 26852 40852 26908
rect 40012 25452 40292 25508
rect 39564 25394 39620 25406
rect 39564 25342 39566 25394
rect 39618 25342 39620 25394
rect 39564 25284 39620 25342
rect 39564 25218 39620 25228
rect 40012 25060 40068 25452
rect 40236 25394 40292 25452
rect 40236 25342 40238 25394
rect 40290 25342 40292 25394
rect 40236 25330 40292 25342
rect 39116 23938 39284 23940
rect 39116 23886 39118 23938
rect 39170 23886 39284 23938
rect 39116 23884 39284 23886
rect 39340 24892 39508 24948
rect 39564 25004 40068 25060
rect 40124 25284 40180 25294
rect 39116 23874 39172 23884
rect 38780 23326 38782 23378
rect 38834 23326 38836 23378
rect 38556 23212 38724 23268
rect 38444 22878 38446 22930
rect 38498 22878 38500 22930
rect 38444 22866 38500 22878
rect 38668 22708 38724 23212
rect 38780 22932 38836 23326
rect 38780 22866 38836 22876
rect 38892 23714 38948 23726
rect 38892 23662 38894 23714
rect 38946 23662 38948 23714
rect 38668 22652 38836 22708
rect 38556 22372 38612 22382
rect 38220 22146 38276 22158
rect 38220 22094 38222 22146
rect 38274 22094 38276 22146
rect 38220 21588 38276 22094
rect 38220 21532 38500 21588
rect 38108 21522 38164 21532
rect 37772 21474 37828 21486
rect 37772 21422 37774 21474
rect 37826 21422 37828 21474
rect 37772 20244 37828 21422
rect 38332 21362 38388 21374
rect 38332 21310 38334 21362
rect 38386 21310 38388 21362
rect 38108 20804 38164 20814
rect 37772 20178 37828 20188
rect 37884 20802 38164 20804
rect 37884 20750 38110 20802
rect 38162 20750 38164 20802
rect 37884 20748 38164 20750
rect 37884 20020 37940 20748
rect 38108 20738 38164 20748
rect 38220 20804 38276 20814
rect 38332 20804 38388 21310
rect 38220 20802 38388 20804
rect 38220 20750 38222 20802
rect 38274 20750 38388 20802
rect 38220 20748 38388 20750
rect 38444 20914 38500 21532
rect 38444 20862 38446 20914
rect 38498 20862 38500 20914
rect 38220 20738 38276 20748
rect 38444 20692 38500 20862
rect 38444 20626 38500 20636
rect 37996 20578 38052 20590
rect 37996 20526 37998 20578
rect 38050 20526 38052 20578
rect 37996 20244 38052 20526
rect 38444 20468 38500 20478
rect 38220 20244 38276 20254
rect 37996 20242 38276 20244
rect 37996 20190 38222 20242
rect 38274 20190 38276 20242
rect 37996 20188 38276 20190
rect 38220 20178 38276 20188
rect 38220 20020 38276 20030
rect 37884 19954 37940 19964
rect 38108 20018 38276 20020
rect 38108 19966 38222 20018
rect 38274 19966 38276 20018
rect 38108 19964 38276 19966
rect 36988 19180 37492 19236
rect 37884 19796 37940 19806
rect 36540 17666 36708 17668
rect 36540 17614 36542 17666
rect 36594 17614 36708 17666
rect 36540 17612 36708 17614
rect 36540 17602 36596 17612
rect 36652 17332 36708 17612
rect 36876 18788 36932 18798
rect 36876 17668 36932 18732
rect 36988 18450 37044 19180
rect 37548 19010 37604 19022
rect 37548 18958 37550 19010
rect 37602 18958 37604 19010
rect 36988 18398 36990 18450
rect 37042 18398 37044 18450
rect 36988 18004 37044 18398
rect 36988 17938 37044 17948
rect 37100 18564 37156 18574
rect 37548 18564 37604 18958
rect 36876 17666 37044 17668
rect 36876 17614 36878 17666
rect 36930 17614 37044 17666
rect 36876 17612 37044 17614
rect 36876 17602 36932 17612
rect 36988 17556 37044 17612
rect 36988 17332 37044 17500
rect 36652 17276 36932 17332
rect 36764 17108 36820 17118
rect 36764 17014 36820 17052
rect 35868 16566 35924 16604
rect 36316 16604 36484 16660
rect 36540 16882 36596 16894
rect 36540 16830 36542 16882
rect 36594 16830 36596 16882
rect 35644 15596 35812 15652
rect 35644 14756 35700 15596
rect 35980 15540 36036 15550
rect 35980 15314 36036 15484
rect 35980 15262 35982 15314
rect 36034 15262 36036 15314
rect 35980 15250 36036 15262
rect 35756 15202 35812 15214
rect 35756 15150 35758 15202
rect 35810 15150 35812 15202
rect 35756 15148 35812 15150
rect 36316 15148 36372 16604
rect 36428 16324 36484 16334
rect 36428 16230 36484 16268
rect 36540 15988 36596 16830
rect 36764 16884 36820 16894
rect 36652 16770 36708 16782
rect 36652 16718 36654 16770
rect 36706 16718 36708 16770
rect 36652 16212 36708 16718
rect 36764 16322 36820 16828
rect 36764 16270 36766 16322
rect 36818 16270 36820 16322
rect 36764 16258 36820 16270
rect 36652 16146 36708 16156
rect 36652 15988 36708 15998
rect 36540 15932 36652 15988
rect 36652 15856 36708 15932
rect 36764 15876 36820 15886
rect 36764 15428 36820 15820
rect 36876 15652 36932 17276
rect 36988 17266 37044 17276
rect 36876 15586 36932 15596
rect 36988 16548 37044 16558
rect 36428 15372 36820 15428
rect 36428 15314 36484 15372
rect 36428 15262 36430 15314
rect 36482 15262 36484 15314
rect 36428 15250 36484 15262
rect 36652 15204 36708 15214
rect 35756 15092 36260 15148
rect 36316 15092 36484 15148
rect 35644 14700 36036 14756
rect 35644 14532 35700 14542
rect 35644 14530 35812 14532
rect 35644 14478 35646 14530
rect 35698 14478 35812 14530
rect 35644 14476 35812 14478
rect 35644 14466 35700 14476
rect 35420 14418 35588 14420
rect 35420 14366 35422 14418
rect 35474 14366 35588 14418
rect 35420 14364 35588 14366
rect 35756 14420 35812 14476
rect 35196 13972 35252 13982
rect 35084 13916 35196 13972
rect 35084 12962 35140 13916
rect 35196 13878 35252 13916
rect 35420 13636 35476 14364
rect 35756 14354 35812 14364
rect 35868 14306 35924 14318
rect 35868 14254 35870 14306
rect 35922 14254 35924 14306
rect 35868 14196 35924 14254
rect 35868 14130 35924 14140
rect 35980 14084 36036 14700
rect 36204 14754 36260 15092
rect 36204 14702 36206 14754
rect 36258 14702 36260 14754
rect 36204 14690 36260 14702
rect 36316 14530 36372 14542
rect 36316 14478 36318 14530
rect 36370 14478 36372 14530
rect 36316 14308 36372 14478
rect 36316 14242 36372 14252
rect 35980 14028 36148 14084
rect 35756 13748 35812 13758
rect 35756 13654 35812 13692
rect 35420 13570 35476 13580
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 36092 13188 36148 14028
rect 36204 13858 36260 13870
rect 36204 13806 36206 13858
rect 36258 13806 36260 13858
rect 36204 13636 36260 13806
rect 36204 13570 36260 13580
rect 36428 13300 36484 15092
rect 36540 13748 36596 13758
rect 36540 13654 36596 13692
rect 36428 13244 36596 13300
rect 35084 12910 35086 12962
rect 35138 12910 35140 12962
rect 35084 12404 35140 12910
rect 35980 13186 36148 13188
rect 35980 13134 36094 13186
rect 36146 13134 36148 13186
rect 35980 13132 36148 13134
rect 35308 12850 35364 12862
rect 35308 12798 35310 12850
rect 35362 12798 35364 12850
rect 35084 12338 35140 12348
rect 35196 12404 35252 12414
rect 35308 12404 35364 12798
rect 35868 12850 35924 12862
rect 35868 12798 35870 12850
rect 35922 12798 35924 12850
rect 35196 12402 35364 12404
rect 35196 12350 35198 12402
rect 35250 12350 35364 12402
rect 35196 12348 35364 12350
rect 35532 12404 35588 12414
rect 35196 12338 35252 12348
rect 35532 12178 35588 12348
rect 35868 12404 35924 12798
rect 35868 12338 35924 12348
rect 35868 12180 35924 12190
rect 35532 12126 35534 12178
rect 35586 12126 35588 12178
rect 35532 12114 35588 12126
rect 35756 12178 35924 12180
rect 35756 12126 35870 12178
rect 35922 12126 35924 12178
rect 35756 12124 35924 12126
rect 35308 11956 35364 11966
rect 35308 11954 35700 11956
rect 35308 11902 35310 11954
rect 35362 11902 35700 11954
rect 35308 11900 35700 11902
rect 35308 11890 35364 11900
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35084 11284 35140 11294
rect 35084 10052 35140 11228
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35084 9986 35140 9996
rect 35532 9940 35588 9950
rect 35644 9940 35700 11900
rect 35756 10724 35812 12124
rect 35868 12114 35924 12124
rect 35980 11956 36036 13132
rect 36092 13122 36148 13132
rect 36428 12738 36484 12750
rect 36428 12686 36430 12738
rect 36482 12686 36484 12738
rect 36428 12292 36484 12686
rect 36428 12226 36484 12236
rect 36204 12180 36260 12190
rect 35868 11900 36036 11956
rect 36092 11956 36148 11966
rect 35868 11282 35924 11900
rect 36092 11862 36148 11900
rect 36204 11506 36260 12124
rect 36204 11454 36206 11506
rect 36258 11454 36260 11506
rect 36204 11442 36260 11454
rect 35868 11230 35870 11282
rect 35922 11230 35924 11282
rect 35868 11218 35924 11230
rect 35980 11284 36036 11294
rect 35980 11190 36036 11228
rect 36092 11170 36148 11182
rect 36092 11118 36094 11170
rect 36146 11118 36148 11170
rect 36092 11060 36148 11118
rect 35868 11004 36148 11060
rect 36316 11170 36372 11182
rect 36316 11118 36318 11170
rect 36370 11118 36372 11170
rect 35868 10724 35924 11004
rect 36316 10948 36372 11118
rect 36540 11172 36596 13244
rect 36652 12852 36708 15148
rect 36764 14642 36820 15372
rect 36764 14590 36766 14642
rect 36818 14590 36820 14642
rect 36764 14578 36820 14590
rect 36876 15092 36932 15102
rect 36876 13188 36932 15036
rect 36988 14308 37044 16492
rect 36988 14242 37044 14252
rect 37100 15540 37156 18508
rect 37212 18508 37604 18564
rect 37212 18228 37268 18508
rect 37548 18452 37604 18508
rect 37884 18674 37940 19740
rect 37996 19012 38052 19022
rect 37996 18918 38052 18956
rect 37884 18622 37886 18674
rect 37938 18622 37940 18674
rect 37884 18564 37940 18622
rect 37884 18498 37940 18508
rect 37548 18386 37604 18396
rect 38108 18452 38164 19964
rect 38220 19954 38276 19964
rect 38332 19236 38388 19246
rect 38332 19142 38388 19180
rect 38220 19010 38276 19022
rect 38220 18958 38222 19010
rect 38274 18958 38276 19010
rect 38220 18564 38276 18958
rect 38220 18498 38276 18508
rect 38108 18386 38164 18396
rect 37436 18340 37492 18350
rect 37436 18246 37492 18284
rect 37996 18340 38052 18350
rect 37212 16660 37268 18172
rect 37436 18004 37492 18014
rect 37436 16996 37492 17948
rect 37660 17556 37716 17566
rect 37660 17462 37716 17500
rect 37548 17442 37604 17454
rect 37548 17390 37550 17442
rect 37602 17390 37604 17442
rect 37548 17108 37604 17390
rect 37548 17042 37604 17052
rect 37660 17332 37716 17342
rect 37436 16902 37492 16940
rect 37212 16594 37268 16604
rect 37436 16660 37492 16670
rect 37100 15204 37156 15484
rect 37100 13972 37156 15148
rect 37212 15764 37268 15774
rect 37212 15148 37268 15708
rect 37436 15540 37492 16604
rect 37324 15484 37492 15540
rect 37660 15540 37716 17276
rect 37772 17220 37828 17230
rect 37772 16100 37828 17164
rect 37996 17108 38052 18284
rect 37996 16994 38052 17052
rect 37996 16942 37998 16994
rect 38050 16942 38052 16994
rect 37996 16930 38052 16942
rect 38108 17220 38164 17230
rect 38108 16994 38164 17164
rect 38108 16942 38110 16994
rect 38162 16942 38164 16994
rect 38108 16930 38164 16942
rect 38220 16996 38276 17006
rect 38220 16902 38276 16940
rect 37772 15986 37828 16044
rect 37772 15934 37774 15986
rect 37826 15934 37828 15986
rect 37772 15922 37828 15934
rect 37884 15988 37940 15998
rect 37772 15540 37828 15550
rect 37660 15538 37828 15540
rect 37660 15486 37774 15538
rect 37826 15486 37828 15538
rect 37660 15484 37828 15486
rect 37324 15426 37380 15484
rect 37772 15474 37828 15484
rect 37324 15374 37326 15426
rect 37378 15374 37380 15426
rect 37324 15362 37380 15374
rect 37212 15092 37380 15148
rect 37212 13972 37268 13982
rect 37100 13970 37268 13972
rect 37100 13918 37214 13970
rect 37266 13918 37268 13970
rect 37100 13916 37268 13918
rect 37212 13906 37268 13916
rect 36876 13122 36932 13132
rect 36652 12796 36932 12852
rect 36652 12628 36708 12638
rect 36652 12402 36708 12572
rect 36652 12350 36654 12402
rect 36706 12350 36708 12402
rect 36652 12338 36708 12350
rect 36764 12404 36820 12414
rect 36764 11508 36820 12348
rect 36540 11106 36596 11116
rect 36652 11506 36820 11508
rect 36652 11454 36766 11506
rect 36818 11454 36820 11506
rect 36652 11452 36820 11454
rect 36316 10882 36372 10892
rect 36652 10836 36708 11452
rect 36764 11442 36820 11452
rect 36428 10780 36708 10836
rect 35756 10722 35924 10724
rect 35756 10670 35758 10722
rect 35810 10670 35924 10722
rect 35756 10668 35924 10670
rect 35756 10658 35812 10668
rect 35756 9940 35812 9950
rect 35644 9884 35756 9940
rect 35532 9846 35588 9884
rect 35756 9846 35812 9884
rect 34972 9772 35252 9828
rect 34748 9762 34804 9772
rect 35196 9492 35252 9772
rect 35868 9716 35924 10668
rect 36092 10724 36148 10734
rect 36428 10724 36484 10780
rect 36092 10722 36484 10724
rect 36092 10670 36094 10722
rect 36146 10670 36484 10722
rect 36092 10668 36484 10670
rect 36092 10658 36148 10668
rect 36316 10386 36372 10668
rect 36876 10612 36932 12796
rect 37324 12740 37380 15092
rect 37436 14644 37492 14654
rect 37884 14644 37940 15932
rect 38108 15986 38164 15998
rect 38108 15934 38110 15986
rect 38162 15934 38164 15986
rect 38108 15540 38164 15934
rect 38108 15148 38164 15484
rect 38220 15652 38276 15662
rect 38220 15538 38276 15596
rect 38220 15486 38222 15538
rect 38274 15486 38276 15538
rect 38220 15316 38276 15486
rect 38220 15250 38276 15260
rect 38444 15148 38500 20412
rect 38556 20018 38612 22316
rect 38668 22148 38724 22158
rect 38668 22054 38724 22092
rect 38780 22146 38836 22652
rect 38892 22372 38948 23662
rect 38892 22306 38948 22316
rect 39228 22260 39284 22270
rect 39228 22166 39284 22204
rect 38780 22094 38782 22146
rect 38834 22094 38836 22146
rect 38780 21812 38836 22094
rect 39004 22148 39060 22158
rect 39340 22148 39396 24892
rect 39452 24724 39508 24734
rect 39564 24724 39620 25004
rect 40124 24834 40180 25228
rect 40348 25172 40404 25182
rect 40460 25172 40516 26852
rect 40796 26850 40852 26852
rect 40796 26798 40798 26850
rect 40850 26798 40852 26850
rect 40572 26180 40628 26190
rect 40572 25506 40628 26124
rect 40572 25454 40574 25506
rect 40626 25454 40628 25506
rect 40572 25442 40628 25454
rect 40684 26178 40740 26190
rect 40684 26126 40686 26178
rect 40738 26126 40740 26178
rect 40684 25508 40740 26126
rect 40796 25732 40852 26798
rect 41356 26180 41412 26910
rect 41468 26516 41524 28140
rect 41580 27972 41636 27982
rect 41580 27878 41636 27916
rect 41916 27860 41972 27870
rect 41916 27766 41972 27804
rect 41916 27412 41972 27422
rect 41580 27076 41636 27114
rect 41580 27010 41636 27020
rect 41916 27074 41972 27356
rect 41916 27022 41918 27074
rect 41970 27022 41972 27074
rect 41580 26852 41636 26862
rect 41580 26850 41748 26852
rect 41580 26798 41582 26850
rect 41634 26798 41748 26850
rect 41580 26796 41748 26798
rect 41580 26786 41636 26796
rect 41580 26516 41636 26526
rect 41468 26514 41636 26516
rect 41468 26462 41582 26514
rect 41634 26462 41636 26514
rect 41468 26460 41636 26462
rect 41580 26450 41636 26460
rect 41356 26114 41412 26124
rect 41132 25844 41188 25854
rect 40796 25676 41076 25732
rect 40684 25442 40740 25452
rect 40908 25396 40964 25406
rect 40460 25116 40740 25172
rect 40348 24948 40404 25116
rect 40572 24948 40628 24958
rect 40348 24946 40628 24948
rect 40348 24894 40574 24946
rect 40626 24894 40628 24946
rect 40348 24892 40628 24894
rect 40124 24782 40126 24834
rect 40178 24782 40180 24834
rect 40124 24770 40180 24782
rect 40572 24836 40628 24892
rect 40572 24770 40628 24780
rect 39452 24722 39620 24724
rect 39452 24670 39454 24722
rect 39506 24670 39620 24722
rect 39452 24668 39620 24670
rect 39676 24722 39732 24734
rect 39676 24670 39678 24722
rect 39730 24670 39732 24722
rect 39452 23938 39508 24668
rect 39452 23886 39454 23938
rect 39506 23886 39508 23938
rect 39452 22260 39508 23886
rect 39676 23492 39732 24670
rect 39900 24722 39956 24734
rect 39900 24670 39902 24722
rect 39954 24670 39956 24722
rect 39788 24610 39844 24622
rect 39788 24558 39790 24610
rect 39842 24558 39844 24610
rect 39788 24052 39844 24558
rect 39788 23986 39844 23996
rect 39900 24162 39956 24670
rect 39900 24110 39902 24162
rect 39954 24110 39956 24162
rect 39564 23380 39620 23390
rect 39676 23380 39732 23436
rect 39564 23378 39732 23380
rect 39564 23326 39566 23378
rect 39618 23326 39732 23378
rect 39564 23324 39732 23326
rect 39564 23314 39620 23324
rect 39900 22370 39956 24110
rect 40236 23938 40292 23950
rect 40236 23886 40238 23938
rect 40290 23886 40292 23938
rect 40236 23604 40292 23886
rect 40236 23538 40292 23548
rect 40460 23938 40516 23950
rect 40460 23886 40462 23938
rect 40514 23886 40516 23938
rect 40460 23380 40516 23886
rect 40684 23548 40740 25116
rect 40908 23938 40964 25340
rect 40908 23886 40910 23938
rect 40962 23886 40964 23938
rect 40908 23874 40964 23886
rect 41020 25172 41076 25676
rect 41132 25396 41188 25788
rect 41132 25302 41188 25340
rect 41244 25282 41300 25294
rect 41468 25284 41524 25294
rect 41244 25230 41246 25282
rect 41298 25230 41300 25282
rect 41244 25172 41300 25230
rect 41020 25116 41300 25172
rect 41356 25282 41524 25284
rect 41356 25230 41470 25282
rect 41522 25230 41524 25282
rect 41356 25228 41524 25230
rect 41020 23716 41076 25116
rect 41244 23940 41300 23950
rect 41356 23940 41412 25228
rect 41468 25218 41524 25228
rect 41468 24612 41524 24622
rect 41468 24518 41524 24556
rect 41692 23940 41748 26796
rect 41804 25956 41860 25966
rect 41804 25618 41860 25900
rect 41804 25566 41806 25618
rect 41858 25566 41860 25618
rect 41804 25554 41860 25566
rect 41916 24724 41972 27022
rect 42028 26740 42084 29708
rect 42028 26674 42084 26684
rect 42140 26180 42196 26190
rect 42140 26086 42196 26124
rect 42252 25284 42308 30828
rect 43260 30322 43316 31052
rect 44268 31106 44548 31108
rect 44268 31054 44270 31106
rect 44322 31054 44548 31106
rect 44268 31052 44548 31054
rect 44268 31042 44324 31052
rect 44044 30994 44100 31006
rect 44044 30942 44046 30994
rect 44098 30942 44100 30994
rect 43260 30270 43262 30322
rect 43314 30270 43316 30322
rect 43260 30258 43316 30270
rect 43820 30772 43876 30782
rect 42364 30212 42420 30222
rect 42364 29652 42420 30156
rect 42364 29520 42420 29596
rect 42476 30100 42532 30110
rect 42476 28866 42532 30044
rect 43820 30100 43876 30716
rect 43932 30212 43988 30222
rect 43932 30118 43988 30156
rect 43708 29764 43764 29774
rect 43260 29652 43316 29662
rect 43260 29558 43316 29596
rect 43708 29650 43764 29708
rect 43708 29598 43710 29650
rect 43762 29598 43764 29650
rect 43708 29586 43764 29598
rect 42924 29540 42980 29550
rect 42476 28814 42478 28866
rect 42530 28814 42532 28866
rect 42476 28802 42532 28814
rect 42700 29538 42980 29540
rect 42700 29486 42926 29538
rect 42978 29486 42980 29538
rect 42700 29484 42980 29486
rect 42700 28868 42756 29484
rect 42924 29474 42980 29484
rect 42588 28642 42644 28654
rect 42588 28590 42590 28642
rect 42642 28590 42644 28642
rect 42476 28420 42532 28430
rect 42364 28418 42532 28420
rect 42364 28366 42478 28418
rect 42530 28366 42532 28418
rect 42364 28364 42532 28366
rect 42364 27188 42420 28364
rect 42476 28354 42532 28364
rect 42588 28420 42644 28590
rect 42476 27972 42532 27982
rect 42588 27972 42644 28364
rect 42476 27970 42644 27972
rect 42476 27918 42478 27970
rect 42530 27918 42644 27970
rect 42476 27916 42644 27918
rect 42476 27906 42532 27916
rect 42700 27858 42756 28812
rect 42700 27806 42702 27858
rect 42754 27806 42756 27858
rect 42588 27746 42644 27758
rect 42588 27694 42590 27746
rect 42642 27694 42644 27746
rect 42588 27412 42644 27694
rect 42700 27748 42756 27806
rect 42700 27682 42756 27692
rect 42812 28642 42868 28654
rect 43820 28644 43876 30044
rect 44044 29764 44100 30942
rect 44492 30996 44548 31052
rect 44492 30210 44548 30940
rect 45388 30994 45444 31006
rect 45388 30942 45390 30994
rect 45442 30942 45444 30994
rect 44492 30158 44494 30210
rect 44546 30158 44548 30210
rect 44156 30100 44212 30110
rect 44156 30006 44212 30044
rect 44044 29698 44100 29708
rect 44268 29986 44324 29998
rect 44268 29934 44270 29986
rect 44322 29934 44324 29986
rect 44268 29428 44324 29934
rect 44380 29652 44436 29662
rect 44492 29652 44548 30158
rect 44716 30882 44772 30894
rect 44716 30830 44718 30882
rect 44770 30830 44772 30882
rect 44716 29764 44772 30830
rect 45388 30884 45444 30942
rect 45724 30996 45780 31006
rect 45724 30902 45780 30940
rect 45948 30994 46004 31006
rect 45948 30942 45950 30994
rect 46002 30942 46004 30994
rect 45388 30818 45444 30828
rect 45388 30100 45444 30110
rect 45388 29988 45444 30044
rect 44716 29698 44772 29708
rect 45276 29986 45444 29988
rect 45276 29934 45390 29986
rect 45442 29934 45444 29986
rect 45276 29932 45444 29934
rect 44604 29652 44660 29662
rect 44492 29650 44660 29652
rect 44492 29598 44606 29650
rect 44658 29598 44660 29650
rect 44492 29596 44660 29598
rect 44380 29558 44436 29596
rect 44604 29586 44660 29596
rect 44828 29540 44884 29550
rect 44828 29446 44884 29484
rect 42812 28590 42814 28642
rect 42866 28590 42868 28642
rect 42812 27636 42868 28590
rect 43708 28588 43876 28644
rect 44156 29372 44324 29428
rect 43484 28532 43540 28542
rect 42812 27570 42868 27580
rect 42924 28420 42980 28430
rect 42588 27346 42644 27356
rect 42364 27132 42868 27188
rect 42364 26964 42420 26974
rect 42364 26870 42420 26908
rect 42700 26962 42756 26974
rect 42700 26910 42702 26962
rect 42754 26910 42756 26962
rect 42588 26852 42644 26862
rect 42588 26758 42644 26796
rect 42252 25190 42308 25228
rect 42364 26740 42420 26750
rect 42364 26180 42420 26684
rect 42588 26180 42644 26190
rect 42700 26180 42756 26910
rect 42364 26178 42756 26180
rect 42364 26126 42590 26178
rect 42642 26126 42756 26178
rect 42364 26124 42756 26126
rect 42252 24724 42308 24734
rect 41916 24722 42308 24724
rect 41916 24670 42254 24722
rect 42306 24670 42308 24722
rect 41916 24668 42308 24670
rect 42252 24658 42308 24668
rect 42364 24500 42420 26124
rect 42588 26114 42644 26124
rect 42588 24836 42644 24846
rect 42252 24444 42420 24500
rect 42476 24500 42532 24510
rect 42588 24500 42644 24780
rect 42812 24724 42868 27132
rect 42924 26964 42980 28364
rect 43036 27972 43092 27982
rect 43036 27634 43092 27916
rect 43372 27972 43428 27982
rect 43036 27582 43038 27634
rect 43090 27582 43092 27634
rect 43036 27570 43092 27582
rect 43148 27860 43204 27870
rect 42924 26898 42980 26908
rect 43148 27186 43204 27804
rect 43148 27134 43150 27186
rect 43202 27134 43204 27186
rect 43148 26404 43204 27134
rect 43260 27858 43316 27870
rect 43260 27806 43262 27858
rect 43314 27806 43316 27858
rect 43260 26964 43316 27806
rect 43260 26898 43316 26908
rect 43372 26514 43428 27916
rect 43372 26462 43374 26514
rect 43426 26462 43428 26514
rect 43372 26450 43428 26462
rect 43148 26338 43204 26348
rect 43148 25620 43204 25630
rect 43148 25526 43204 25564
rect 43260 25508 43316 25518
rect 43036 25396 43092 25406
rect 43036 25394 43204 25396
rect 43036 25342 43038 25394
rect 43090 25342 43204 25394
rect 43036 25340 43204 25342
rect 43036 25330 43092 25340
rect 42924 24724 42980 24734
rect 42812 24722 42980 24724
rect 42812 24670 42926 24722
rect 42978 24670 42980 24722
rect 42812 24668 42980 24670
rect 42476 24498 42644 24500
rect 42476 24446 42478 24498
rect 42530 24446 42644 24498
rect 42476 24444 42644 24446
rect 41916 23940 41972 23950
rect 41244 23938 41636 23940
rect 41244 23886 41246 23938
rect 41298 23886 41636 23938
rect 41244 23884 41636 23886
rect 41692 23938 41972 23940
rect 41692 23886 41918 23938
rect 41970 23886 41972 23938
rect 41692 23884 41972 23886
rect 41244 23874 41300 23884
rect 41020 23650 41076 23660
rect 41132 23714 41188 23726
rect 41132 23662 41134 23714
rect 41186 23662 41188 23714
rect 40684 23492 41076 23548
rect 40460 23314 40516 23324
rect 40124 23154 40180 23166
rect 40124 23102 40126 23154
rect 40178 23102 40180 23154
rect 40012 22484 40068 22494
rect 40012 22390 40068 22428
rect 39900 22318 39902 22370
rect 39954 22318 39956 22370
rect 39900 22306 39956 22318
rect 39452 22204 39732 22260
rect 39004 22146 39172 22148
rect 39004 22094 39006 22146
rect 39058 22094 39172 22146
rect 39004 22092 39172 22094
rect 39004 22082 39060 22092
rect 39116 21812 39172 22092
rect 39340 22082 39396 22092
rect 39452 21812 39508 21822
rect 39116 21756 39396 21812
rect 38780 21746 38836 21756
rect 38668 21700 38724 21710
rect 38668 21476 38724 21644
rect 39340 21698 39396 21756
rect 39452 21718 39508 21756
rect 39340 21646 39342 21698
rect 39394 21646 39396 21698
rect 38780 21476 38836 21486
rect 38668 21474 38836 21476
rect 38668 21422 38782 21474
rect 38834 21422 38836 21474
rect 38668 21420 38836 21422
rect 38780 21140 38836 21420
rect 38780 21074 38836 21084
rect 39340 21026 39396 21646
rect 39564 21698 39620 21710
rect 39564 21646 39566 21698
rect 39618 21646 39620 21698
rect 39340 20974 39342 21026
rect 39394 20974 39396 21026
rect 39340 20962 39396 20974
rect 39452 21588 39508 21598
rect 39452 20914 39508 21532
rect 39452 20862 39454 20914
rect 39506 20862 39508 20914
rect 39452 20850 39508 20862
rect 39564 21476 39620 21646
rect 38668 20804 38724 20814
rect 38668 20710 38724 20748
rect 38892 20802 38948 20814
rect 38892 20750 38894 20802
rect 38946 20750 38948 20802
rect 38556 19966 38558 20018
rect 38610 19966 38612 20018
rect 38556 19954 38612 19966
rect 38780 20018 38836 20030
rect 38780 19966 38782 20018
rect 38834 19966 38836 20018
rect 38780 19572 38836 19966
rect 38892 19684 38948 20750
rect 39340 20804 39396 20814
rect 39004 20132 39060 20142
rect 39004 20038 39060 20076
rect 39340 19908 39396 20748
rect 39452 20356 39508 20366
rect 39452 20130 39508 20300
rect 39452 20078 39454 20130
rect 39506 20078 39508 20130
rect 39452 20066 39508 20078
rect 39564 20132 39620 21420
rect 39564 20066 39620 20076
rect 39340 19852 39620 19908
rect 38892 19628 39172 19684
rect 38780 19506 38836 19516
rect 38892 19236 38948 19246
rect 38780 19012 38836 19022
rect 38668 19010 38836 19012
rect 38668 18958 38782 19010
rect 38834 18958 38836 19010
rect 38668 18956 38836 18958
rect 38108 15092 38276 15148
rect 37436 14642 37940 14644
rect 37436 14590 37438 14642
rect 37490 14590 37886 14642
rect 37938 14590 37940 14642
rect 37436 14588 37940 14590
rect 37436 14578 37492 14588
rect 37884 14578 37940 14588
rect 37548 14308 37604 14318
rect 37548 13074 37604 14252
rect 38108 13858 38164 13870
rect 38108 13806 38110 13858
rect 38162 13806 38164 13858
rect 38108 13748 38164 13806
rect 37548 13022 37550 13074
rect 37602 13022 37604 13074
rect 37548 13010 37604 13022
rect 37996 13522 38052 13534
rect 37996 13470 37998 13522
rect 38050 13470 38052 13522
rect 37996 12964 38052 13470
rect 37996 12898 38052 12908
rect 37884 12740 37940 12750
rect 38108 12740 38164 13692
rect 38220 13076 38276 15092
rect 38332 15092 38500 15148
rect 38556 18564 38612 18574
rect 38556 17554 38612 18508
rect 38668 18228 38724 18956
rect 38780 18946 38836 18956
rect 38892 18788 38948 19180
rect 39116 19124 39172 19628
rect 39340 19460 39396 19470
rect 39116 19030 39172 19068
rect 39228 19348 39284 19358
rect 39004 19012 39060 19022
rect 39004 18918 39060 18956
rect 38780 18732 38948 18788
rect 38780 18562 38836 18732
rect 38780 18510 38782 18562
rect 38834 18510 38836 18562
rect 38780 18498 38836 18510
rect 39004 18676 39060 18686
rect 39228 18676 39284 19292
rect 39004 18674 39284 18676
rect 39004 18622 39006 18674
rect 39058 18622 39284 18674
rect 39004 18620 39284 18622
rect 39340 18674 39396 19404
rect 39564 19346 39620 19852
rect 39564 19294 39566 19346
rect 39618 19294 39620 19346
rect 39564 18900 39620 19294
rect 39676 19236 39732 22204
rect 39900 22148 39956 22158
rect 40124 22148 40180 23102
rect 40348 23156 40404 23166
rect 40348 23062 40404 23100
rect 40572 23154 40628 23166
rect 40572 23102 40574 23154
rect 40626 23102 40628 23154
rect 40460 23042 40516 23054
rect 40460 22990 40462 23042
rect 40514 22990 40516 23042
rect 40348 22370 40404 22382
rect 40348 22318 40350 22370
rect 40402 22318 40404 22370
rect 40236 22260 40292 22270
rect 40236 22166 40292 22204
rect 39956 22092 40068 22148
rect 39900 22082 39956 22092
rect 39788 20580 39844 20590
rect 39788 20578 39956 20580
rect 39788 20526 39790 20578
rect 39842 20526 39956 20578
rect 39788 20524 39956 20526
rect 39788 20514 39844 20524
rect 39900 20244 39956 20524
rect 39900 19906 39956 20188
rect 39900 19854 39902 19906
rect 39954 19854 39956 19906
rect 39900 19796 39956 19854
rect 39900 19730 39956 19740
rect 40012 19348 40068 22092
rect 40012 19282 40068 19292
rect 39676 19170 39732 19180
rect 40012 19124 40068 19134
rect 40012 19030 40068 19068
rect 40124 18900 40180 22092
rect 40236 21812 40292 21822
rect 40348 21812 40404 22318
rect 40460 22036 40516 22990
rect 40572 22484 40628 23102
rect 40572 22418 40628 22428
rect 40796 23154 40852 23166
rect 40796 23102 40798 23154
rect 40850 23102 40852 23154
rect 40796 23044 40852 23102
rect 40460 21970 40516 21980
rect 40684 22372 40740 22382
rect 40292 21756 40404 21812
rect 40236 21680 40292 21756
rect 40460 21588 40516 21598
rect 40460 21494 40516 21532
rect 40348 21474 40404 21486
rect 40348 21422 40350 21474
rect 40402 21422 40404 21474
rect 40236 21026 40292 21038
rect 40236 20974 40238 21026
rect 40290 20974 40292 21026
rect 40236 20914 40292 20974
rect 40236 20862 40238 20914
rect 40290 20862 40292 20914
rect 40236 20356 40292 20862
rect 40348 20580 40404 21422
rect 40684 21140 40740 22316
rect 40796 21588 40852 22988
rect 40908 22260 40964 22270
rect 40908 22166 40964 22204
rect 40908 21588 40964 21598
rect 40796 21586 40964 21588
rect 40796 21534 40910 21586
rect 40962 21534 40964 21586
rect 40796 21532 40964 21534
rect 40908 21364 40964 21532
rect 40908 21298 40964 21308
rect 40684 21084 40964 21140
rect 40908 20802 40964 21084
rect 40908 20750 40910 20802
rect 40962 20750 40964 20802
rect 40908 20738 40964 20750
rect 40348 20514 40404 20524
rect 40908 20356 40964 20366
rect 40236 20300 40516 20356
rect 40348 20132 40404 20142
rect 40460 20132 40516 20300
rect 40796 20132 40852 20142
rect 40460 20130 40852 20132
rect 40460 20078 40798 20130
rect 40850 20078 40852 20130
rect 40460 20076 40852 20078
rect 40348 20038 40404 20076
rect 39564 18834 39620 18844
rect 39900 18844 40180 18900
rect 40684 19572 40740 19582
rect 39900 18788 39956 18844
rect 39340 18622 39342 18674
rect 39394 18622 39396 18674
rect 39004 18564 39060 18620
rect 39004 18498 39060 18508
rect 39228 18450 39284 18462
rect 39228 18398 39230 18450
rect 39282 18398 39284 18450
rect 38892 18340 38948 18350
rect 38668 18172 38836 18228
rect 38556 17502 38558 17554
rect 38610 17502 38612 17554
rect 38556 15092 38612 17502
rect 38668 17444 38724 17454
rect 38668 17350 38724 17388
rect 38780 16996 38836 18172
rect 38892 17666 38948 18284
rect 39116 18338 39172 18350
rect 39116 18286 39118 18338
rect 39170 18286 39172 18338
rect 39116 18228 39172 18286
rect 39228 18340 39284 18398
rect 39228 18274 39284 18284
rect 39116 18162 39172 18172
rect 39340 18004 39396 18622
rect 39116 17948 39396 18004
rect 39676 18732 39956 18788
rect 39004 17892 39060 17902
rect 39004 17798 39060 17836
rect 38892 17614 38894 17666
rect 38946 17614 38948 17666
rect 38892 17602 38948 17614
rect 38780 16930 38836 16940
rect 38668 16660 38724 16670
rect 38668 16658 38948 16660
rect 38668 16606 38670 16658
rect 38722 16606 38948 16658
rect 38668 16604 38948 16606
rect 38668 16594 38724 16604
rect 38668 16100 38724 16110
rect 38668 16006 38724 16044
rect 38892 15202 38948 16604
rect 39116 15652 39172 17948
rect 39228 17668 39284 17678
rect 39676 17668 39732 18732
rect 40124 18676 40180 18686
rect 39900 18674 40180 18676
rect 39900 18622 40126 18674
rect 40178 18622 40180 18674
rect 39900 18620 40180 18622
rect 39900 18340 39956 18620
rect 40124 18610 40180 18620
rect 40236 18562 40292 18574
rect 40236 18510 40238 18562
rect 40290 18510 40292 18562
rect 39900 18274 39956 18284
rect 40012 18452 40068 18462
rect 40012 18228 40068 18396
rect 40012 18226 40180 18228
rect 40012 18174 40014 18226
rect 40066 18174 40180 18226
rect 40012 18172 40180 18174
rect 40012 18162 40068 18172
rect 39900 17892 39956 17902
rect 39900 17798 39956 17836
rect 39676 17612 39956 17668
rect 39228 17574 39284 17612
rect 39900 17444 39956 17612
rect 40012 17444 40068 17454
rect 39900 17442 40068 17444
rect 39900 17390 40014 17442
rect 40066 17390 40068 17442
rect 39900 17388 40068 17390
rect 40124 17444 40180 18172
rect 40236 18116 40292 18510
rect 40236 18050 40292 18060
rect 40348 18452 40404 18462
rect 40684 18452 40740 19516
rect 40796 19460 40852 20076
rect 40796 19394 40852 19404
rect 40796 19010 40852 19022
rect 40796 18958 40798 19010
rect 40850 18958 40852 19010
rect 40796 18676 40852 18958
rect 40796 18610 40852 18620
rect 40796 18452 40852 18462
rect 40684 18450 40852 18452
rect 40684 18398 40798 18450
rect 40850 18398 40852 18450
rect 40684 18396 40852 18398
rect 40236 17668 40292 17678
rect 40348 17668 40404 18396
rect 40796 18386 40852 18396
rect 40236 17666 40404 17668
rect 40236 17614 40238 17666
rect 40290 17614 40404 17666
rect 40236 17612 40404 17614
rect 40236 17602 40292 17612
rect 40460 17556 40516 17566
rect 40124 17388 40292 17444
rect 39900 17220 39956 17230
rect 39340 17106 39396 17118
rect 39340 17054 39342 17106
rect 39394 17054 39396 17106
rect 39340 16100 39396 17054
rect 39676 16996 39732 17006
rect 39452 16884 39508 16894
rect 39452 16790 39508 16828
rect 39340 16034 39396 16044
rect 39676 16098 39732 16940
rect 39900 16882 39956 17164
rect 39900 16830 39902 16882
rect 39954 16830 39956 16882
rect 39900 16818 39956 16830
rect 39676 16046 39678 16098
rect 39730 16046 39732 16098
rect 39676 16034 39732 16046
rect 39788 15876 39844 15886
rect 39116 15586 39172 15596
rect 39340 15874 39844 15876
rect 39340 15822 39790 15874
rect 39842 15822 39844 15874
rect 39340 15820 39844 15822
rect 39340 15314 39396 15820
rect 39788 15810 39844 15820
rect 39340 15262 39342 15314
rect 39394 15262 39396 15314
rect 39340 15250 39396 15262
rect 39564 15428 39620 15438
rect 39564 15314 39620 15372
rect 39564 15262 39566 15314
rect 39618 15262 39620 15314
rect 39564 15250 39620 15262
rect 38892 15150 38894 15202
rect 38946 15150 38948 15202
rect 38892 15138 38948 15150
rect 38332 13748 38388 15092
rect 38556 15036 38724 15092
rect 38444 14420 38500 14430
rect 38444 14308 38500 14364
rect 38444 14306 38612 14308
rect 38444 14254 38446 14306
rect 38498 14254 38612 14306
rect 38444 14252 38612 14254
rect 38444 14242 38500 14252
rect 38332 13746 38500 13748
rect 38332 13694 38334 13746
rect 38386 13694 38500 13746
rect 38332 13692 38500 13694
rect 38332 13682 38388 13692
rect 38332 13076 38388 13086
rect 38220 13074 38388 13076
rect 38220 13022 38334 13074
rect 38386 13022 38388 13074
rect 38220 13020 38388 13022
rect 38332 13010 38388 13020
rect 38444 12964 38500 13692
rect 38444 12898 38500 12908
rect 37324 12684 37492 12740
rect 37100 12292 37156 12302
rect 37100 12198 37156 12236
rect 37212 12180 37268 12190
rect 37212 12086 37268 12124
rect 37324 12178 37380 12190
rect 37324 12126 37326 12178
rect 37378 12126 37380 12178
rect 37324 11956 37380 12126
rect 37100 10948 37156 10958
rect 37100 10834 37156 10892
rect 37100 10782 37102 10834
rect 37154 10782 37156 10834
rect 37100 10770 37156 10782
rect 36652 10556 36932 10612
rect 37324 10612 37380 11900
rect 37436 10834 37492 12684
rect 37884 12738 38164 12740
rect 37884 12686 37886 12738
rect 37938 12686 38164 12738
rect 37884 12684 38164 12686
rect 37884 12180 37940 12684
rect 37884 12114 37940 12124
rect 37548 11844 37604 11854
rect 37548 11282 37604 11788
rect 38556 11844 38612 14252
rect 38668 13972 38724 15036
rect 38780 15090 38836 15102
rect 38780 15038 38782 15090
rect 38834 15038 38836 15090
rect 38780 14196 38836 15038
rect 39228 14532 39284 14542
rect 39228 14438 39284 14476
rect 39004 14418 39060 14430
rect 39004 14366 39006 14418
rect 39058 14366 39060 14418
rect 38780 14130 38836 14140
rect 38892 14308 38948 14318
rect 38668 13906 38724 13916
rect 38892 13860 38948 14252
rect 39004 13972 39060 14366
rect 39004 13906 39060 13916
rect 39452 14306 39508 14318
rect 39452 14254 39454 14306
rect 39506 14254 39508 14306
rect 39452 14084 39508 14254
rect 39564 14308 39620 14318
rect 39564 14214 39620 14252
rect 40012 14196 40068 17388
rect 40124 15986 40180 15998
rect 40124 15934 40126 15986
rect 40178 15934 40180 15986
rect 40124 14980 40180 15934
rect 40236 15764 40292 17388
rect 40460 17106 40516 17500
rect 40684 17442 40740 17454
rect 40684 17390 40686 17442
rect 40738 17390 40740 17442
rect 40684 17220 40740 17390
rect 40684 17154 40740 17164
rect 40460 17054 40462 17106
rect 40514 17054 40516 17106
rect 40460 17042 40516 17054
rect 40684 16996 40740 17006
rect 40684 16098 40740 16940
rect 40684 16046 40686 16098
rect 40738 16046 40740 16098
rect 40684 16034 40740 16046
rect 40796 16996 40852 17006
rect 40908 16996 40964 20300
rect 40796 16994 40964 16996
rect 40796 16942 40798 16994
rect 40850 16942 40964 16994
rect 40796 16940 40964 16942
rect 40796 15986 40852 16940
rect 40796 15934 40798 15986
rect 40850 15934 40852 15986
rect 40796 15922 40852 15934
rect 40236 15698 40292 15708
rect 40348 15652 40404 15662
rect 40348 15538 40404 15596
rect 40348 15486 40350 15538
rect 40402 15486 40404 15538
rect 40348 15474 40404 15486
rect 40796 15316 40852 15326
rect 40684 15314 40852 15316
rect 40684 15262 40798 15314
rect 40850 15262 40852 15314
rect 40684 15260 40852 15262
rect 40124 14914 40180 14924
rect 40236 15090 40292 15102
rect 40236 15038 40238 15090
rect 40290 15038 40292 15090
rect 40236 14530 40292 15038
rect 40684 15092 40740 15260
rect 40796 15250 40852 15260
rect 40684 14644 40740 15036
rect 40236 14478 40238 14530
rect 40290 14478 40292 14530
rect 40236 14466 40292 14478
rect 40348 14588 40740 14644
rect 41020 15090 41076 23492
rect 41132 23044 41188 23662
rect 41468 23492 41524 23502
rect 41132 22978 41188 22988
rect 41356 23380 41412 23390
rect 41356 22372 41412 23324
rect 41468 23378 41524 23436
rect 41468 23326 41470 23378
rect 41522 23326 41524 23378
rect 41468 23314 41524 23326
rect 41356 22306 41412 22316
rect 41132 22260 41188 22270
rect 41132 22146 41188 22204
rect 41132 22094 41134 22146
rect 41186 22094 41188 22146
rect 41132 19796 41188 22094
rect 41244 22258 41300 22270
rect 41244 22206 41246 22258
rect 41298 22206 41300 22258
rect 41244 22036 41300 22206
rect 41244 21970 41300 21980
rect 41468 22036 41524 22046
rect 41356 21140 41412 21150
rect 41244 21028 41300 21038
rect 41244 20802 41300 20972
rect 41244 20750 41246 20802
rect 41298 20750 41300 20802
rect 41244 20738 41300 20750
rect 41132 19730 41188 19740
rect 41244 20578 41300 20590
rect 41244 20526 41246 20578
rect 41298 20526 41300 20578
rect 41132 19010 41188 19022
rect 41132 18958 41134 19010
rect 41186 18958 41188 19010
rect 41132 18004 41188 18958
rect 41132 17668 41188 17948
rect 41244 17892 41300 20526
rect 41244 17826 41300 17836
rect 41244 17668 41300 17678
rect 41132 17666 41300 17668
rect 41132 17614 41246 17666
rect 41298 17614 41300 17666
rect 41132 17612 41300 17614
rect 41244 17444 41300 17612
rect 41244 17378 41300 17388
rect 41356 15148 41412 21084
rect 41468 20802 41524 21980
rect 41580 21812 41636 23884
rect 41916 23874 41972 23884
rect 41804 23716 41860 23726
rect 41804 22482 41860 23660
rect 42028 23716 42084 23726
rect 42028 23622 42084 23660
rect 42140 23714 42196 23726
rect 42140 23662 42142 23714
rect 42194 23662 42196 23714
rect 42140 23268 42196 23662
rect 42252 23716 42308 24444
rect 42476 24434 42532 24444
rect 42364 23940 42420 23950
rect 42364 23846 42420 23884
rect 42252 23660 42420 23716
rect 42140 23202 42196 23212
rect 41804 22430 41806 22482
rect 41858 22430 41860 22482
rect 41804 22418 41860 22430
rect 41916 23042 41972 23054
rect 41916 22990 41918 23042
rect 41970 22990 41972 23042
rect 41692 21812 41748 21822
rect 41580 21810 41748 21812
rect 41580 21758 41694 21810
rect 41746 21758 41748 21810
rect 41580 21756 41748 21758
rect 41692 21746 41748 21756
rect 41916 21812 41972 22990
rect 42252 22820 42308 22830
rect 42028 22708 42084 22718
rect 42028 21812 42084 22652
rect 42140 22594 42196 22606
rect 42140 22542 42142 22594
rect 42194 22542 42196 22594
rect 42140 22482 42196 22542
rect 42140 22430 42142 22482
rect 42194 22430 42196 22482
rect 42140 22418 42196 22430
rect 42140 21812 42196 21822
rect 42028 21810 42196 21812
rect 42028 21758 42142 21810
rect 42194 21758 42196 21810
rect 42028 21756 42196 21758
rect 41916 21746 41972 21756
rect 41916 21588 41972 21598
rect 41916 21586 42084 21588
rect 41916 21534 41918 21586
rect 41970 21534 42084 21586
rect 41916 21532 42084 21534
rect 41916 21522 41972 21532
rect 41468 20750 41470 20802
rect 41522 20750 41524 20802
rect 41468 20738 41524 20750
rect 41804 21474 41860 21486
rect 41804 21422 41806 21474
rect 41858 21422 41860 21474
rect 41468 19906 41524 19918
rect 41468 19854 41470 19906
rect 41522 19854 41524 19906
rect 41468 19796 41524 19854
rect 41468 19730 41524 19740
rect 41580 19012 41636 19022
rect 41580 18918 41636 18956
rect 41804 18676 41860 21422
rect 41692 18620 41860 18676
rect 41916 21364 41972 21374
rect 41916 20132 41972 21308
rect 42028 21028 42084 21532
rect 42028 20962 42084 20972
rect 42028 20132 42084 20142
rect 41916 20130 42084 20132
rect 41916 20078 42030 20130
rect 42082 20078 42084 20130
rect 41916 20076 42084 20078
rect 41580 17108 41636 17118
rect 41468 16884 41524 16894
rect 41468 16790 41524 16828
rect 41020 15038 41022 15090
rect 41074 15038 41076 15090
rect 40012 14130 40068 14140
rect 40348 14084 40404 14588
rect 40796 14532 40852 14542
rect 40796 14438 40852 14476
rect 40684 14420 40740 14430
rect 39452 14028 39844 14084
rect 38780 13804 38948 13860
rect 39340 13860 39396 13870
rect 39452 13860 39508 14028
rect 39340 13858 39508 13860
rect 39340 13806 39342 13858
rect 39394 13806 39508 13858
rect 39340 13804 39508 13806
rect 39564 13858 39620 13870
rect 39564 13806 39566 13858
rect 39618 13806 39620 13858
rect 38668 13748 38724 13758
rect 38780 13748 38836 13804
rect 39340 13794 39396 13804
rect 39564 13748 39620 13806
rect 39676 13860 39732 13870
rect 39676 13766 39732 13804
rect 38668 13746 38836 13748
rect 38668 13694 38670 13746
rect 38722 13694 38836 13746
rect 38668 13692 38836 13694
rect 39452 13692 39620 13748
rect 38668 13682 38724 13692
rect 39116 13634 39172 13646
rect 39116 13582 39118 13634
rect 39170 13582 39172 13634
rect 39116 12852 39172 13582
rect 39452 13412 39508 13692
rect 39452 13346 39508 13356
rect 39676 13524 39732 13534
rect 39116 12786 39172 12796
rect 39228 13300 39284 13310
rect 39228 13074 39284 13244
rect 39228 13022 39230 13074
rect 39282 13022 39284 13074
rect 39116 12628 39172 12638
rect 38780 12180 38836 12190
rect 38780 12086 38836 12124
rect 38556 11778 38612 11788
rect 38892 11732 38948 11742
rect 38780 11508 38836 11518
rect 38892 11508 38948 11676
rect 38780 11506 38948 11508
rect 38780 11454 38782 11506
rect 38834 11454 38948 11506
rect 38780 11452 38948 11454
rect 39116 11506 39172 12572
rect 39228 11618 39284 13022
rect 39452 13076 39508 13086
rect 39452 12982 39508 13020
rect 39340 12964 39396 12974
rect 39340 12402 39396 12908
rect 39340 12350 39342 12402
rect 39394 12350 39396 12402
rect 39340 12338 39396 12350
rect 39676 12402 39732 13468
rect 39788 13076 39844 14028
rect 40236 14028 40404 14084
rect 40460 14306 40516 14318
rect 40460 14254 40462 14306
rect 40514 14254 40516 14306
rect 40236 13972 40292 14028
rect 39900 13748 39956 13758
rect 39900 13654 39956 13692
rect 39788 13010 39844 13020
rect 39788 12740 39844 12750
rect 39788 12738 40068 12740
rect 39788 12686 39790 12738
rect 39842 12686 40068 12738
rect 39788 12684 40068 12686
rect 39788 12674 39844 12684
rect 39676 12350 39678 12402
rect 39730 12350 39732 12402
rect 39676 12338 39732 12350
rect 39228 11566 39230 11618
rect 39282 11566 39284 11618
rect 39228 11554 39284 11566
rect 39788 11618 39844 11630
rect 39788 11566 39790 11618
rect 39842 11566 39844 11618
rect 39116 11454 39118 11506
rect 39170 11454 39172 11506
rect 38780 11442 38836 11452
rect 37548 11230 37550 11282
rect 37602 11230 37604 11282
rect 37548 11218 37604 11230
rect 37884 11282 37940 11294
rect 37884 11230 37886 11282
rect 37938 11230 37940 11282
rect 37436 10782 37438 10834
rect 37490 10782 37492 10834
rect 37436 10770 37492 10782
rect 37660 10722 37716 10734
rect 37660 10670 37662 10722
rect 37714 10670 37716 10722
rect 37660 10612 37716 10670
rect 37324 10556 37716 10612
rect 36316 10334 36318 10386
rect 36370 10334 36372 10386
rect 36316 10322 36372 10334
rect 36540 10498 36596 10510
rect 36540 10446 36542 10498
rect 36594 10446 36596 10498
rect 35868 9650 35924 9660
rect 35980 10052 36036 10062
rect 35084 9436 35252 9492
rect 35420 9602 35476 9614
rect 35420 9550 35422 9602
rect 35474 9550 35476 9602
rect 35420 9492 35476 9550
rect 35084 9380 35140 9436
rect 35420 9426 35476 9436
rect 35868 9492 35924 9502
rect 34636 9202 34692 9212
rect 34972 9324 35140 9380
rect 34972 9154 35028 9324
rect 35196 9268 35252 9278
rect 35196 9156 35252 9212
rect 34972 9102 34974 9154
rect 35026 9102 35028 9154
rect 34636 8372 34692 8382
rect 34636 8278 34692 8316
rect 34972 8258 35028 9102
rect 34972 8206 34974 8258
rect 35026 8206 35028 8258
rect 34972 8194 35028 8206
rect 35084 9154 35252 9156
rect 35084 9102 35198 9154
rect 35250 9102 35252 9154
rect 35084 9100 35252 9102
rect 34636 8146 34692 8158
rect 34636 8094 34638 8146
rect 34690 8094 34692 8146
rect 34636 7924 34692 8094
rect 35084 8146 35140 9100
rect 35196 9090 35252 9100
rect 35532 9156 35588 9166
rect 35532 9062 35588 9100
rect 35868 9156 35924 9436
rect 35980 9266 36036 9996
rect 36540 9828 36596 10446
rect 36540 9762 36596 9772
rect 36092 9716 36148 9726
rect 36092 9622 36148 9660
rect 36316 9714 36372 9726
rect 36316 9662 36318 9714
rect 36370 9662 36372 9714
rect 36316 9492 36372 9662
rect 36652 9604 36708 10556
rect 36876 10386 36932 10398
rect 36876 10334 36878 10386
rect 36930 10334 36932 10386
rect 36764 9828 36820 9838
rect 36764 9734 36820 9772
rect 36876 9716 36932 10334
rect 36876 9660 37268 9716
rect 36652 9548 36932 9604
rect 35980 9214 35982 9266
rect 36034 9214 36036 9266
rect 35980 9202 36036 9214
rect 36092 9436 36372 9492
rect 35868 9090 35924 9100
rect 35420 8930 35476 8942
rect 35420 8878 35422 8930
rect 35474 8878 35476 8930
rect 35420 8820 35476 8878
rect 35420 8764 35588 8820
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35532 8372 35588 8764
rect 35532 8306 35588 8316
rect 36092 8484 36148 9436
rect 36204 9268 36260 9278
rect 36204 9266 36596 9268
rect 36204 9214 36206 9266
rect 36258 9214 36596 9266
rect 36204 9212 36596 9214
rect 36204 9202 36260 9212
rect 36316 9044 36372 9054
rect 36316 8950 36372 8988
rect 35084 8094 35086 8146
rect 35138 8094 35140 8146
rect 35084 8036 35140 8094
rect 35084 7970 35140 7980
rect 35196 8148 35252 8158
rect 34636 7858 34692 7868
rect 35196 7476 35252 8092
rect 35980 8034 36036 8046
rect 35980 7982 35982 8034
rect 36034 7982 36036 8034
rect 34524 7410 34580 7420
rect 34972 7474 35252 7476
rect 34972 7422 35198 7474
rect 35250 7422 35252 7474
rect 34972 7420 35252 7422
rect 34972 6916 35028 7420
rect 35196 7410 35252 7420
rect 35644 7474 35700 7486
rect 35644 7422 35646 7474
rect 35698 7422 35700 7474
rect 35084 7252 35140 7262
rect 35084 7158 35140 7196
rect 35420 7252 35476 7262
rect 35420 7250 35588 7252
rect 35420 7198 35422 7250
rect 35474 7198 35588 7250
rect 35420 7196 35588 7198
rect 35420 7186 35476 7196
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 34972 6860 35364 6916
rect 35308 6804 35364 6860
rect 33740 6692 33796 6702
rect 33740 6468 33796 6636
rect 34636 6692 34692 6702
rect 34636 6598 34692 6636
rect 35308 6690 35364 6748
rect 35308 6638 35310 6690
rect 35362 6638 35364 6690
rect 35308 6626 35364 6638
rect 33852 6468 33908 6478
rect 33740 6466 33908 6468
rect 33740 6414 33854 6466
rect 33906 6414 33908 6466
rect 33740 6412 33908 6414
rect 33740 6132 33796 6412
rect 33852 6402 33908 6412
rect 35084 6468 35140 6478
rect 35084 6374 35140 6412
rect 35196 6466 35252 6478
rect 35196 6414 35198 6466
rect 35250 6414 35252 6466
rect 33628 6020 33684 6030
rect 33628 5926 33684 5964
rect 33740 5348 33796 6076
rect 33964 5908 34020 5918
rect 33964 5814 34020 5852
rect 35196 5908 35252 6414
rect 35532 6468 35588 7196
rect 35644 6692 35700 7422
rect 35756 6692 35812 6702
rect 35644 6690 35812 6692
rect 35644 6638 35758 6690
rect 35810 6638 35812 6690
rect 35644 6636 35812 6638
rect 35532 6402 35588 6412
rect 35196 5842 35252 5852
rect 35756 5908 35812 6636
rect 35756 5814 35812 5852
rect 35980 6468 36036 7982
rect 36092 7588 36148 8428
rect 36540 8482 36596 9212
rect 36764 8932 36820 8942
rect 36764 8838 36820 8876
rect 36540 8430 36542 8482
rect 36594 8430 36596 8482
rect 36428 8372 36484 8382
rect 36428 8278 36484 8316
rect 36540 8260 36596 8430
rect 36540 8194 36596 8204
rect 36204 7588 36260 7598
rect 36092 7586 36260 7588
rect 36092 7534 36206 7586
rect 36258 7534 36260 7586
rect 36092 7532 36260 7534
rect 36204 7522 36260 7532
rect 36540 7588 36596 7598
rect 36540 7494 36596 7532
rect 36204 6804 36260 6814
rect 36204 6578 36260 6748
rect 36540 6804 36596 6814
rect 36204 6526 36206 6578
rect 36258 6526 36260 6578
rect 36204 6514 36260 6526
rect 36316 6692 36372 6702
rect 36540 6692 36596 6748
rect 36372 6690 36596 6692
rect 36372 6638 36542 6690
rect 36594 6638 36596 6690
rect 36372 6636 36596 6638
rect 34188 5796 34244 5806
rect 34188 5702 34244 5740
rect 34636 5794 34692 5806
rect 34636 5742 34638 5794
rect 34690 5742 34692 5794
rect 33740 5234 33796 5292
rect 34636 5572 34692 5742
rect 35308 5796 35364 5806
rect 35308 5702 35364 5740
rect 35980 5796 36036 6412
rect 36204 5908 36260 5918
rect 36316 5908 36372 6636
rect 36540 6626 36596 6636
rect 36204 5906 36372 5908
rect 36204 5854 36206 5906
rect 36258 5854 36372 5906
rect 36204 5852 36372 5854
rect 36204 5842 36260 5852
rect 35980 5702 36036 5740
rect 36652 5796 36708 5806
rect 36652 5702 36708 5740
rect 33740 5182 33742 5234
rect 33794 5182 33796 5234
rect 33740 5170 33796 5182
rect 34524 5236 34580 5246
rect 33516 4946 33572 4956
rect 33516 4676 33572 4686
rect 33516 4562 33572 4620
rect 33516 4510 33518 4562
rect 33570 4510 33572 4562
rect 33516 4498 33572 4510
rect 33852 4452 33908 4462
rect 33292 1474 33348 1484
rect 33628 3668 33684 3678
rect 33628 800 33684 3612
rect 33852 3554 33908 4396
rect 34524 4338 34580 5180
rect 34636 5010 34692 5516
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 36540 5236 36596 5246
rect 36540 5142 36596 5180
rect 34636 4958 34638 5010
rect 34690 4958 34692 5010
rect 34636 4946 34692 4958
rect 34524 4286 34526 4338
rect 34578 4286 34580 4338
rect 34524 4274 34580 4286
rect 34972 4340 35028 4350
rect 34972 4246 35028 4284
rect 35644 4340 35700 4350
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 34524 3668 34580 3678
rect 34524 3574 34580 3612
rect 35644 3666 35700 4284
rect 35644 3614 35646 3666
rect 35698 3614 35700 3666
rect 35644 3602 35700 3614
rect 36876 4340 36932 9548
rect 37212 9266 37268 9660
rect 37212 9214 37214 9266
rect 37266 9214 37268 9266
rect 36988 8372 37044 8382
rect 36988 7812 37044 8316
rect 37212 8372 37268 9214
rect 37212 8306 37268 8316
rect 37548 8260 37604 8270
rect 37548 8166 37604 8204
rect 36988 7698 37044 7756
rect 36988 7646 36990 7698
rect 37042 7646 37044 7698
rect 36988 7634 37044 7646
rect 37660 7588 37716 10556
rect 37772 10610 37828 10622
rect 37772 10558 37774 10610
rect 37826 10558 37828 10610
rect 37772 9940 37828 10558
rect 37884 10612 37940 11230
rect 38668 10724 38724 10734
rect 38444 10612 38500 10622
rect 37884 10610 38500 10612
rect 37884 10558 38446 10610
rect 38498 10558 38500 10610
rect 37884 10556 38500 10558
rect 37884 9940 37940 9950
rect 37772 9938 37940 9940
rect 37772 9886 37886 9938
rect 37938 9886 37940 9938
rect 37772 9884 37940 9886
rect 37884 9874 37940 9884
rect 38332 9938 38388 9950
rect 38332 9886 38334 9938
rect 38386 9886 38388 9938
rect 38332 9268 38388 9886
rect 38444 9492 38500 10556
rect 38668 10276 38724 10668
rect 38668 10210 38724 10220
rect 38556 9828 38612 9838
rect 38556 9734 38612 9772
rect 39116 9828 39172 11454
rect 39788 11506 39844 11566
rect 39788 11454 39790 11506
rect 39842 11454 39844 11506
rect 39788 11442 39844 11454
rect 39340 10836 39396 10846
rect 40012 10836 40068 12684
rect 40236 12402 40292 13916
rect 40348 13860 40404 13870
rect 40348 13766 40404 13804
rect 40460 13748 40516 14254
rect 40572 13972 40628 13982
rect 40684 13972 40740 14364
rect 40572 13970 40740 13972
rect 40572 13918 40574 13970
rect 40626 13918 40740 13970
rect 40572 13916 40740 13918
rect 40572 13906 40628 13916
rect 40684 13748 40740 13758
rect 41020 13748 41076 15038
rect 40460 13746 40852 13748
rect 40460 13694 40686 13746
rect 40738 13694 40852 13746
rect 40460 13692 40852 13694
rect 40684 13682 40740 13692
rect 40684 13524 40740 13534
rect 40236 12350 40238 12402
rect 40290 12350 40292 12402
rect 40236 12338 40292 12350
rect 40348 13412 40404 13422
rect 40348 12740 40404 13356
rect 40348 12180 40404 12684
rect 40124 12124 40404 12180
rect 40572 13076 40628 13086
rect 40572 12292 40628 13020
rect 40124 11506 40180 12124
rect 40124 11454 40126 11506
rect 40178 11454 40180 11506
rect 40124 11442 40180 11454
rect 40572 11506 40628 12236
rect 40684 12738 40740 13468
rect 40684 12686 40686 12738
rect 40738 12686 40740 12738
rect 40684 11956 40740 12686
rect 40684 11890 40740 11900
rect 40796 13524 40852 13692
rect 41020 13682 41076 13692
rect 41132 15092 41412 15148
rect 41468 15314 41524 15326
rect 41468 15262 41470 15314
rect 41522 15262 41524 15314
rect 41468 15092 41524 15262
rect 41132 13524 41188 15092
rect 41468 15026 41524 15036
rect 41580 14980 41636 17052
rect 41580 14914 41636 14924
rect 41692 14756 41748 18620
rect 41804 18452 41860 18462
rect 41804 16884 41860 18396
rect 41916 18450 41972 20076
rect 42028 20066 42084 20076
rect 42028 19348 42084 19358
rect 42028 19254 42084 19292
rect 42140 18788 42196 21756
rect 42140 18722 42196 18732
rect 42252 18676 42308 22764
rect 42364 21700 42420 23660
rect 42476 23154 42532 23166
rect 42476 23102 42478 23154
rect 42530 23102 42532 23154
rect 42476 23044 42532 23102
rect 42476 22978 42532 22988
rect 42588 22596 42644 24444
rect 42700 24610 42756 24622
rect 42700 24558 42702 24610
rect 42754 24558 42756 24610
rect 42700 23938 42756 24558
rect 42700 23886 42702 23938
rect 42754 23886 42756 23938
rect 42700 23874 42756 23886
rect 42924 23716 42980 24668
rect 42812 23266 42868 23278
rect 42812 23214 42814 23266
rect 42866 23214 42868 23266
rect 42588 22530 42644 22540
rect 42700 23156 42756 23166
rect 42588 22372 42644 22382
rect 42588 22278 42644 22316
rect 42700 21810 42756 23100
rect 42812 22820 42868 23214
rect 42812 22754 42868 22764
rect 42700 21758 42702 21810
rect 42754 21758 42756 21810
rect 42700 21746 42756 21758
rect 42364 21634 42420 21644
rect 42476 21476 42532 21486
rect 42364 20804 42420 20814
rect 42476 20804 42532 21420
rect 42588 20804 42644 20814
rect 42924 20804 42980 23660
rect 43036 24498 43092 24510
rect 43036 24446 43038 24498
rect 43090 24446 43092 24498
rect 43036 23044 43092 24446
rect 43036 22978 43092 22988
rect 43148 22372 43204 25340
rect 43260 25394 43316 25452
rect 43260 25342 43262 25394
rect 43314 25342 43316 25394
rect 43260 25330 43316 25342
rect 43372 25396 43428 25406
rect 43148 22306 43204 22316
rect 43260 23044 43316 23054
rect 43372 23044 43428 25340
rect 43260 23042 43428 23044
rect 43260 22990 43262 23042
rect 43314 22990 43428 23042
rect 43260 22988 43428 22990
rect 43260 22594 43316 22988
rect 43260 22542 43262 22594
rect 43314 22542 43316 22594
rect 43036 22148 43092 22158
rect 43260 22148 43316 22542
rect 43036 22054 43092 22092
rect 43148 22092 43316 22148
rect 43148 21476 43204 22092
rect 43484 21924 43540 28476
rect 43596 27636 43652 27646
rect 43596 27412 43652 27580
rect 43596 27186 43652 27356
rect 43708 27298 43764 28588
rect 43820 28420 43876 28430
rect 43876 28364 44100 28420
rect 43820 28326 43876 28364
rect 44044 28082 44100 28364
rect 44044 28030 44046 28082
rect 44098 28030 44100 28082
rect 44044 28018 44100 28030
rect 43708 27246 43710 27298
rect 43762 27246 43764 27298
rect 43708 27234 43764 27246
rect 43820 27858 43876 27870
rect 43820 27806 43822 27858
rect 43874 27806 43876 27858
rect 43820 27748 43876 27806
rect 43596 27134 43598 27186
rect 43650 27134 43652 27186
rect 43596 27122 43652 27134
rect 43820 27188 43876 27692
rect 43820 27122 43876 27132
rect 43932 27746 43988 27758
rect 43932 27694 43934 27746
rect 43986 27694 43988 27746
rect 43932 26402 43988 27694
rect 44156 27412 44212 29372
rect 44716 29204 44772 29214
rect 44716 29202 44884 29204
rect 44716 29150 44718 29202
rect 44770 29150 44884 29202
rect 44716 29148 44884 29150
rect 44716 29138 44772 29148
rect 44716 28530 44772 28542
rect 44716 28478 44718 28530
rect 44770 28478 44772 28530
rect 44380 28418 44436 28430
rect 44380 28366 44382 28418
rect 44434 28366 44436 28418
rect 44156 27356 44324 27412
rect 44044 27300 44100 27310
rect 44044 27298 44212 27300
rect 44044 27246 44046 27298
rect 44098 27246 44212 27298
rect 44044 27244 44212 27246
rect 44044 27234 44100 27244
rect 44156 27186 44212 27244
rect 44156 27134 44158 27186
rect 44210 27134 44212 27186
rect 44156 27122 44212 27134
rect 43932 26350 43934 26402
rect 43986 26350 43988 26402
rect 43932 26338 43988 26350
rect 44156 26852 44212 26862
rect 43820 26292 43876 26302
rect 43708 25620 43764 25630
rect 43708 24724 43764 25564
rect 43820 25506 43876 26236
rect 43820 25454 43822 25506
rect 43874 25454 43876 25506
rect 43820 25442 43876 25454
rect 44156 25508 44212 26796
rect 44268 26290 44324 27356
rect 44380 26740 44436 28366
rect 44492 27972 44548 27982
rect 44492 27858 44548 27916
rect 44716 27972 44772 28478
rect 44716 27906 44772 27916
rect 44492 27806 44494 27858
rect 44546 27806 44548 27858
rect 44492 27524 44548 27806
rect 44492 27458 44548 27468
rect 44492 26964 44548 26974
rect 44492 26870 44548 26908
rect 44828 26908 44884 29148
rect 45276 26964 45332 29932
rect 45388 29922 45444 29932
rect 45948 29876 46004 30942
rect 46060 30996 46116 31006
rect 46060 30210 46116 30940
rect 46060 30158 46062 30210
rect 46114 30158 46116 30210
rect 46060 30146 46116 30158
rect 46172 30436 46228 30446
rect 45948 29820 46116 29876
rect 45948 29652 46004 29662
rect 45948 29540 46004 29596
rect 45724 29538 46004 29540
rect 45724 29486 45950 29538
rect 46002 29486 46004 29538
rect 45724 29484 46004 29486
rect 45724 29092 45780 29484
rect 45948 29474 46004 29484
rect 46060 29426 46116 29820
rect 46060 29374 46062 29426
rect 46114 29374 46116 29426
rect 45612 29036 45780 29092
rect 45836 29316 45892 29326
rect 45612 28530 45668 29036
rect 45612 28478 45614 28530
rect 45666 28478 45668 28530
rect 45612 28466 45668 28478
rect 45724 28532 45780 28542
rect 45836 28532 45892 29260
rect 45948 29314 46004 29326
rect 45948 29262 45950 29314
rect 46002 29262 46004 29314
rect 45948 28980 46004 29262
rect 46060 29316 46116 29374
rect 46060 29250 46116 29260
rect 45948 28914 46004 28924
rect 46172 28754 46228 30380
rect 46284 29988 46340 33628
rect 46620 33236 46676 33246
rect 46620 32786 46676 33180
rect 46732 32900 46788 55412
rect 47180 55188 47236 55198
rect 47180 55094 47236 55132
rect 47516 55186 47572 56028
rect 51772 55972 51828 59200
rect 55804 57204 55860 57214
rect 55804 56194 55860 57148
rect 55804 56142 55806 56194
rect 55858 56142 55860 56194
rect 55804 56130 55860 56142
rect 52780 56084 52836 56094
rect 52780 55990 52836 56028
rect 54684 56082 54740 56094
rect 54684 56030 54686 56082
rect 54738 56030 54740 56082
rect 51772 55906 51828 55916
rect 53452 55972 53508 55982
rect 53452 55878 53508 55916
rect 47516 55134 47518 55186
rect 47570 55134 47572 55186
rect 47516 55122 47572 55134
rect 53900 55522 53956 55534
rect 53900 55470 53902 55522
rect 53954 55470 53956 55522
rect 53900 55074 53956 55470
rect 54684 55522 54740 56030
rect 54684 55470 54686 55522
rect 54738 55470 54740 55522
rect 54684 55458 54740 55470
rect 56028 55412 56084 55422
rect 56028 55318 56084 55356
rect 57148 55412 57204 59200
rect 57148 55346 57204 55356
rect 54908 55300 54964 55310
rect 54348 55298 54964 55300
rect 54348 55246 54910 55298
rect 54962 55246 54964 55298
rect 54348 55244 54964 55246
rect 54348 55076 54404 55244
rect 54908 55234 54964 55244
rect 53900 55022 53902 55074
rect 53954 55022 53956 55074
rect 47068 54964 47124 54974
rect 46844 40404 46900 40414
rect 46844 40310 46900 40348
rect 47068 34916 47124 54908
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 49532 53844 49588 53854
rect 48748 52164 48804 52174
rect 48748 51602 48804 52108
rect 48748 51550 48750 51602
rect 48802 51550 48804 51602
rect 48748 51538 48804 51550
rect 48412 51378 48468 51390
rect 48412 51326 48414 51378
rect 48466 51326 48468 51378
rect 47852 51268 47908 51278
rect 48412 51268 48468 51326
rect 47852 51266 48468 51268
rect 47852 51214 47854 51266
rect 47906 51214 48468 51266
rect 47852 51212 48468 51214
rect 47404 48916 47460 48926
rect 47404 48822 47460 48860
rect 47852 40516 47908 51212
rect 47852 40450 47908 40460
rect 47516 40290 47572 40302
rect 47516 40238 47518 40290
rect 47570 40238 47572 40290
rect 47516 39618 47572 40238
rect 47516 39566 47518 39618
rect 47570 39566 47572 39618
rect 47516 39554 47572 39566
rect 47852 39394 47908 39406
rect 47852 39342 47854 39394
rect 47906 39342 47908 39394
rect 47852 35924 47908 39342
rect 47852 35858 47908 35868
rect 47068 34850 47124 34860
rect 49532 34580 49588 53788
rect 53900 53844 53956 55022
rect 53900 53778 53956 53788
rect 54236 55074 54404 55076
rect 54236 55022 54350 55074
rect 54402 55022 54404 55074
rect 54236 55020 54404 55022
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 52892 52836 52948 52846
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 52780 35812 52836 35822
rect 49532 34514 49588 34524
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 52332 33684 52388 33694
rect 46732 32834 46788 32844
rect 47516 33236 47572 33246
rect 46620 32734 46622 32786
rect 46674 32734 46676 32786
rect 46620 32722 46676 32734
rect 47516 32564 47572 33180
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 51660 32676 51716 32686
rect 47516 32432 47572 32508
rect 48076 32562 48132 32574
rect 48076 32510 48078 32562
rect 48130 32510 48132 32562
rect 48076 32452 48132 32510
rect 48076 32386 48132 32396
rect 48188 32450 48244 32462
rect 48188 32398 48190 32450
rect 48242 32398 48244 32450
rect 47628 31780 47684 31790
rect 48188 31780 48244 32398
rect 51100 32452 51156 32462
rect 51100 32358 51156 32396
rect 47628 31778 48244 31780
rect 47628 31726 47630 31778
rect 47682 31726 48190 31778
rect 48242 31726 48244 31778
rect 47628 31724 48244 31726
rect 47628 31714 47684 31724
rect 48188 31714 48244 31724
rect 51548 31780 51604 31790
rect 51548 31686 51604 31724
rect 46508 31668 46564 31678
rect 46284 29894 46340 29932
rect 46396 31666 46564 31668
rect 46396 31614 46510 31666
rect 46562 31614 46564 31666
rect 46396 31612 46564 31614
rect 46396 29652 46452 31612
rect 46508 31602 46564 31612
rect 47292 31556 47348 31566
rect 47180 31554 47348 31556
rect 47180 31502 47294 31554
rect 47346 31502 47348 31554
rect 47180 31500 47348 31502
rect 46508 30996 46564 31006
rect 46564 30940 46676 30996
rect 46508 30902 46564 30940
rect 46620 30212 46676 30940
rect 46844 30884 46900 30894
rect 46844 30790 46900 30828
rect 47180 30884 47236 31500
rect 47292 31490 47348 31500
rect 47516 31556 47572 31566
rect 47516 31462 47572 31500
rect 47852 31556 47908 31566
rect 47852 31218 47908 31500
rect 47852 31166 47854 31218
rect 47906 31166 47908 31218
rect 47852 31154 47908 31166
rect 48524 31554 48580 31566
rect 48524 31502 48526 31554
rect 48578 31502 48580 31554
rect 48188 31108 48244 31118
rect 48076 31106 48244 31108
rect 48076 31054 48190 31106
rect 48242 31054 48244 31106
rect 48076 31052 48244 31054
rect 48076 30996 48132 31052
rect 48188 31042 48244 31052
rect 47180 30818 47236 30828
rect 47292 30882 47348 30894
rect 47292 30830 47294 30882
rect 47346 30830 47348 30882
rect 47292 30212 47348 30830
rect 46620 30146 46676 30156
rect 47180 30156 47348 30212
rect 46172 28702 46174 28754
rect 46226 28702 46228 28754
rect 46172 28644 46228 28702
rect 46172 28578 46228 28588
rect 46284 29596 46452 29652
rect 46508 30098 46564 30110
rect 46508 30046 46510 30098
rect 46562 30046 46564 30098
rect 46508 29652 46564 30046
rect 45724 28530 45892 28532
rect 45724 28478 45726 28530
rect 45778 28478 45892 28530
rect 45724 28476 45892 28478
rect 44828 26852 44996 26908
rect 45276 26898 45332 26908
rect 45388 28418 45444 28430
rect 45388 28366 45390 28418
rect 45442 28366 45444 28418
rect 44380 26684 44660 26740
rect 44268 26238 44270 26290
rect 44322 26238 44324 26290
rect 44268 26226 44324 26238
rect 44268 26068 44324 26078
rect 44268 25974 44324 26012
rect 44156 25376 44212 25452
rect 44492 25394 44548 25406
rect 44492 25342 44494 25394
rect 44546 25342 44548 25394
rect 44044 25282 44100 25294
rect 44044 25230 44046 25282
rect 44098 25230 44100 25282
rect 44044 25172 44100 25230
rect 44044 25106 44100 25116
rect 43820 24948 43876 24958
rect 43820 24946 44324 24948
rect 43820 24894 43822 24946
rect 43874 24894 44324 24946
rect 43820 24892 44324 24894
rect 43820 24882 43876 24892
rect 43708 24668 43876 24724
rect 43708 23940 43764 23950
rect 43708 23846 43764 23884
rect 43820 23826 43876 24668
rect 43932 24722 43988 24734
rect 43932 24670 43934 24722
rect 43986 24670 43988 24722
rect 43932 24612 43988 24670
rect 44156 24722 44212 24734
rect 44156 24670 44158 24722
rect 44210 24670 44212 24722
rect 43932 24546 43988 24556
rect 44044 24610 44100 24622
rect 44044 24558 44046 24610
rect 44098 24558 44100 24610
rect 44044 24164 44100 24558
rect 44044 24098 44100 24108
rect 44156 24276 44212 24670
rect 43820 23774 43822 23826
rect 43874 23774 43876 23826
rect 43820 23762 43876 23774
rect 43932 23826 43988 23838
rect 43932 23774 43934 23826
rect 43986 23774 43988 23826
rect 43596 23714 43652 23726
rect 43596 23662 43598 23714
rect 43650 23662 43652 23714
rect 43596 23156 43652 23662
rect 43596 23090 43652 23100
rect 43708 23604 43764 23614
rect 43708 23042 43764 23548
rect 43932 23604 43988 23774
rect 43932 23538 43988 23548
rect 44044 23826 44100 23838
rect 44044 23774 44046 23826
rect 44098 23774 44100 23826
rect 43708 22990 43710 23042
rect 43762 22990 43764 23042
rect 43708 22708 43764 22990
rect 43708 22642 43764 22652
rect 43820 23380 43876 23390
rect 43596 22596 43652 22606
rect 43596 22482 43652 22540
rect 43596 22430 43598 22482
rect 43650 22430 43652 22482
rect 43596 22418 43652 22430
rect 43148 21410 43204 21420
rect 43260 21868 43540 21924
rect 43596 22260 43652 22270
rect 42476 20802 42644 20804
rect 42476 20750 42590 20802
rect 42642 20750 42644 20802
rect 42476 20748 42644 20750
rect 42364 20710 42420 20748
rect 42588 20738 42644 20748
rect 42700 20748 42980 20804
rect 43036 21364 43092 21374
rect 42476 20578 42532 20590
rect 42700 20580 42756 20748
rect 42476 20526 42478 20578
rect 42530 20526 42532 20578
rect 42476 20356 42532 20526
rect 42476 20290 42532 20300
rect 42588 20524 42756 20580
rect 42812 20578 42868 20590
rect 42812 20526 42814 20578
rect 42866 20526 42868 20578
rect 42364 20020 42420 20030
rect 42364 20018 42532 20020
rect 42364 19966 42366 20018
rect 42418 19966 42532 20018
rect 42364 19964 42532 19966
rect 42364 19954 42420 19964
rect 42252 18610 42308 18620
rect 42364 19572 42420 19582
rect 42140 18564 42196 18574
rect 41916 18398 41918 18450
rect 41970 18398 41972 18450
rect 41916 18386 41972 18398
rect 42028 18450 42084 18462
rect 42028 18398 42030 18450
rect 42082 18398 42084 18450
rect 41916 18228 41972 18238
rect 41916 17554 41972 18172
rect 41916 17502 41918 17554
rect 41970 17502 41972 17554
rect 41916 17108 41972 17502
rect 42028 17108 42084 18398
rect 42140 17666 42196 18508
rect 42364 18562 42420 19516
rect 42364 18510 42366 18562
rect 42418 18510 42420 18562
rect 42364 18498 42420 18510
rect 42252 18340 42308 18350
rect 42252 18246 42308 18284
rect 42476 18228 42532 19964
rect 42476 18162 42532 18172
rect 42588 18004 42644 20524
rect 42812 19348 42868 20526
rect 43036 20468 43092 21308
rect 42924 20244 42980 20254
rect 43036 20244 43092 20412
rect 42924 20242 43092 20244
rect 42924 20190 42926 20242
rect 42978 20190 43092 20242
rect 42924 20188 43092 20190
rect 42924 20178 42980 20188
rect 43148 20020 43204 20030
rect 42812 19282 42868 19292
rect 43036 20018 43204 20020
rect 43036 19966 43150 20018
rect 43202 19966 43204 20018
rect 43036 19964 43204 19966
rect 42812 19012 42868 19022
rect 43036 19012 43092 19964
rect 43148 19954 43204 19964
rect 43148 19236 43204 19246
rect 43260 19236 43316 21868
rect 43596 21812 43652 22204
rect 43820 21812 43876 23324
rect 44044 22372 44100 23774
rect 44156 23268 44212 24220
rect 44268 23492 44324 24892
rect 44380 24724 44436 24734
rect 44380 24630 44436 24668
rect 44492 23828 44548 25342
rect 44492 23762 44548 23772
rect 44604 24612 44660 26684
rect 44828 26516 44884 26526
rect 44828 26290 44884 26460
rect 44828 26238 44830 26290
rect 44882 26238 44884 26290
rect 44828 26226 44884 26238
rect 44268 23426 44324 23436
rect 44380 23604 44436 23614
rect 44156 23212 44324 23268
rect 43484 21756 43652 21812
rect 43708 21756 43876 21812
rect 43932 22316 44100 22372
rect 44156 23042 44212 23054
rect 44156 22990 44158 23042
rect 44210 22990 44212 23042
rect 44156 22932 44212 22990
rect 44156 22372 44212 22876
rect 43932 22148 43988 22316
rect 44156 22306 44212 22316
rect 43484 21698 43540 21756
rect 43708 21700 43764 21756
rect 43484 21646 43486 21698
rect 43538 21646 43540 21698
rect 43484 21634 43540 21646
rect 43596 21644 43764 21700
rect 43596 21642 43652 21644
rect 43596 21590 43598 21642
rect 43650 21590 43652 21642
rect 43596 21578 43652 21590
rect 43484 21362 43540 21374
rect 43484 21310 43486 21362
rect 43538 21310 43540 21362
rect 43484 20804 43540 21310
rect 43484 20738 43540 20748
rect 43820 20804 43876 20814
rect 43820 20710 43876 20748
rect 43708 20692 43764 20702
rect 43708 20356 43764 20636
rect 43708 20290 43764 20300
rect 43932 20242 43988 22092
rect 44044 22146 44100 22158
rect 44044 22094 44046 22146
rect 44098 22094 44100 22146
rect 44044 21812 44100 22094
rect 44044 21746 44100 21756
rect 44156 22036 44212 22046
rect 44044 21588 44100 21598
rect 44156 21588 44212 21980
rect 44044 21586 44212 21588
rect 44044 21534 44046 21586
rect 44098 21534 44212 21586
rect 44044 21532 44212 21534
rect 44044 21522 44100 21532
rect 44044 20692 44100 20702
rect 44044 20598 44100 20636
rect 44156 20580 44212 20590
rect 44156 20486 44212 20524
rect 44268 20578 44324 23212
rect 44380 22370 44436 23548
rect 44604 23380 44660 24556
rect 44604 23314 44660 23324
rect 44716 25508 44772 25518
rect 44716 23378 44772 25452
rect 44716 23326 44718 23378
rect 44770 23326 44772 23378
rect 44716 23314 44772 23326
rect 44380 22318 44382 22370
rect 44434 22318 44436 22370
rect 44380 22306 44436 22318
rect 44492 22596 44548 22606
rect 44492 22036 44548 22540
rect 44716 22036 44772 22046
rect 44548 21980 44660 22036
rect 44492 21970 44548 21980
rect 44268 20526 44270 20578
rect 44322 20526 44324 20578
rect 43932 20190 43934 20242
rect 43986 20190 43988 20242
rect 43932 20178 43988 20190
rect 44156 20356 44212 20366
rect 44156 20242 44212 20300
rect 44156 20190 44158 20242
rect 44210 20190 44212 20242
rect 44156 20178 44212 20190
rect 43820 19908 43876 19918
rect 43820 19814 43876 19852
rect 44268 19908 44324 20526
rect 44380 21812 44436 21822
rect 44380 20356 44436 21756
rect 44492 21588 44548 21598
rect 44492 21474 44548 21532
rect 44492 21422 44494 21474
rect 44546 21422 44548 21474
rect 44492 20916 44548 21422
rect 44492 20850 44548 20860
rect 44380 20290 44436 20300
rect 44268 19842 44324 19852
rect 44380 20018 44436 20030
rect 44380 19966 44382 20018
rect 44434 19966 44436 20018
rect 44268 19460 44324 19470
rect 44380 19460 44436 19966
rect 44268 19458 44436 19460
rect 44268 19406 44270 19458
rect 44322 19406 44436 19458
rect 44268 19404 44436 19406
rect 44268 19394 44324 19404
rect 43148 19234 43260 19236
rect 43148 19182 43150 19234
rect 43202 19182 43260 19234
rect 43148 19180 43260 19182
rect 43148 19170 43204 19180
rect 43260 19104 43316 19180
rect 44380 19236 44436 19246
rect 43596 19124 43652 19134
rect 42812 19010 43092 19012
rect 42812 18958 42814 19010
rect 42866 18958 43092 19010
rect 42812 18956 43092 18958
rect 43596 19010 43652 19068
rect 43596 18958 43598 19010
rect 43650 18958 43652 19010
rect 42812 18946 42868 18956
rect 42812 18788 42868 18798
rect 42812 18674 42868 18732
rect 42812 18622 42814 18674
rect 42866 18622 42868 18674
rect 42364 17948 42644 18004
rect 42700 18340 42756 18350
rect 42140 17614 42142 17666
rect 42194 17614 42196 17666
rect 42140 17602 42196 17614
rect 42252 17668 42308 17678
rect 42028 17052 42196 17108
rect 41916 17042 41972 17052
rect 42028 16884 42084 16894
rect 41804 16882 42084 16884
rect 41804 16830 42030 16882
rect 42082 16830 42084 16882
rect 41804 16828 42084 16830
rect 41692 14690 41748 14700
rect 41804 16210 41860 16222
rect 41804 16158 41806 16210
rect 41858 16158 41860 16210
rect 41692 14532 41748 14542
rect 41692 14438 41748 14476
rect 41804 14530 41860 16158
rect 41916 16100 41972 16110
rect 41916 15986 41972 16044
rect 41916 15934 41918 15986
rect 41970 15934 41972 15986
rect 41916 15922 41972 15934
rect 42028 15652 42084 16828
rect 42140 16212 42196 17052
rect 42252 17106 42308 17612
rect 42252 17054 42254 17106
rect 42306 17054 42308 17106
rect 42252 17042 42308 17054
rect 42140 16146 42196 16156
rect 42140 15988 42196 15998
rect 42364 15988 42420 17948
rect 42700 17666 42756 18284
rect 42700 17614 42702 17666
rect 42754 17614 42756 17666
rect 42700 17602 42756 17614
rect 42812 17668 42868 18622
rect 42812 17602 42868 17612
rect 42588 17554 42644 17566
rect 42588 17502 42590 17554
rect 42642 17502 42644 17554
rect 42588 17220 42644 17502
rect 42588 16996 42644 17164
rect 42588 16930 42644 16940
rect 42924 17332 42980 18956
rect 43596 18788 43652 18958
rect 44268 19010 44324 19022
rect 44268 18958 44270 19010
rect 44322 18958 44324 19010
rect 43596 18722 43652 18732
rect 44156 18900 44212 18910
rect 42924 16994 42980 17276
rect 42924 16942 42926 16994
rect 42978 16942 42980 16994
rect 42924 16930 42980 16942
rect 43148 18676 43204 18686
rect 42700 16884 42756 16894
rect 42700 16660 42756 16828
rect 43148 16884 43204 18620
rect 43932 18676 43988 18714
rect 43932 18610 43988 18620
rect 44156 18674 44212 18844
rect 44156 18622 44158 18674
rect 44210 18622 44212 18674
rect 44156 18610 44212 18622
rect 44044 18564 44100 18574
rect 44044 18470 44100 18508
rect 43820 18452 43876 18462
rect 43820 18358 43876 18396
rect 44268 18452 44324 18958
rect 44380 18788 44436 19180
rect 44604 19012 44660 21980
rect 44716 21252 44772 21980
rect 44716 21196 44884 21252
rect 44716 21028 44772 21038
rect 44716 20914 44772 20972
rect 44716 20862 44718 20914
rect 44770 20862 44772 20914
rect 44716 20850 44772 20862
rect 44828 19572 44884 21196
rect 44828 19506 44884 19516
rect 44940 19236 44996 26852
rect 45276 24276 45332 24286
rect 45052 23044 45108 23054
rect 45052 22260 45108 22988
rect 45052 22194 45108 22204
rect 45164 21698 45220 21710
rect 45164 21646 45166 21698
rect 45218 21646 45220 21698
rect 45052 21588 45108 21598
rect 45052 21494 45108 21532
rect 45164 21476 45220 21646
rect 45164 21410 45220 21420
rect 44940 19170 44996 19180
rect 45052 19572 45108 19582
rect 44604 18956 44996 19012
rect 44380 18732 44660 18788
rect 44380 18564 44436 18574
rect 44380 18470 44436 18508
rect 44268 18386 44324 18396
rect 44492 18452 44548 18462
rect 43708 18228 43764 18238
rect 43372 17220 43428 17230
rect 43148 16882 43316 16884
rect 43148 16830 43150 16882
rect 43202 16830 43316 16882
rect 43148 16828 43316 16830
rect 43148 16818 43204 16828
rect 42140 15986 42420 15988
rect 42140 15934 42142 15986
rect 42194 15934 42420 15986
rect 42140 15932 42420 15934
rect 42588 16604 42756 16660
rect 42140 15922 42196 15932
rect 42028 15586 42084 15596
rect 41916 15202 41972 15214
rect 41916 15150 41918 15202
rect 41970 15150 41972 15202
rect 41916 14980 41972 15150
rect 41916 14914 41972 14924
rect 41804 14478 41806 14530
rect 41858 14478 41860 14530
rect 41804 14466 41860 14478
rect 41916 14756 41972 14766
rect 41356 14308 41412 14318
rect 41356 14214 41412 14252
rect 41468 14306 41524 14318
rect 41468 14254 41470 14306
rect 41522 14254 41524 14306
rect 41468 14196 41524 14254
rect 41580 14308 41636 14318
rect 41580 14306 41748 14308
rect 41580 14254 41582 14306
rect 41634 14254 41748 14306
rect 41580 14252 41748 14254
rect 41580 14242 41636 14252
rect 41356 13972 41412 13982
rect 40796 13468 41188 13524
rect 41244 13524 41300 13534
rect 40572 11454 40574 11506
rect 40626 11454 40628 11506
rect 40572 11442 40628 11454
rect 40796 11284 40852 13468
rect 41244 13074 41300 13468
rect 41244 13022 41246 13074
rect 41298 13022 41300 13074
rect 41244 13010 41300 13022
rect 41356 12740 41412 13916
rect 41468 13636 41524 14140
rect 41468 13570 41524 13580
rect 41580 13412 41636 13422
rect 41580 13074 41636 13356
rect 41580 13022 41582 13074
rect 41634 13022 41636 13074
rect 41580 13010 41636 13022
rect 41356 12684 41636 12740
rect 40796 11218 40852 11228
rect 41468 12066 41524 12078
rect 41468 12014 41470 12066
rect 41522 12014 41524 12066
rect 41468 11284 41524 12014
rect 41580 11506 41636 12684
rect 41580 11454 41582 11506
rect 41634 11454 41636 11506
rect 41580 11442 41636 11454
rect 41468 11218 41524 11228
rect 41132 11170 41188 11182
rect 41132 11118 41134 11170
rect 41186 11118 41188 11170
rect 39340 10834 40068 10836
rect 39340 10782 39342 10834
rect 39394 10782 40068 10834
rect 39340 10780 40068 10782
rect 39340 10770 39396 10780
rect 39452 10612 39508 10622
rect 39452 10518 39508 10556
rect 40012 10610 40068 10780
rect 40012 10558 40014 10610
rect 40066 10558 40068 10610
rect 40012 10546 40068 10558
rect 40236 11060 40292 11070
rect 40236 10612 40292 11004
rect 41132 10836 41188 11118
rect 41692 11060 41748 14252
rect 41916 14084 41972 14700
rect 41916 14028 42084 14084
rect 41916 13860 41972 13870
rect 41916 13766 41972 13804
rect 41692 10994 41748 11004
rect 41804 13748 41860 13758
rect 41580 10836 41636 10846
rect 41804 10836 41860 13692
rect 42028 13076 42084 14028
rect 42252 13972 42308 15932
rect 42476 15876 42532 15886
rect 42364 15764 42420 15774
rect 42364 15538 42420 15708
rect 42364 15486 42366 15538
rect 42418 15486 42420 15538
rect 42364 15474 42420 15486
rect 42476 15428 42532 15820
rect 42476 15362 42532 15372
rect 42476 15204 42532 15214
rect 42476 15092 42532 15148
rect 42476 15026 42532 15036
rect 42588 14532 42644 16604
rect 43260 16548 43316 16828
rect 43148 16492 43316 16548
rect 42924 16324 42980 16334
rect 42924 16098 42980 16268
rect 42924 16046 42926 16098
rect 42978 16046 42980 16098
rect 42924 16034 42980 16046
rect 42700 15986 42756 15998
rect 42700 15934 42702 15986
rect 42754 15934 42756 15986
rect 42700 15204 42756 15934
rect 42812 15876 42868 15886
rect 42812 15782 42868 15820
rect 42812 15428 42868 15438
rect 42812 15334 42868 15372
rect 42700 15138 42756 15148
rect 43148 15090 43204 16492
rect 43260 16324 43316 16362
rect 43260 16258 43316 16268
rect 43148 15038 43150 15090
rect 43202 15038 43204 15090
rect 43148 15026 43204 15038
rect 43260 15652 43316 15662
rect 43260 15202 43316 15596
rect 43372 15316 43428 17164
rect 43708 16884 43764 18172
rect 44156 18116 44212 18126
rect 44156 17666 44212 18060
rect 44380 17892 44436 17930
rect 44380 17826 44436 17836
rect 44156 17614 44158 17666
rect 44210 17614 44212 17666
rect 44156 17602 44212 17614
rect 43932 17554 43988 17566
rect 43932 17502 43934 17554
rect 43986 17502 43988 17554
rect 43932 17332 43988 17502
rect 43932 17266 43988 17276
rect 44380 17556 44436 17566
rect 43932 17108 43988 17118
rect 43932 17106 44100 17108
rect 43932 17054 43934 17106
rect 43986 17054 44100 17106
rect 43932 17052 44100 17054
rect 43932 17042 43988 17052
rect 43932 16884 43988 16894
rect 43764 16882 43988 16884
rect 43764 16830 43934 16882
rect 43986 16830 43988 16882
rect 43764 16828 43988 16830
rect 43708 16752 43764 16828
rect 43932 16818 43988 16828
rect 43596 16212 43652 16222
rect 43484 16100 43540 16110
rect 43484 16006 43540 16044
rect 43596 15428 43652 16156
rect 43708 15652 43764 15662
rect 43708 15538 43764 15596
rect 43708 15486 43710 15538
rect 43762 15486 43764 15538
rect 43708 15474 43764 15486
rect 43372 15260 43540 15316
rect 43260 15150 43262 15202
rect 43314 15150 43316 15202
rect 43260 14756 43316 15150
rect 43260 14690 43316 14700
rect 42812 14532 42868 14542
rect 43148 14532 43204 14542
rect 42588 14530 42756 14532
rect 42588 14478 42590 14530
rect 42642 14478 42756 14530
rect 42588 14476 42756 14478
rect 42588 14466 42644 14476
rect 42588 13972 42644 13982
rect 42252 13970 42644 13972
rect 42252 13918 42590 13970
rect 42642 13918 42644 13970
rect 42252 13916 42644 13918
rect 42588 13906 42644 13916
rect 42028 13010 42084 13020
rect 42140 13746 42196 13758
rect 42140 13694 42142 13746
rect 42194 13694 42196 13746
rect 42140 12964 42196 13694
rect 42476 13748 42532 13758
rect 42140 12898 42196 12908
rect 42252 13636 42308 13646
rect 41916 12740 41972 12750
rect 41916 11396 41972 12684
rect 42028 12404 42084 12414
rect 42252 12404 42308 13580
rect 42028 12402 42308 12404
rect 42028 12350 42030 12402
rect 42082 12350 42308 12402
rect 42028 12348 42308 12350
rect 42364 12850 42420 12862
rect 42364 12798 42366 12850
rect 42418 12798 42420 12850
rect 42028 12338 42084 12348
rect 42364 12180 42420 12798
rect 41916 11340 42196 11396
rect 41132 10834 41860 10836
rect 41132 10782 41582 10834
rect 41634 10782 41860 10834
rect 41132 10780 41860 10782
rect 41916 11172 41972 11182
rect 41580 10770 41636 10780
rect 41916 10724 41972 11116
rect 42028 11170 42084 11182
rect 42028 11118 42030 11170
rect 42082 11118 42084 11170
rect 42028 11060 42084 11118
rect 42028 10836 42084 11004
rect 42028 10770 42084 10780
rect 40236 10480 40292 10556
rect 41804 10668 41972 10724
rect 39340 10388 39396 10398
rect 40572 10388 40628 10398
rect 39116 9762 39172 9772
rect 39228 10386 39396 10388
rect 39228 10334 39342 10386
rect 39394 10334 39396 10386
rect 39228 10332 39396 10334
rect 38668 9604 38724 9614
rect 38444 9436 38612 9492
rect 38444 9268 38500 9278
rect 38332 9266 38500 9268
rect 38332 9214 38446 9266
rect 38498 9214 38500 9266
rect 38332 9212 38500 9214
rect 38444 9202 38500 9212
rect 38220 9044 38276 9054
rect 38220 8950 38276 8988
rect 38332 9042 38388 9054
rect 38332 8990 38334 9042
rect 38386 8990 38388 9042
rect 37772 8932 37828 8942
rect 37772 8484 37828 8876
rect 37772 7700 37828 8428
rect 37884 8036 37940 8046
rect 37884 7942 37940 7980
rect 38332 8036 38388 8990
rect 38332 7970 38388 7980
rect 38444 8148 38500 8158
rect 37884 7700 37940 7710
rect 37772 7698 37940 7700
rect 37772 7646 37886 7698
rect 37938 7646 37940 7698
rect 37772 7644 37940 7646
rect 37884 7634 37940 7644
rect 38332 7700 38388 7710
rect 38444 7700 38500 8092
rect 38332 7698 38500 7700
rect 38332 7646 38334 7698
rect 38386 7646 38500 7698
rect 38332 7644 38500 7646
rect 37436 7362 37492 7374
rect 37436 7310 37438 7362
rect 37490 7310 37492 7362
rect 36876 3668 36932 4284
rect 36876 3602 36932 3612
rect 37100 6580 37156 6590
rect 37100 5796 37156 6524
rect 37436 6468 37492 7310
rect 37324 6466 37492 6468
rect 37324 6414 37438 6466
rect 37490 6414 37492 6466
rect 37324 6412 37492 6414
rect 37100 3666 37156 5740
rect 37212 5906 37268 5918
rect 37212 5854 37214 5906
rect 37266 5854 37268 5906
rect 37212 5236 37268 5854
rect 37212 5170 37268 5180
rect 37324 5908 37380 6412
rect 37436 6402 37492 6412
rect 37100 3614 37102 3666
rect 37154 3614 37156 3666
rect 37100 3602 37156 3614
rect 37324 3668 37380 5852
rect 37660 5010 37716 7532
rect 37884 7364 37940 7374
rect 37884 5906 37940 7308
rect 38332 6804 38388 7644
rect 38332 6738 38388 6748
rect 37884 5854 37886 5906
rect 37938 5854 37940 5906
rect 37772 5124 37828 5134
rect 37772 5030 37828 5068
rect 37660 4958 37662 5010
rect 37714 4958 37716 5010
rect 37660 4946 37716 4958
rect 37436 4900 37492 4910
rect 37436 4898 37604 4900
rect 37436 4846 37438 4898
rect 37490 4846 37604 4898
rect 37436 4844 37604 4846
rect 37436 4834 37492 4844
rect 37436 4564 37492 4574
rect 37436 4470 37492 4508
rect 37548 4452 37604 4844
rect 37548 4386 37604 4396
rect 37884 4340 37940 5854
rect 37996 6692 38052 6702
rect 37996 4562 38052 6636
rect 38220 6690 38276 6702
rect 38220 6638 38222 6690
rect 38274 6638 38276 6690
rect 38220 5236 38276 6638
rect 38556 6692 38612 9436
rect 38668 8932 38724 9548
rect 39228 9268 39284 10332
rect 39340 10322 39396 10332
rect 40348 10386 40628 10388
rect 40348 10334 40574 10386
rect 40626 10334 40628 10386
rect 40348 10332 40628 10334
rect 40012 9828 40068 9838
rect 40068 9772 40180 9828
rect 40012 9734 40068 9772
rect 39900 9714 39956 9726
rect 39900 9662 39902 9714
rect 39954 9662 39956 9714
rect 39340 9604 39396 9614
rect 39340 9510 39396 9548
rect 39900 9492 39956 9662
rect 40124 9492 40180 9772
rect 40236 9716 40292 9726
rect 40348 9716 40404 10332
rect 40572 10322 40628 10332
rect 40684 9828 40740 9838
rect 41468 9828 41524 9838
rect 40684 9826 40852 9828
rect 40684 9774 40686 9826
rect 40738 9774 40852 9826
rect 40684 9772 40852 9774
rect 40684 9762 40740 9772
rect 40236 9714 40348 9716
rect 40236 9662 40238 9714
rect 40290 9662 40348 9714
rect 40236 9660 40348 9662
rect 40236 9650 40292 9660
rect 40348 9584 40404 9660
rect 40124 9436 40404 9492
rect 39900 9426 39956 9436
rect 38780 9266 39284 9268
rect 38780 9214 39230 9266
rect 39282 9214 39284 9266
rect 38780 9212 39284 9214
rect 38780 9042 38836 9212
rect 38780 8990 38782 9042
rect 38834 8990 38836 9042
rect 38780 8978 38836 8990
rect 38668 8866 38724 8876
rect 39004 8260 39060 8270
rect 39004 8166 39060 8204
rect 38780 8148 38836 8158
rect 39116 8148 39172 9212
rect 39228 9202 39284 9212
rect 40348 9268 40404 9436
rect 39340 9156 39396 9166
rect 39340 9062 39396 9100
rect 39676 9154 39732 9166
rect 39676 9102 39678 9154
rect 39730 9102 39732 9154
rect 40348 9136 40404 9212
rect 39452 9044 39508 9054
rect 39228 8372 39284 8382
rect 39228 8278 39284 8316
rect 39452 8260 39508 8988
rect 39676 8372 39732 9102
rect 39676 8306 39732 8316
rect 40796 8372 40852 9772
rect 40908 9268 40964 9278
rect 40908 9174 40964 9212
rect 40796 8260 40852 8316
rect 40908 8260 40964 8270
rect 40796 8258 40964 8260
rect 40796 8206 40910 8258
rect 40962 8206 40964 8258
rect 40796 8204 40964 8206
rect 39452 8194 39508 8204
rect 40908 8194 40964 8204
rect 41132 8260 41188 8270
rect 41132 8166 41188 8204
rect 41356 8260 41412 8270
rect 41468 8260 41524 9772
rect 41692 9828 41748 9838
rect 41692 9266 41748 9772
rect 41692 9214 41694 9266
rect 41746 9214 41748 9266
rect 41692 9202 41748 9214
rect 41356 8258 41524 8260
rect 41356 8206 41358 8258
rect 41410 8206 41524 8258
rect 41356 8204 41524 8206
rect 41356 8194 41412 8204
rect 39340 8148 39396 8158
rect 39116 8146 39396 8148
rect 39116 8094 39342 8146
rect 39394 8094 39396 8146
rect 39116 8092 39396 8094
rect 38780 8054 38836 8092
rect 39340 8082 39396 8092
rect 39900 8148 39956 8158
rect 39900 8034 39956 8092
rect 39900 7982 39902 8034
rect 39954 7982 39956 8034
rect 39900 7028 39956 7982
rect 41468 7700 41524 8204
rect 41580 8146 41636 8158
rect 41580 8094 41582 8146
rect 41634 8094 41636 8146
rect 41580 7812 41636 8094
rect 41580 7746 41636 7756
rect 41468 7634 41524 7644
rect 39900 6962 39956 6972
rect 38556 6626 38612 6636
rect 38780 6692 38836 6702
rect 38780 6598 38836 6636
rect 41132 6466 41188 6478
rect 41132 6414 41134 6466
rect 41186 6414 41188 6466
rect 38220 5122 38276 5180
rect 40124 6018 40180 6030
rect 40124 5966 40126 6018
rect 40178 5966 40180 6018
rect 38220 5070 38222 5122
rect 38274 5070 38276 5122
rect 38220 5058 38276 5070
rect 38892 5122 38948 5134
rect 38892 5070 38894 5122
rect 38946 5070 38948 5122
rect 37996 4510 37998 4562
rect 38050 4510 38052 4562
rect 37996 4498 38052 4510
rect 38444 5012 38500 5022
rect 38444 4562 38500 4956
rect 38444 4510 38446 4562
rect 38498 4510 38500 4562
rect 37996 4340 38052 4350
rect 37884 4284 37996 4340
rect 37548 3668 37604 3678
rect 37324 3666 37604 3668
rect 37324 3614 37550 3666
rect 37602 3614 37604 3666
rect 37324 3612 37604 3614
rect 37548 3602 37604 3612
rect 37996 3666 38052 4284
rect 37996 3614 37998 3666
rect 38050 3614 38052 3666
rect 37996 3602 38052 3614
rect 38444 3666 38500 4510
rect 38780 4564 38836 4574
rect 38780 4470 38836 4508
rect 38892 4116 38948 5070
rect 40124 4564 40180 5966
rect 40908 6020 40964 6030
rect 40908 5926 40964 5964
rect 40124 4498 40180 4508
rect 41132 4898 41188 6414
rect 41132 4846 41134 4898
rect 41186 4846 41188 4898
rect 41132 4564 41188 4846
rect 41132 4498 41188 4508
rect 39340 4452 39396 4462
rect 39340 4358 39396 4396
rect 39452 4450 39508 4462
rect 39452 4398 39454 4450
rect 39506 4398 39508 4450
rect 39452 4340 39508 4398
rect 39452 4274 39508 4284
rect 40012 4340 40068 4350
rect 40012 4246 40068 4284
rect 39452 4116 39508 4126
rect 38892 4114 39508 4116
rect 38892 4062 39454 4114
rect 39506 4062 39508 4114
rect 38892 4060 39508 4062
rect 39452 4050 39508 4060
rect 38444 3614 38446 3666
rect 38498 3614 38500 3666
rect 38444 3602 38500 3614
rect 33852 3502 33854 3554
rect 33906 3502 33908 3554
rect 33852 3490 33908 3502
rect 40012 3556 40068 3566
rect 40012 3462 40068 3500
rect 40908 3556 40964 3566
rect 40908 3462 40964 3500
rect 39116 3442 39172 3454
rect 39116 3390 39118 3442
rect 39170 3390 39172 3442
rect 39116 3388 39172 3390
rect 39004 3332 39172 3388
rect 41804 3332 41860 10668
rect 42140 10612 42196 11340
rect 42364 10836 42420 12124
rect 42364 10770 42420 10780
rect 42476 10834 42532 13692
rect 42700 13636 42756 14476
rect 42812 14530 42980 14532
rect 42812 14478 42814 14530
rect 42866 14478 42980 14530
rect 42812 14476 42980 14478
rect 42812 14466 42868 14476
rect 42812 14306 42868 14318
rect 42812 14254 42814 14306
rect 42866 14254 42868 14306
rect 42812 13860 42868 14254
rect 42924 13972 42980 14476
rect 43204 14476 43428 14532
rect 43148 14400 43204 14476
rect 42924 13906 42980 13916
rect 43260 13972 43316 13982
rect 42812 13794 42868 13804
rect 42700 13570 42756 13580
rect 42924 13748 42980 13758
rect 42924 13634 42980 13692
rect 42924 13582 42926 13634
rect 42978 13582 42980 13634
rect 42924 13524 42980 13582
rect 42924 13458 42980 13468
rect 42924 13076 42980 13086
rect 42700 12962 42756 12974
rect 42700 12910 42702 12962
rect 42754 12910 42756 12962
rect 42700 12516 42756 12910
rect 42924 12964 42980 13020
rect 42924 12962 43092 12964
rect 42924 12910 42926 12962
rect 42978 12910 43092 12962
rect 42924 12908 43092 12910
rect 42924 12898 42980 12908
rect 42700 12450 42756 12460
rect 42812 12738 42868 12750
rect 42812 12686 42814 12738
rect 42866 12686 42868 12738
rect 42812 12402 42868 12686
rect 42812 12350 42814 12402
rect 42866 12350 42868 12402
rect 42812 12338 42868 12350
rect 42588 12178 42644 12190
rect 42588 12126 42590 12178
rect 42642 12126 42644 12178
rect 42588 11732 42644 12126
rect 42700 12068 42756 12078
rect 42700 11974 42756 12012
rect 42588 11676 42868 11732
rect 42812 11618 42868 11676
rect 42812 11566 42814 11618
rect 42866 11566 42868 11618
rect 42812 11554 42868 11566
rect 42924 11394 42980 11406
rect 42924 11342 42926 11394
rect 42978 11342 42980 11394
rect 42924 11284 42980 11342
rect 42924 11218 42980 11228
rect 42476 10782 42478 10834
rect 42530 10782 42532 10834
rect 42476 10770 42532 10782
rect 42924 10836 42980 10846
rect 43036 10836 43092 12908
rect 43260 12404 43316 13916
rect 43372 13746 43428 14476
rect 43372 13694 43374 13746
rect 43426 13694 43428 13746
rect 43372 13682 43428 13694
rect 43484 13748 43540 15260
rect 43484 13682 43540 13692
rect 43484 13300 43540 13310
rect 43484 13074 43540 13244
rect 43484 13022 43486 13074
rect 43538 13022 43540 13074
rect 43484 13010 43540 13022
rect 43260 12348 43540 12404
rect 43260 12180 43316 12190
rect 43260 12178 43428 12180
rect 43260 12126 43262 12178
rect 43314 12126 43428 12178
rect 43260 12124 43428 12126
rect 43260 12114 43316 12124
rect 43148 11620 43204 11630
rect 43148 11526 43204 11564
rect 43260 11508 43316 11518
rect 43260 11414 43316 11452
rect 43372 11284 43428 12124
rect 42924 10834 43092 10836
rect 42924 10782 42926 10834
rect 42978 10782 43092 10834
rect 42924 10780 43092 10782
rect 43148 11228 43428 11284
rect 42924 10770 42980 10780
rect 41916 10556 42196 10612
rect 41916 10498 41972 10556
rect 41916 10446 41918 10498
rect 41970 10446 41972 10498
rect 41916 10434 41972 10446
rect 43148 10052 43204 11228
rect 43484 11172 43540 12348
rect 43596 11508 43652 15372
rect 43820 14980 43876 14990
rect 43708 13748 43764 13758
rect 43708 13654 43764 13692
rect 43708 12404 43764 12414
rect 43820 12404 43876 14924
rect 44044 14980 44100 17052
rect 44156 16658 44212 16670
rect 44156 16606 44158 16658
rect 44210 16606 44212 16658
rect 44156 16324 44212 16606
rect 44156 16210 44212 16268
rect 44156 16158 44158 16210
rect 44210 16158 44212 16210
rect 44156 16146 44212 16158
rect 44380 16322 44436 17500
rect 44492 16882 44548 18396
rect 44604 17108 44660 18732
rect 44828 18564 44884 18574
rect 44716 18340 44772 18350
rect 44716 17666 44772 18284
rect 44716 17614 44718 17666
rect 44770 17614 44772 17666
rect 44716 17602 44772 17614
rect 44828 17556 44884 18508
rect 44940 18450 44996 18956
rect 44940 18398 44942 18450
rect 44994 18398 44996 18450
rect 44940 18386 44996 18398
rect 44828 17490 44884 17500
rect 44716 17442 44772 17454
rect 44716 17390 44718 17442
rect 44770 17390 44772 17442
rect 44716 17220 44772 17390
rect 44716 17164 44884 17220
rect 44604 17052 44772 17108
rect 44492 16830 44494 16882
rect 44546 16830 44548 16882
rect 44716 16996 44772 17052
rect 44716 16864 44772 16940
rect 44492 16548 44548 16830
rect 44492 16492 44772 16548
rect 44380 16270 44382 16322
rect 44434 16270 44436 16322
rect 44156 15988 44212 15998
rect 44156 15894 44212 15932
rect 44268 15652 44324 15662
rect 44268 15538 44324 15596
rect 44268 15486 44270 15538
rect 44322 15486 44324 15538
rect 44268 15204 44324 15486
rect 44268 15138 44324 15148
rect 44380 15148 44436 16270
rect 44604 15428 44660 15438
rect 44604 15334 44660 15372
rect 44044 14914 44100 14924
rect 44156 15090 44212 15102
rect 44380 15092 44548 15148
rect 44156 15038 44158 15090
rect 44210 15038 44212 15090
rect 44044 14306 44100 14318
rect 44044 14254 44046 14306
rect 44098 14254 44100 14306
rect 43932 13972 43988 13982
rect 43932 13878 43988 13916
rect 44044 13970 44100 14254
rect 44044 13918 44046 13970
rect 44098 13918 44100 13970
rect 44044 13906 44100 13918
rect 43708 12402 43876 12404
rect 43708 12350 43710 12402
rect 43762 12350 43876 12402
rect 43708 12348 43876 12350
rect 43932 13636 43988 13646
rect 43708 12338 43764 12348
rect 43932 12292 43988 13580
rect 44156 13636 44212 15038
rect 44268 14420 44324 14430
rect 44268 13860 44324 14364
rect 44380 14306 44436 14318
rect 44380 14254 44382 14306
rect 44434 14254 44436 14306
rect 44380 13860 44436 14254
rect 44492 14306 44548 15092
rect 44492 14254 44494 14306
rect 44546 14254 44548 14306
rect 44492 14196 44548 14254
rect 44492 14130 44548 14140
rect 44604 14980 44660 14990
rect 44380 13804 44548 13860
rect 44268 13794 44324 13804
rect 44380 13636 44436 13646
rect 44156 13634 44436 13636
rect 44156 13582 44382 13634
rect 44434 13582 44436 13634
rect 44156 13580 44436 13582
rect 44156 13300 44212 13580
rect 44380 13570 44436 13580
rect 44156 13234 44212 13244
rect 44156 12962 44212 12974
rect 44156 12910 44158 12962
rect 44210 12910 44212 12962
rect 44156 12852 44212 12910
rect 44156 12786 44212 12796
rect 44380 12962 44436 12974
rect 44380 12910 44382 12962
rect 44434 12910 44436 12962
rect 44380 12852 44436 12910
rect 44380 12786 44436 12796
rect 44268 12404 44324 12414
rect 43820 12236 43988 12292
rect 44044 12402 44324 12404
rect 44044 12350 44270 12402
rect 44322 12350 44324 12402
rect 44044 12348 44324 12350
rect 43596 11452 43764 11508
rect 43260 11116 43540 11172
rect 43596 11284 43652 11294
rect 43260 10834 43316 11116
rect 43260 10782 43262 10834
rect 43314 10782 43316 10834
rect 43260 10770 43316 10782
rect 43148 9986 43204 9996
rect 41916 9940 41972 9950
rect 41916 9846 41972 9884
rect 42140 9826 42196 9838
rect 42140 9774 42142 9826
rect 42194 9774 42196 9826
rect 42140 9268 42196 9774
rect 42812 9828 42868 9838
rect 42812 9734 42868 9772
rect 42476 9716 42532 9726
rect 42700 9716 42756 9726
rect 42476 9622 42532 9660
rect 42588 9714 42756 9716
rect 42588 9662 42702 9714
rect 42754 9662 42756 9714
rect 42588 9660 42756 9662
rect 42140 9202 42196 9212
rect 42476 9380 42532 9390
rect 42476 9154 42532 9324
rect 42476 9102 42478 9154
rect 42530 9102 42532 9154
rect 42476 9090 42532 9102
rect 42028 9042 42084 9054
rect 42028 8990 42030 9042
rect 42082 8990 42084 9042
rect 42028 8484 42084 8990
rect 42364 8484 42420 8494
rect 42084 8428 42196 8484
rect 42028 8418 42084 8428
rect 42140 8370 42196 8428
rect 42140 8318 42142 8370
rect 42194 8318 42196 8370
rect 42140 8306 42196 8318
rect 41916 8260 41972 8270
rect 41916 6914 41972 8204
rect 42364 7364 42420 8428
rect 42588 8372 42644 9660
rect 42700 9604 42756 9660
rect 43484 9604 43540 9614
rect 42700 9602 43540 9604
rect 42700 9550 43486 9602
rect 43538 9550 43540 9602
rect 42700 9548 43540 9550
rect 43484 9538 43540 9548
rect 42924 9380 42980 9390
rect 43596 9380 43652 11228
rect 42924 9154 42980 9324
rect 43484 9324 43652 9380
rect 43372 9156 43428 9166
rect 42924 9102 42926 9154
rect 42978 9102 42980 9154
rect 42924 8820 42980 9102
rect 42924 8754 42980 8764
rect 43036 9154 43428 9156
rect 43036 9102 43374 9154
rect 43426 9102 43428 9154
rect 43036 9100 43428 9102
rect 42924 8484 42980 8494
rect 42924 8390 42980 8428
rect 42476 7700 42532 7710
rect 42476 7606 42532 7644
rect 42588 7476 42644 8316
rect 42700 8260 42756 8270
rect 42700 8166 42756 8204
rect 42700 7812 42756 7822
rect 42700 7698 42756 7756
rect 42700 7646 42702 7698
rect 42754 7646 42756 7698
rect 42700 7634 42756 7646
rect 42812 7700 42868 7710
rect 43036 7700 43092 9100
rect 43372 9090 43428 9100
rect 43148 8932 43204 8942
rect 43484 8932 43540 9324
rect 43148 8370 43204 8876
rect 43372 8876 43540 8932
rect 43596 9042 43652 9054
rect 43596 8990 43598 9042
rect 43650 8990 43652 9042
rect 43148 8318 43150 8370
rect 43202 8318 43204 8370
rect 43148 8306 43204 8318
rect 43260 8820 43316 8830
rect 42812 7698 43092 7700
rect 42812 7646 42814 7698
rect 42866 7646 43092 7698
rect 42812 7644 43092 7646
rect 42812 7634 42868 7644
rect 42924 7476 42980 7486
rect 42588 7474 42980 7476
rect 42588 7422 42926 7474
rect 42978 7422 42980 7474
rect 42588 7420 42980 7422
rect 42924 7410 42980 7420
rect 42364 7308 42756 7364
rect 41916 6862 41918 6914
rect 41970 6862 41972 6914
rect 41916 6850 41972 6862
rect 42700 6802 42756 7308
rect 42700 6750 42702 6802
rect 42754 6750 42756 6802
rect 42700 6738 42756 6750
rect 43036 6468 43092 6478
rect 43260 6468 43316 8764
rect 43372 7700 43428 8876
rect 43596 8482 43652 8990
rect 43596 8430 43598 8482
rect 43650 8430 43652 8482
rect 43596 8418 43652 8430
rect 43372 7634 43428 7644
rect 43484 8260 43540 8270
rect 43708 8260 43764 11452
rect 43820 10834 43876 12236
rect 43932 11394 43988 11406
rect 43932 11342 43934 11394
rect 43986 11342 43988 11394
rect 43932 11284 43988 11342
rect 44044 11396 44100 12348
rect 44268 12338 44324 12348
rect 44492 12292 44548 13804
rect 44492 12226 44548 12236
rect 44604 12068 44660 14924
rect 44716 14532 44772 16492
rect 44828 15428 44884 17164
rect 45052 15652 45108 19516
rect 45276 19572 45332 24220
rect 45388 24164 45444 28366
rect 45612 27972 45668 27982
rect 45612 27858 45668 27916
rect 45612 27806 45614 27858
rect 45666 27806 45668 27858
rect 45612 27794 45668 27806
rect 45724 27746 45780 28476
rect 45724 27694 45726 27746
rect 45778 27694 45780 27746
rect 45500 27634 45556 27646
rect 45500 27582 45502 27634
rect 45554 27582 45556 27634
rect 45500 25508 45556 27582
rect 45612 27524 45668 27534
rect 45612 26962 45668 27468
rect 45724 27076 45780 27694
rect 46060 27076 46116 27086
rect 45724 27074 46116 27076
rect 45724 27022 46062 27074
rect 46114 27022 46116 27074
rect 45724 27020 46116 27022
rect 46060 27010 46116 27020
rect 45612 26910 45614 26962
rect 45666 26910 45668 26962
rect 45612 26898 45668 26910
rect 46284 26908 46340 29596
rect 46508 29586 46564 29596
rect 46732 30098 46788 30110
rect 46732 30046 46734 30098
rect 46786 30046 46788 30098
rect 46732 29540 46788 30046
rect 46732 29484 47012 29540
rect 46620 29428 46676 29438
rect 46620 29334 46676 29372
rect 46620 28868 46676 28878
rect 46620 28754 46676 28812
rect 46620 28702 46622 28754
rect 46674 28702 46676 28754
rect 46620 28690 46676 28702
rect 46956 27970 47012 29484
rect 47180 29316 47236 30156
rect 47292 29986 47348 29998
rect 47292 29934 47294 29986
rect 47346 29934 47348 29986
rect 47292 29540 47348 29934
rect 47628 29988 47684 29998
rect 47628 29894 47684 29932
rect 47404 29652 47460 29662
rect 47404 29558 47460 29596
rect 47292 29474 47348 29484
rect 47180 29250 47236 29260
rect 47740 29426 47796 29438
rect 47740 29374 47742 29426
rect 47794 29374 47796 29426
rect 47740 28868 47796 29374
rect 47740 28802 47796 28812
rect 47964 29428 48020 29438
rect 47180 28418 47236 28430
rect 47180 28366 47182 28418
rect 47234 28366 47236 28418
rect 46956 27918 46958 27970
rect 47010 27918 47012 27970
rect 45836 26852 45892 26862
rect 45836 26758 45892 26796
rect 45948 26850 46004 26862
rect 45948 26798 45950 26850
rect 46002 26798 46004 26850
rect 45836 26290 45892 26302
rect 45836 26238 45838 26290
rect 45890 26238 45892 26290
rect 45836 26180 45892 26238
rect 45836 26114 45892 26124
rect 45500 25442 45556 25452
rect 45500 25284 45556 25294
rect 45500 24722 45556 25228
rect 45836 25282 45892 25294
rect 45836 25230 45838 25282
rect 45890 25230 45892 25282
rect 45500 24670 45502 24722
rect 45554 24670 45556 24722
rect 45500 24658 45556 24670
rect 45724 24722 45780 24734
rect 45724 24670 45726 24722
rect 45778 24670 45780 24722
rect 45388 24098 45444 24108
rect 45612 24498 45668 24510
rect 45612 24446 45614 24498
rect 45666 24446 45668 24498
rect 45388 23716 45444 23726
rect 45388 23622 45444 23660
rect 45612 23716 45668 24446
rect 45724 24500 45780 24670
rect 45724 24434 45780 24444
rect 45612 23650 45668 23660
rect 45724 23828 45780 23838
rect 45500 23268 45556 23278
rect 45500 23044 45556 23212
rect 45500 22950 45556 22988
rect 45612 22932 45668 22942
rect 45388 22260 45444 22336
rect 45444 22204 45556 22260
rect 45388 22194 45444 22204
rect 45500 21812 45556 22204
rect 45500 21746 45556 21756
rect 45388 21700 45444 21710
rect 45388 21606 45444 21644
rect 45388 21140 45444 21150
rect 45388 20914 45444 21084
rect 45388 20862 45390 20914
rect 45442 20862 45444 20914
rect 45388 20850 45444 20862
rect 45500 20244 45556 20282
rect 45500 20178 45556 20188
rect 45276 19506 45332 19516
rect 45388 20130 45444 20142
rect 45388 20078 45390 20130
rect 45442 20078 45444 20130
rect 45164 19348 45220 19358
rect 45164 17556 45220 19292
rect 45276 19236 45332 19246
rect 45388 19236 45444 20078
rect 45500 20020 45556 20030
rect 45500 19926 45556 19964
rect 45612 19908 45668 22876
rect 45612 19842 45668 19852
rect 45388 19180 45556 19236
rect 45276 19124 45332 19180
rect 45276 19068 45444 19124
rect 45388 19010 45444 19068
rect 45388 18958 45390 19010
rect 45442 18958 45444 19010
rect 45388 18946 45444 18958
rect 45164 17106 45220 17500
rect 45164 17054 45166 17106
rect 45218 17054 45220 17106
rect 45164 17042 45220 17054
rect 45388 17108 45444 17118
rect 45388 16210 45444 17052
rect 45388 16158 45390 16210
rect 45442 16158 45444 16210
rect 45388 16146 45444 16158
rect 45500 16772 45556 19180
rect 45612 18788 45668 18798
rect 45724 18788 45780 23772
rect 45836 23492 45892 25230
rect 45948 24836 46004 26798
rect 45948 24770 46004 24780
rect 46060 26852 46340 26908
rect 46396 27858 46452 27870
rect 46396 27806 46398 27858
rect 46450 27806 46452 27858
rect 46396 26964 46452 27806
rect 46844 27858 46900 27870
rect 46844 27806 46846 27858
rect 46898 27806 46900 27858
rect 46844 27748 46900 27806
rect 46956 27860 47012 27918
rect 46956 27794 47012 27804
rect 47068 28084 47124 28094
rect 46844 27682 46900 27692
rect 46956 27636 47012 27646
rect 46956 27542 47012 27580
rect 46060 24834 46116 26852
rect 46172 26290 46228 26302
rect 46172 26238 46174 26290
rect 46226 26238 46228 26290
rect 46172 26068 46228 26238
rect 46172 26002 46228 26012
rect 46060 24782 46062 24834
rect 46114 24782 46116 24834
rect 46060 24770 46116 24782
rect 46172 25394 46228 25406
rect 46172 25342 46174 25394
rect 46226 25342 46228 25394
rect 45948 24612 46004 24622
rect 45948 24518 46004 24556
rect 45836 23426 45892 23436
rect 45948 23828 46004 23838
rect 45948 23378 46004 23772
rect 45948 23326 45950 23378
rect 46002 23326 46004 23378
rect 45948 23314 46004 23326
rect 45836 23268 45892 23278
rect 45836 18900 45892 23212
rect 46172 23044 46228 25342
rect 46284 23826 46340 23838
rect 46284 23774 46286 23826
rect 46338 23774 46340 23826
rect 46284 23492 46340 23774
rect 46284 23426 46340 23436
rect 46396 23268 46452 26908
rect 46620 27524 46676 27534
rect 46508 26740 46564 26750
rect 46508 24500 46564 26684
rect 46620 26514 46676 27468
rect 47068 27074 47124 28028
rect 47180 27748 47236 28366
rect 47628 28420 47684 28430
rect 47628 28418 47796 28420
rect 47628 28366 47630 28418
rect 47682 28366 47796 28418
rect 47628 28364 47796 28366
rect 47628 28354 47684 28364
rect 47628 27860 47684 27870
rect 47628 27766 47684 27804
rect 47180 27682 47236 27692
rect 47628 27636 47684 27646
rect 47068 27022 47070 27074
rect 47122 27022 47124 27074
rect 47068 27010 47124 27022
rect 47516 27524 47572 27534
rect 46620 26462 46622 26514
rect 46674 26462 46676 26514
rect 46620 26450 46676 26462
rect 46844 26850 46900 26862
rect 46844 26798 46846 26850
rect 46898 26798 46900 26850
rect 46844 26068 46900 26798
rect 47516 26514 47572 27468
rect 47516 26462 47518 26514
rect 47570 26462 47572 26514
rect 47516 26450 47572 26462
rect 47068 26292 47124 26302
rect 47068 26198 47124 26236
rect 46844 26002 46900 26012
rect 47404 25618 47460 25630
rect 47404 25566 47406 25618
rect 47458 25566 47460 25618
rect 46844 25394 46900 25406
rect 46844 25342 46846 25394
rect 46898 25342 46900 25394
rect 46732 25284 46788 25294
rect 46732 25190 46788 25228
rect 46844 24946 46900 25342
rect 47404 25396 47460 25566
rect 47404 25330 47460 25340
rect 47628 25396 47684 27580
rect 47740 26964 47796 28364
rect 47740 26870 47796 26908
rect 47852 28082 47908 28094
rect 47852 28030 47854 28082
rect 47906 28030 47908 28082
rect 47628 25302 47684 25340
rect 47740 25508 47796 25518
rect 46844 24894 46846 24946
rect 46898 24894 46900 24946
rect 46844 24882 46900 24894
rect 46956 25284 47012 25294
rect 46956 24836 47012 25228
rect 47740 24948 47796 25452
rect 47852 25060 47908 28030
rect 47964 27972 48020 29372
rect 47964 27840 48020 27916
rect 48076 27188 48132 30940
rect 48524 30324 48580 31502
rect 48636 31556 48692 31566
rect 48636 31218 48692 31500
rect 49084 31556 49140 31566
rect 49084 31462 49140 31500
rect 50204 31556 50260 31566
rect 50764 31556 50820 31566
rect 51212 31556 51268 31566
rect 48636 31166 48638 31218
rect 48690 31166 48692 31218
rect 48636 31154 48692 31166
rect 49532 31108 49588 31118
rect 49532 31014 49588 31052
rect 49868 30996 49924 31006
rect 50204 30996 50260 31500
rect 49868 30994 50260 30996
rect 49868 30942 49870 30994
rect 49922 30942 50260 30994
rect 49868 30940 50260 30942
rect 50428 31554 50820 31556
rect 50428 31502 50766 31554
rect 50818 31502 50820 31554
rect 50428 31500 50820 31502
rect 50428 30996 50484 31500
rect 50764 31490 50820 31500
rect 51100 31554 51268 31556
rect 51100 31502 51214 31554
rect 51266 31502 51268 31554
rect 51100 31500 51268 31502
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50652 31220 50708 31230
rect 50652 31126 50708 31164
rect 48524 30268 48692 30324
rect 48524 30098 48580 30110
rect 48524 30046 48526 30098
rect 48578 30046 48580 30098
rect 48188 29988 48244 29998
rect 48524 29988 48580 30046
rect 48188 29986 48356 29988
rect 48188 29934 48190 29986
rect 48242 29934 48356 29986
rect 48188 29932 48356 29934
rect 48188 29922 48244 29932
rect 48188 29316 48244 29326
rect 48188 29222 48244 29260
rect 48188 28532 48244 28542
rect 48188 27970 48244 28476
rect 48188 27918 48190 27970
rect 48242 27918 48244 27970
rect 48188 27906 48244 27918
rect 48300 27860 48356 29932
rect 48524 29922 48580 29932
rect 48524 28868 48580 28878
rect 48412 28756 48468 28766
rect 48412 28662 48468 28700
rect 48524 28530 48580 28812
rect 48524 28478 48526 28530
rect 48578 28478 48580 28530
rect 48524 28466 48580 28478
rect 48636 28084 48692 30268
rect 49756 30212 49812 30222
rect 49308 30100 49364 30110
rect 49308 30006 49364 30044
rect 49644 30100 49700 30110
rect 49644 30006 49700 30044
rect 48748 29652 48804 29662
rect 48748 28866 48804 29596
rect 49644 29652 49700 29662
rect 49756 29652 49812 30156
rect 49700 29596 49812 29652
rect 49644 29520 49700 29596
rect 49756 29428 49812 29438
rect 49868 29428 49924 30940
rect 50428 30864 50484 30940
rect 50764 30772 50820 30782
rect 50652 30770 50820 30772
rect 50652 30718 50766 30770
rect 50818 30718 50820 30770
rect 50652 30716 50820 30718
rect 50652 30548 50708 30716
rect 50764 30706 50820 30716
rect 50652 30322 50708 30492
rect 50652 30270 50654 30322
rect 50706 30270 50708 30322
rect 50652 30258 50708 30270
rect 50876 30210 50932 30222
rect 50876 30158 50878 30210
rect 50930 30158 50932 30210
rect 50204 30100 50260 30110
rect 50204 29540 50260 30044
rect 50428 30098 50484 30110
rect 50428 30046 50430 30098
rect 50482 30046 50484 30098
rect 50428 29652 50484 30046
rect 50876 29988 50932 30158
rect 50876 29922 50932 29932
rect 50988 30212 51044 30222
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50428 29586 50484 29596
rect 49756 29426 49924 29428
rect 49756 29374 49758 29426
rect 49810 29374 49924 29426
rect 49756 29372 49924 29374
rect 49980 29484 50204 29540
rect 48748 28814 48750 28866
rect 48802 28814 48804 28866
rect 48748 28802 48804 28814
rect 48860 29314 48916 29326
rect 48860 29262 48862 29314
rect 48914 29262 48916 29314
rect 48692 28028 48804 28084
rect 48636 28018 48692 28028
rect 48300 27794 48356 27804
rect 48524 27860 48580 27870
rect 48188 27188 48244 27198
rect 48076 27132 48188 27188
rect 48188 27094 48244 27132
rect 47964 27076 48020 27086
rect 47964 25394 48020 27020
rect 47964 25342 47966 25394
rect 48018 25342 48020 25394
rect 47964 25330 48020 25342
rect 48076 26852 48132 26862
rect 48076 25172 48132 26796
rect 48524 26514 48580 27804
rect 48524 26462 48526 26514
rect 48578 26462 48580 26514
rect 48524 26450 48580 26462
rect 48636 27748 48692 27758
rect 48300 26292 48356 26302
rect 48636 26292 48692 27692
rect 48748 27188 48804 28028
rect 48860 27972 48916 29262
rect 48860 27906 48916 27916
rect 48972 29316 49028 29326
rect 48748 27132 48916 27188
rect 48300 26290 48692 26292
rect 48300 26238 48302 26290
rect 48354 26238 48692 26290
rect 48300 26236 48692 26238
rect 48300 26226 48356 26236
rect 48300 26068 48356 26078
rect 48188 25284 48244 25294
rect 48188 25190 48244 25228
rect 47852 25004 48020 25060
rect 47404 24892 47796 24948
rect 46956 24742 47012 24780
rect 47180 24836 47236 24846
rect 47180 24742 47236 24780
rect 46732 24722 46788 24734
rect 46732 24670 46734 24722
rect 46786 24670 46788 24722
rect 46732 24612 46788 24670
rect 47292 24724 47348 24734
rect 46732 24556 47012 24612
rect 46508 24444 46900 24500
rect 46620 24052 46676 24062
rect 46620 23938 46676 23996
rect 46620 23886 46622 23938
rect 46674 23886 46676 23938
rect 46620 23874 46676 23886
rect 46732 23938 46788 23950
rect 46732 23886 46734 23938
rect 46786 23886 46788 23938
rect 46620 23716 46676 23726
rect 46620 23622 46676 23660
rect 46396 23202 46452 23212
rect 46508 23492 46564 23502
rect 46060 22372 46116 22382
rect 46172 22372 46228 22988
rect 46396 23044 46452 23054
rect 46508 23044 46564 23436
rect 46396 23042 46564 23044
rect 46396 22990 46398 23042
rect 46450 22990 46564 23042
rect 46396 22988 46564 22990
rect 46396 22932 46452 22988
rect 46396 22866 46452 22876
rect 46284 22372 46340 22382
rect 46172 22370 46340 22372
rect 46172 22318 46286 22370
rect 46338 22318 46340 22370
rect 46172 22316 46340 22318
rect 45948 22148 46004 22158
rect 45948 22054 46004 22092
rect 45948 21700 46004 21710
rect 45948 21606 46004 21644
rect 45948 19124 46004 19134
rect 45948 19030 46004 19068
rect 46060 19012 46116 22316
rect 46284 22306 46340 22316
rect 46732 22372 46788 23886
rect 46844 23716 46900 24444
rect 46956 24164 47012 24556
rect 46956 24108 47124 24164
rect 46956 23940 47012 23950
rect 46956 23846 47012 23884
rect 46844 23660 47012 23716
rect 46844 23492 46900 23502
rect 46844 23378 46900 23436
rect 46844 23326 46846 23378
rect 46898 23326 46900 23378
rect 46844 22820 46900 23326
rect 46844 22754 46900 22764
rect 46732 22306 46788 22316
rect 46956 22260 47012 23660
rect 47068 23268 47124 24108
rect 47180 23828 47236 23838
rect 47180 23734 47236 23772
rect 47292 23716 47348 24668
rect 47292 23378 47348 23660
rect 47292 23326 47294 23378
rect 47346 23326 47348 23378
rect 47292 23314 47348 23326
rect 47180 23268 47236 23278
rect 47068 23212 47180 23268
rect 47180 23202 47236 23212
rect 46172 22146 46228 22158
rect 46844 22148 46900 22158
rect 46172 22094 46174 22146
rect 46226 22094 46228 22146
rect 46172 21700 46228 22094
rect 46172 21028 46228 21644
rect 46396 22146 46900 22148
rect 46396 22094 46846 22146
rect 46898 22094 46900 22146
rect 46396 22092 46900 22094
rect 46284 21588 46340 21598
rect 46396 21588 46452 22092
rect 46844 22082 46900 22092
rect 46956 21924 47012 22204
rect 46844 21868 47012 21924
rect 47180 22820 47236 22830
rect 47404 22820 47460 24892
rect 47852 24836 47908 24846
rect 47628 24612 47684 24622
rect 47628 24518 47684 24556
rect 47516 24498 47572 24510
rect 47516 24446 47518 24498
rect 47570 24446 47572 24498
rect 47516 24276 47572 24446
rect 47516 24210 47572 24220
rect 47740 24500 47796 24510
rect 47628 24052 47684 24062
rect 47740 24052 47796 24444
rect 47628 24050 47796 24052
rect 47628 23998 47630 24050
rect 47682 23998 47796 24050
rect 47628 23996 47796 23998
rect 47628 23986 47684 23996
rect 47740 23380 47796 23390
rect 47740 23286 47796 23324
rect 46284 21586 46452 21588
rect 46284 21534 46286 21586
rect 46338 21534 46452 21586
rect 46284 21532 46452 21534
rect 46732 21812 46788 21822
rect 46284 21522 46340 21532
rect 46508 21474 46564 21486
rect 46508 21422 46510 21474
rect 46562 21422 46564 21474
rect 46172 20972 46452 21028
rect 46284 20804 46340 20814
rect 46284 20710 46340 20748
rect 46396 20692 46452 20972
rect 46508 20916 46564 21422
rect 46732 21474 46788 21756
rect 46732 21422 46734 21474
rect 46786 21422 46788 21474
rect 46732 21410 46788 21422
rect 46844 21140 46900 21868
rect 46844 21074 46900 21084
rect 46956 21586 47012 21598
rect 46956 21534 46958 21586
rect 47010 21534 47012 21586
rect 46508 20860 46676 20916
rect 46508 20692 46564 20702
rect 46396 20690 46564 20692
rect 46396 20638 46510 20690
rect 46562 20638 46564 20690
rect 46396 20636 46564 20638
rect 46508 20626 46564 20636
rect 46396 20020 46452 20030
rect 46172 19908 46228 19918
rect 46172 19236 46228 19852
rect 46284 19684 46340 19694
rect 46284 19346 46340 19628
rect 46284 19294 46286 19346
rect 46338 19294 46340 19346
rect 46284 19282 46340 19294
rect 46396 19348 46452 19964
rect 46620 20020 46676 20860
rect 46732 20804 46788 20842
rect 46732 20738 46788 20748
rect 46732 20580 46788 20590
rect 46956 20580 47012 21534
rect 46732 20578 47012 20580
rect 46732 20526 46734 20578
rect 46786 20526 47012 20578
rect 46732 20524 47012 20526
rect 47068 20802 47124 20814
rect 47068 20750 47070 20802
rect 47122 20750 47124 20802
rect 46732 20514 46788 20524
rect 46620 19954 46676 19964
rect 46732 20356 46788 20366
rect 47068 20356 47124 20750
rect 46396 19282 46452 19292
rect 46732 19346 46788 20300
rect 46732 19294 46734 19346
rect 46786 19294 46788 19346
rect 46732 19282 46788 19294
rect 46956 20300 47124 20356
rect 46956 19458 47012 20300
rect 46956 19406 46958 19458
rect 47010 19406 47012 19458
rect 46172 19170 46228 19180
rect 46060 18956 46452 19012
rect 45836 18844 46004 18900
rect 45724 18732 45892 18788
rect 45612 18340 45668 18732
rect 45836 18452 45892 18732
rect 45836 18386 45892 18396
rect 45724 18340 45780 18350
rect 45612 18338 45780 18340
rect 45612 18286 45726 18338
rect 45778 18286 45780 18338
rect 45612 18284 45780 18286
rect 45724 18228 45780 18284
rect 45724 18162 45780 18172
rect 45836 18226 45892 18238
rect 45836 18174 45838 18226
rect 45890 18174 45892 18226
rect 45836 17892 45892 18174
rect 45724 17836 45892 17892
rect 45724 17554 45780 17836
rect 45724 17502 45726 17554
rect 45778 17502 45780 17554
rect 45724 17490 45780 17502
rect 45836 17108 45892 17118
rect 45052 15586 45108 15596
rect 45276 15988 45332 15998
rect 44828 15372 45108 15428
rect 44828 14532 44884 14542
rect 44716 14476 44828 14532
rect 44828 13970 44884 14476
rect 44828 13918 44830 13970
rect 44882 13918 44884 13970
rect 44828 13906 44884 13918
rect 44716 12738 44772 12750
rect 44716 12686 44718 12738
rect 44770 12686 44772 12738
rect 44716 12628 44772 12686
rect 44716 12562 44772 12572
rect 44156 12012 44660 12068
rect 44828 12178 44884 12190
rect 44828 12126 44830 12178
rect 44882 12126 44884 12178
rect 44156 11620 44212 12012
rect 44492 11844 44548 11854
rect 44156 11488 44212 11564
rect 44268 11732 44324 11742
rect 44044 11330 44100 11340
rect 43932 11218 43988 11228
rect 44268 11060 44324 11676
rect 44380 11620 44436 11630
rect 44380 11526 44436 11564
rect 44268 10994 44324 11004
rect 43820 10782 43822 10834
rect 43874 10782 43876 10834
rect 43820 10770 43876 10782
rect 44492 10834 44548 11788
rect 44492 10782 44494 10834
rect 44546 10782 44548 10834
rect 44492 10770 44548 10782
rect 44828 11618 44884 12126
rect 45052 11956 45108 15372
rect 44828 11566 44830 11618
rect 44882 11566 44884 11618
rect 44828 10724 44884 11566
rect 44940 11900 45108 11956
rect 45164 14196 45220 14206
rect 45164 13636 45220 14140
rect 45276 14084 45332 15932
rect 45500 15538 45556 16716
rect 45500 15486 45502 15538
rect 45554 15486 45556 15538
rect 45500 15474 45556 15486
rect 45724 16884 45780 16894
rect 45724 15426 45780 16828
rect 45836 16100 45892 17052
rect 45836 16034 45892 16044
rect 45724 15374 45726 15426
rect 45778 15374 45780 15426
rect 45724 15362 45780 15374
rect 45388 15090 45444 15102
rect 45388 15038 45390 15090
rect 45442 15038 45444 15090
rect 45388 14308 45444 15038
rect 45724 15092 45780 15102
rect 45500 14420 45556 14430
rect 45500 14326 45556 14364
rect 45724 14420 45780 15036
rect 45724 14354 45780 14364
rect 45836 14532 45892 14542
rect 45948 14532 46004 18844
rect 46060 17780 46116 17790
rect 46060 17666 46116 17724
rect 46060 17614 46062 17666
rect 46114 17614 46116 17666
rect 46060 16884 46116 17614
rect 46172 17668 46228 17678
rect 46172 16994 46228 17612
rect 46172 16942 46174 16994
rect 46226 16942 46228 16994
rect 46172 16930 46228 16942
rect 46060 16818 46116 16828
rect 46172 16548 46228 16558
rect 46172 15986 46228 16492
rect 46396 16100 46452 18956
rect 46620 18562 46676 18574
rect 46620 18510 46622 18562
rect 46674 18510 46676 18562
rect 46620 18452 46676 18510
rect 46620 18386 46676 18396
rect 46732 18450 46788 18462
rect 46732 18398 46734 18450
rect 46786 18398 46788 18450
rect 46732 18340 46788 18398
rect 46620 18226 46676 18238
rect 46620 18174 46622 18226
rect 46674 18174 46676 18226
rect 46620 17668 46676 18174
rect 46620 17602 46676 17612
rect 46732 17108 46788 18284
rect 46844 17108 46900 17118
rect 46732 17106 46900 17108
rect 46732 17054 46846 17106
rect 46898 17054 46900 17106
rect 46732 17052 46900 17054
rect 46844 17042 46900 17052
rect 46956 16548 47012 19406
rect 46396 16098 46564 16100
rect 46396 16046 46398 16098
rect 46450 16046 46564 16098
rect 46396 16044 46564 16046
rect 46396 16034 46452 16044
rect 46172 15934 46174 15986
rect 46226 15934 46228 15986
rect 46172 15922 46228 15934
rect 46396 15876 46452 15886
rect 46172 15316 46228 15326
rect 46172 15222 46228 15260
rect 46396 14532 46452 15820
rect 45836 14530 46004 14532
rect 45836 14478 45838 14530
rect 45890 14478 46004 14530
rect 45836 14476 46004 14478
rect 46172 14476 46452 14532
rect 45388 14242 45444 14252
rect 45500 14196 45556 14206
rect 45276 14028 45444 14084
rect 45276 13636 45332 13646
rect 45164 13634 45332 13636
rect 45164 13582 45278 13634
rect 45330 13582 45332 13634
rect 45164 13580 45332 13582
rect 45164 12516 45220 13580
rect 45276 13570 45332 13580
rect 45388 12852 45444 14028
rect 45500 13074 45556 14140
rect 45836 14084 45892 14476
rect 46172 14308 46228 14476
rect 46508 14308 46564 16044
rect 46956 15876 47012 16492
rect 47068 19684 47124 19694
rect 47068 15988 47124 19628
rect 47180 19346 47236 22764
rect 47292 22764 47460 22820
rect 47628 22930 47684 22942
rect 47628 22878 47630 22930
rect 47682 22878 47684 22930
rect 47292 22370 47348 22764
rect 47516 22708 47572 22718
rect 47292 22318 47294 22370
rect 47346 22318 47348 22370
rect 47292 22306 47348 22318
rect 47404 22652 47516 22708
rect 47404 22370 47460 22652
rect 47516 22642 47572 22652
rect 47404 22318 47406 22370
rect 47458 22318 47460 22370
rect 47404 22306 47460 22318
rect 47516 22484 47572 22494
rect 47404 22148 47460 22158
rect 47404 19908 47460 22092
rect 47516 20132 47572 22428
rect 47628 22370 47684 22878
rect 47628 22318 47630 22370
rect 47682 22318 47684 22370
rect 47628 22306 47684 22318
rect 47852 21700 47908 24780
rect 47964 24052 48020 25004
rect 48076 24946 48132 25116
rect 48076 24894 48078 24946
rect 48130 24894 48132 24946
rect 48076 24882 48132 24894
rect 48300 24724 48356 26012
rect 48636 25620 48692 26236
rect 48748 26964 48804 26974
rect 48748 26402 48804 26908
rect 48860 26740 48916 27132
rect 48860 26674 48916 26684
rect 48748 26350 48750 26402
rect 48802 26350 48804 26402
rect 48748 25732 48804 26350
rect 48748 25666 48804 25676
rect 48860 26066 48916 26078
rect 48860 26014 48862 26066
rect 48914 26014 48916 26066
rect 48860 25730 48916 26014
rect 48860 25678 48862 25730
rect 48914 25678 48916 25730
rect 48860 25666 48916 25678
rect 48636 25554 48692 25564
rect 47964 23986 48020 23996
rect 48076 24668 48356 24724
rect 48412 25284 48468 25294
rect 48076 21812 48132 24668
rect 48412 23828 48468 25228
rect 48636 25282 48692 25294
rect 48636 25230 48638 25282
rect 48690 25230 48692 25282
rect 48636 25172 48692 25230
rect 48636 25106 48692 25116
rect 48524 24610 48580 24622
rect 48524 24558 48526 24610
rect 48578 24558 48580 24610
rect 48524 24164 48580 24558
rect 48524 24098 48580 24108
rect 48748 24164 48804 24174
rect 48636 23940 48692 23950
rect 48748 23940 48804 24108
rect 48972 24052 49028 29260
rect 49644 29204 49700 29214
rect 49532 29202 49700 29204
rect 49532 29150 49646 29202
rect 49698 29150 49700 29202
rect 49532 29148 49700 29150
rect 49308 28642 49364 28654
rect 49308 28590 49310 28642
rect 49362 28590 49364 28642
rect 49308 28532 49364 28590
rect 49308 27412 49364 28476
rect 49308 27346 49364 27356
rect 49420 27858 49476 27870
rect 49420 27806 49422 27858
rect 49474 27806 49476 27858
rect 49084 27076 49140 27086
rect 49084 26982 49140 27020
rect 49308 27076 49364 27086
rect 49420 27076 49476 27806
rect 49308 27074 49476 27076
rect 49308 27022 49310 27074
rect 49362 27022 49476 27074
rect 49308 27020 49476 27022
rect 49532 27748 49588 29148
rect 49644 29138 49700 29148
rect 49756 29204 49812 29372
rect 49756 29138 49812 29148
rect 49756 28756 49812 28766
rect 49644 28196 49700 28206
rect 49644 28082 49700 28140
rect 49644 28030 49646 28082
rect 49698 28030 49700 28082
rect 49644 28018 49700 28030
rect 49756 28084 49812 28700
rect 49868 28756 49924 28766
rect 49980 28756 50036 29484
rect 50204 29474 50260 29484
rect 50316 29538 50372 29550
rect 50316 29486 50318 29538
rect 50370 29486 50372 29538
rect 50316 29428 50372 29486
rect 50316 29362 50372 29372
rect 50652 29426 50708 29438
rect 50652 29374 50654 29426
rect 50706 29374 50708 29426
rect 49868 28754 50036 28756
rect 49868 28702 49870 28754
rect 49922 28702 50036 28754
rect 49868 28700 50036 28702
rect 50428 29204 50484 29214
rect 50428 28756 50484 29148
rect 49868 28690 49924 28700
rect 50428 28662 50484 28700
rect 50652 28532 50708 29374
rect 50652 28466 50708 28476
rect 50876 28642 50932 28654
rect 50876 28590 50878 28642
rect 50930 28590 50932 28642
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50204 28084 50260 28094
rect 49756 28082 50260 28084
rect 49756 28030 50206 28082
rect 50258 28030 50260 28082
rect 49756 28028 50260 28030
rect 49756 27970 49812 28028
rect 50204 28018 50260 28028
rect 50876 28084 50932 28590
rect 49756 27918 49758 27970
rect 49810 27918 49812 27970
rect 49756 27906 49812 27918
rect 49532 27076 49588 27692
rect 50876 27300 50932 28028
rect 50876 27234 50932 27244
rect 50204 27076 50260 27086
rect 49532 27074 50260 27076
rect 49532 27022 50206 27074
rect 50258 27022 50260 27074
rect 49532 27020 50260 27022
rect 49196 26964 49252 26974
rect 49196 26870 49252 26908
rect 49196 26740 49252 26750
rect 49084 25284 49140 25294
rect 49196 25284 49252 26684
rect 49308 25508 49364 27020
rect 49532 26516 49588 26526
rect 49420 26178 49476 26190
rect 49420 26126 49422 26178
rect 49474 26126 49476 26178
rect 49420 26068 49476 26126
rect 49420 26002 49476 26012
rect 49308 25442 49364 25452
rect 49532 25618 49588 26460
rect 49868 26180 49924 26190
rect 49868 26086 49924 26124
rect 49532 25566 49534 25618
rect 49586 25566 49588 25618
rect 49532 25508 49588 25566
rect 49532 25442 49588 25452
rect 49644 25730 49700 25742
rect 49644 25678 49646 25730
rect 49698 25678 49700 25730
rect 49084 25282 49252 25284
rect 49084 25230 49086 25282
rect 49138 25230 49252 25282
rect 49084 25228 49252 25230
rect 49084 25218 49140 25228
rect 48636 23938 48804 23940
rect 48636 23886 48638 23938
rect 48690 23886 48804 23938
rect 48636 23884 48804 23886
rect 48860 23996 49028 24052
rect 49084 24052 49140 24062
rect 48636 23874 48692 23884
rect 48412 23772 48580 23828
rect 48188 23716 48244 23726
rect 48524 23716 48580 23772
rect 48188 23714 48356 23716
rect 48188 23662 48190 23714
rect 48242 23662 48356 23714
rect 48188 23660 48356 23662
rect 48524 23660 48804 23716
rect 48188 23650 48244 23660
rect 48300 23492 48356 23660
rect 48188 23044 48244 23054
rect 48188 22950 48244 22988
rect 48188 22260 48244 22270
rect 48188 22166 48244 22204
rect 48300 22148 48356 23436
rect 48748 23378 48804 23660
rect 48748 23326 48750 23378
rect 48802 23326 48804 23378
rect 48748 23314 48804 23326
rect 48860 23714 48916 23996
rect 48860 23662 48862 23714
rect 48914 23662 48916 23714
rect 48524 22930 48580 22942
rect 48524 22878 48526 22930
rect 48578 22878 48580 22930
rect 48300 22082 48356 22092
rect 48412 22370 48468 22382
rect 48412 22318 48414 22370
rect 48466 22318 48468 22370
rect 48076 21746 48132 21756
rect 48188 21812 48244 21822
rect 48412 21812 48468 22318
rect 48188 21810 48468 21812
rect 48188 21758 48190 21810
rect 48242 21758 48468 21810
rect 48188 21756 48468 21758
rect 48524 22372 48580 22878
rect 48860 22932 48916 23662
rect 48972 23826 49028 23838
rect 48972 23774 48974 23826
rect 49026 23774 49028 23826
rect 48972 23492 49028 23774
rect 48972 23426 49028 23436
rect 49084 23044 49140 23996
rect 49196 23380 49252 25228
rect 49196 23314 49252 23324
rect 49420 25284 49476 25294
rect 49084 22978 49140 22988
rect 48860 22866 48916 22876
rect 49196 22932 49252 22942
rect 49196 22596 49252 22876
rect 49196 22484 49252 22540
rect 49084 22428 49252 22484
rect 48636 22372 48692 22382
rect 48524 22370 48692 22372
rect 48524 22318 48638 22370
rect 48690 22318 48692 22370
rect 48524 22316 48692 22318
rect 48188 21746 48244 21756
rect 47740 21644 47908 21700
rect 47740 20692 47796 21644
rect 47964 21586 48020 21598
rect 48300 21588 48356 21756
rect 47964 21534 47966 21586
rect 48018 21534 48020 21586
rect 47964 21364 48020 21534
rect 47964 21298 48020 21308
rect 48076 21532 48356 21588
rect 47964 20804 48020 20814
rect 48076 20804 48132 21532
rect 48300 21362 48356 21374
rect 48300 21310 48302 21362
rect 48354 21310 48356 21362
rect 48300 21252 48356 21310
rect 48300 21186 48356 21196
rect 47964 20802 48132 20804
rect 47964 20750 47966 20802
rect 48018 20750 48132 20802
rect 47964 20748 48132 20750
rect 47964 20738 48020 20748
rect 47740 20636 47908 20692
rect 47628 20580 47684 20590
rect 47628 20578 47796 20580
rect 47628 20526 47630 20578
rect 47682 20526 47796 20578
rect 47628 20524 47796 20526
rect 47628 20514 47684 20524
rect 47516 20066 47572 20076
rect 47404 19852 47572 19908
rect 47180 19294 47182 19346
rect 47234 19294 47236 19346
rect 47180 19282 47236 19294
rect 47292 19460 47348 19470
rect 47292 18674 47348 19404
rect 47292 18622 47294 18674
rect 47346 18622 47348 18674
rect 47180 16324 47236 16334
rect 47180 16230 47236 16268
rect 47292 16100 47348 18622
rect 47404 17668 47460 17678
rect 47404 17574 47460 17612
rect 47516 17332 47572 19852
rect 47628 19458 47684 19470
rect 47628 19406 47630 19458
rect 47682 19406 47684 19458
rect 47628 19346 47684 19406
rect 47628 19294 47630 19346
rect 47682 19294 47684 19346
rect 47628 19282 47684 19294
rect 47628 19124 47684 19134
rect 47628 18562 47684 19068
rect 47628 18510 47630 18562
rect 47682 18510 47684 18562
rect 47628 18498 47684 18510
rect 47516 17266 47572 17276
rect 47404 16882 47460 16894
rect 47404 16830 47406 16882
rect 47458 16830 47460 16882
rect 47404 16772 47460 16830
rect 47404 16706 47460 16716
rect 47516 16660 47572 16670
rect 47292 16098 47460 16100
rect 47292 16046 47294 16098
rect 47346 16046 47460 16098
rect 47292 16044 47460 16046
rect 47292 16034 47348 16044
rect 47180 15988 47236 15998
rect 47068 15986 47236 15988
rect 47068 15934 47182 15986
rect 47234 15934 47236 15986
rect 47068 15932 47236 15934
rect 46956 15810 47012 15820
rect 46956 15652 47012 15662
rect 46956 15538 47012 15596
rect 46956 15486 46958 15538
rect 47010 15486 47012 15538
rect 46956 15474 47012 15486
rect 47180 15540 47236 15932
rect 47404 15652 47460 16044
rect 47404 15586 47460 15596
rect 47180 15484 47348 15540
rect 47180 15316 47236 15354
rect 47180 15250 47236 15260
rect 47068 15202 47124 15214
rect 47068 15150 47070 15202
rect 47122 15150 47124 15202
rect 47068 15148 47124 15150
rect 46956 15092 47124 15148
rect 45836 14028 46116 14084
rect 45724 13970 45780 13982
rect 45724 13918 45726 13970
rect 45778 13918 45780 13970
rect 45724 13524 45780 13918
rect 45724 13458 45780 13468
rect 45500 13022 45502 13074
rect 45554 13022 45556 13074
rect 45500 13010 45556 13022
rect 45948 13076 46004 13086
rect 45948 12982 46004 13020
rect 45836 12852 45892 12862
rect 45388 12796 45668 12852
rect 44940 11620 44996 11900
rect 45164 11844 45220 12460
rect 45276 12628 45332 12638
rect 45276 12292 45332 12572
rect 45500 12292 45556 12302
rect 45276 12290 45556 12292
rect 45276 12238 45502 12290
rect 45554 12238 45556 12290
rect 45276 12236 45556 12238
rect 45500 12226 45556 12236
rect 45612 12068 45668 12796
rect 45164 11778 45220 11788
rect 45500 12012 45668 12068
rect 45724 12178 45780 12190
rect 45724 12126 45726 12178
rect 45778 12126 45780 12178
rect 44940 11554 44996 11564
rect 45052 11732 45108 11742
rect 45052 10834 45108 11676
rect 45052 10782 45054 10834
rect 45106 10782 45108 10834
rect 45052 10770 45108 10782
rect 45276 11284 45332 11294
rect 44940 10724 44996 10734
rect 44828 10722 44996 10724
rect 44828 10670 44942 10722
rect 44994 10670 44996 10722
rect 44828 10668 44996 10670
rect 44940 10658 44996 10668
rect 45052 10386 45108 10398
rect 45052 10334 45054 10386
rect 45106 10334 45108 10386
rect 44492 10276 44548 10286
rect 43820 9714 43876 9726
rect 43820 9662 43822 9714
rect 43874 9662 43876 9714
rect 43820 9268 43876 9662
rect 43820 8932 43876 9212
rect 43820 8866 43876 8876
rect 44492 9602 44548 10220
rect 44716 10052 44772 10062
rect 44716 9958 44772 9996
rect 44492 9550 44494 9602
rect 44546 9550 44548 9602
rect 43484 7586 43540 8204
rect 43484 7534 43486 7586
rect 43538 7534 43540 7586
rect 43484 7522 43540 7534
rect 43596 8204 43764 8260
rect 44044 8260 44100 8270
rect 43596 7364 43652 8204
rect 44044 8166 44100 8204
rect 44380 8034 44436 8046
rect 44380 7982 44382 8034
rect 44434 7982 44436 8034
rect 44380 7924 44436 7982
rect 44380 7858 44436 7868
rect 43820 7812 43876 7822
rect 43820 7698 43876 7756
rect 43820 7646 43822 7698
rect 43874 7646 43876 7698
rect 43820 7634 43876 7646
rect 44380 7700 44436 7710
rect 44380 7606 44436 7644
rect 43036 6466 43316 6468
rect 43036 6414 43038 6466
rect 43090 6414 43316 6466
rect 43036 6412 43316 6414
rect 43484 7308 43652 7364
rect 43484 6468 43540 7308
rect 43596 6692 43652 6702
rect 43596 6598 43652 6636
rect 44492 6692 44548 9550
rect 44604 9602 44660 9614
rect 44604 9550 44606 9602
rect 44658 9550 44660 9602
rect 44604 9044 44660 9550
rect 44716 9044 44772 9054
rect 44604 9042 44772 9044
rect 44604 8990 44718 9042
rect 44770 8990 44772 9042
rect 44604 8988 44772 8990
rect 44716 8978 44772 8988
rect 45052 9042 45108 10334
rect 45052 8990 45054 9042
rect 45106 8990 45108 9042
rect 45052 8978 45108 8990
rect 45164 9940 45220 9950
rect 45052 7700 45108 7710
rect 45164 7700 45220 9884
rect 45052 7698 45220 7700
rect 45052 7646 45054 7698
rect 45106 7646 45220 7698
rect 45052 7644 45220 7646
rect 45052 7634 45108 7644
rect 44492 6626 44548 6636
rect 44604 7028 44660 7038
rect 43484 6412 43652 6468
rect 42588 6356 42644 6366
rect 42588 6132 42644 6300
rect 42700 6132 42756 6142
rect 42588 6130 42756 6132
rect 42588 6078 42702 6130
rect 42754 6078 42756 6130
rect 42588 6076 42756 6078
rect 42700 6066 42756 6076
rect 42812 6020 42868 6030
rect 42812 5926 42868 5964
rect 43036 5796 43092 6412
rect 43036 5730 43092 5740
rect 43484 6018 43540 6030
rect 43484 5966 43486 6018
rect 43538 5966 43540 6018
rect 43484 5796 43540 5966
rect 43484 5730 43540 5740
rect 42588 5682 42644 5694
rect 42588 5630 42590 5682
rect 42642 5630 42644 5682
rect 41916 5124 41972 5134
rect 41916 5030 41972 5068
rect 42588 5124 42644 5630
rect 42588 5058 42644 5068
rect 43596 5012 43652 6412
rect 44044 6466 44100 6478
rect 44044 6414 44046 6466
rect 44098 6414 44100 6466
rect 44044 6356 44100 6414
rect 43932 6300 44044 6356
rect 43820 6020 43876 6030
rect 43820 5926 43876 5964
rect 43820 5236 43876 5246
rect 43932 5236 43988 6300
rect 44044 6290 44100 6300
rect 44380 6466 44436 6478
rect 44380 6414 44382 6466
rect 44434 6414 44436 6466
rect 44380 6244 44436 6414
rect 44380 6178 44436 6188
rect 44492 6132 44548 6142
rect 44604 6132 44660 6972
rect 45276 6692 45332 11228
rect 45388 11172 45444 11182
rect 45388 9938 45444 11116
rect 45500 10500 45556 12012
rect 45724 11732 45780 12126
rect 45724 11666 45780 11676
rect 45836 11844 45892 12796
rect 45612 11396 45668 11406
rect 45836 11396 45892 11788
rect 45612 11394 45892 11396
rect 45612 11342 45614 11394
rect 45666 11342 45892 11394
rect 45612 11340 45892 11342
rect 45948 12068 46004 12078
rect 45948 11394 46004 12012
rect 45948 11342 45950 11394
rect 46002 11342 46004 11394
rect 45612 11330 45668 11340
rect 45948 11330 46004 11342
rect 45724 11170 45780 11182
rect 45724 11118 45726 11170
rect 45778 11118 45780 11170
rect 45724 11060 45780 11118
rect 45724 10724 45780 11004
rect 45724 10658 45780 10668
rect 45836 11170 45892 11182
rect 45836 11118 45838 11170
rect 45890 11118 45892 11170
rect 45724 10500 45780 10510
rect 45500 10498 45780 10500
rect 45500 10446 45726 10498
rect 45778 10446 45780 10498
rect 45500 10444 45780 10446
rect 45388 9886 45390 9938
rect 45442 9886 45444 9938
rect 45388 9874 45444 9886
rect 45724 9156 45780 10444
rect 45724 9090 45780 9100
rect 45836 10052 45892 11118
rect 46060 11172 46116 14028
rect 46172 13636 46228 14252
rect 46172 13570 46228 13580
rect 46396 14252 46564 14308
rect 46732 14308 46788 14318
rect 46172 12292 46228 12302
rect 46172 11394 46228 12236
rect 46172 11342 46174 11394
rect 46226 11342 46228 11394
rect 46172 11330 46228 11342
rect 46284 11844 46340 11854
rect 46060 11116 46228 11172
rect 46060 10836 46116 10846
rect 46060 10742 46116 10780
rect 45612 8932 45668 8942
rect 45388 8930 45668 8932
rect 45388 8878 45614 8930
rect 45666 8878 45668 8930
rect 45388 8876 45668 8878
rect 45388 7252 45444 8876
rect 45612 8866 45668 8876
rect 45500 8260 45556 8270
rect 45500 8258 45780 8260
rect 45500 8206 45502 8258
rect 45554 8206 45780 8258
rect 45500 8204 45780 8206
rect 45500 8194 45556 8204
rect 45612 8034 45668 8046
rect 45612 7982 45614 8034
rect 45666 7982 45668 8034
rect 45500 7812 45556 7822
rect 45500 7586 45556 7756
rect 45500 7534 45502 7586
rect 45554 7534 45556 7586
rect 45500 7522 45556 7534
rect 45388 7196 45556 7252
rect 45388 6692 45444 6702
rect 45276 6690 45444 6692
rect 45276 6638 45390 6690
rect 45442 6638 45444 6690
rect 45276 6636 45444 6638
rect 45388 6468 45444 6636
rect 45388 6402 45444 6412
rect 44492 6130 44660 6132
rect 44492 6078 44494 6130
rect 44546 6078 44660 6130
rect 44492 6076 44660 6078
rect 45276 6356 45332 6366
rect 45276 6130 45332 6300
rect 45276 6078 45278 6130
rect 45330 6078 45332 6130
rect 44492 6066 44548 6076
rect 44380 6020 44436 6030
rect 44380 5926 44436 5964
rect 43820 5234 43988 5236
rect 43820 5182 43822 5234
rect 43874 5182 43988 5234
rect 43820 5180 43988 5182
rect 45276 5236 45332 6078
rect 45388 6132 45444 6142
rect 45388 6038 45444 6076
rect 45500 6018 45556 7196
rect 45612 7140 45668 7982
rect 45724 8036 45780 8204
rect 45836 8258 45892 9996
rect 45948 10724 46004 10734
rect 45948 9268 46004 10668
rect 46172 9938 46228 11116
rect 46172 9886 46174 9938
rect 46226 9886 46228 9938
rect 46172 9874 46228 9886
rect 46284 9380 46340 11788
rect 46396 11394 46452 14252
rect 46732 14214 46788 14252
rect 46508 14084 46564 14094
rect 46508 13748 46564 14028
rect 46844 13970 46900 13982
rect 46844 13918 46846 13970
rect 46898 13918 46900 13970
rect 46732 13860 46788 13870
rect 46732 13766 46788 13804
rect 46508 13654 46564 13692
rect 46732 13524 46788 13534
rect 46508 12964 46564 12974
rect 46508 12870 46564 12908
rect 46732 12962 46788 13468
rect 46844 13076 46900 13918
rect 46956 13860 47012 15092
rect 47068 14420 47124 14430
rect 47068 14326 47124 14364
rect 47180 14308 47236 14318
rect 46956 13794 47012 13804
rect 47068 14196 47124 14206
rect 47068 13522 47124 14140
rect 47180 13746 47236 14252
rect 47180 13694 47182 13746
rect 47234 13694 47236 13746
rect 47180 13682 47236 13694
rect 47068 13470 47070 13522
rect 47122 13470 47124 13522
rect 47068 13458 47124 13470
rect 46844 13020 47236 13076
rect 46732 12910 46734 12962
rect 46786 12910 46788 12962
rect 46732 12898 46788 12910
rect 46620 12738 46676 12750
rect 46620 12686 46622 12738
rect 46674 12686 46676 12738
rect 46396 11342 46398 11394
rect 46450 11342 46452 11394
rect 46396 11330 46452 11342
rect 46508 12178 46564 12190
rect 46508 12126 46510 12178
rect 46562 12126 46564 12178
rect 46508 12068 46564 12126
rect 46508 9940 46564 12012
rect 46620 10948 46676 12686
rect 46956 12740 47012 12750
rect 46956 12738 47124 12740
rect 46956 12686 46958 12738
rect 47010 12686 47124 12738
rect 46956 12684 47124 12686
rect 46956 12674 47012 12684
rect 47068 12292 47124 12684
rect 47180 12402 47236 13020
rect 47292 12964 47348 15484
rect 47516 15428 47572 16604
rect 47516 15314 47572 15372
rect 47516 15262 47518 15314
rect 47570 15262 47572 15314
rect 47516 15250 47572 15262
rect 47404 15204 47460 15214
rect 47404 13972 47460 15148
rect 47740 15092 47796 20524
rect 47852 17220 47908 20636
rect 48188 20020 48244 20030
rect 48188 19926 48244 19964
rect 48412 19796 48468 19806
rect 48076 19572 48132 19582
rect 48076 19346 48132 19516
rect 48076 19294 48078 19346
rect 48130 19294 48132 19346
rect 48076 19282 48132 19294
rect 48412 19348 48468 19740
rect 48524 19572 48580 22316
rect 48636 22306 48692 22316
rect 48860 22258 48916 22270
rect 48860 22206 48862 22258
rect 48914 22206 48916 22258
rect 48636 22146 48692 22158
rect 48636 22094 48638 22146
rect 48690 22094 48692 22146
rect 48636 21028 48692 22094
rect 48860 21812 48916 22206
rect 49084 22258 49140 22428
rect 49420 22372 49476 25228
rect 49644 24722 49700 25678
rect 49980 25060 50036 27020
rect 50204 27010 50260 27020
rect 50428 26964 50484 26974
rect 50988 26908 51044 30156
rect 51100 29540 51156 31500
rect 51212 31490 51268 31500
rect 51324 31106 51380 31118
rect 51324 31054 51326 31106
rect 51378 31054 51380 31106
rect 51324 30212 51380 31054
rect 51660 31106 51716 32620
rect 51996 32562 52052 32574
rect 51996 32510 51998 32562
rect 52050 32510 52052 32562
rect 51996 32452 52052 32510
rect 51996 32386 52052 32396
rect 51660 31054 51662 31106
rect 51714 31054 51716 31106
rect 51660 31042 51716 31054
rect 52108 31554 52164 31566
rect 52108 31502 52110 31554
rect 52162 31502 52164 31554
rect 52108 30884 52164 31502
rect 52332 31556 52388 33628
rect 52668 32676 52724 32686
rect 52556 32338 52612 32350
rect 52556 32286 52558 32338
rect 52610 32286 52612 32338
rect 52444 31780 52500 31790
rect 52556 31780 52612 32286
rect 52500 31724 52612 31780
rect 52444 31648 52500 31724
rect 52332 31500 52500 31556
rect 52108 30818 52164 30828
rect 52332 30772 52388 30782
rect 52332 30678 52388 30716
rect 51324 30146 51380 30156
rect 51436 30324 51492 30334
rect 51324 29986 51380 29998
rect 51324 29934 51326 29986
rect 51378 29934 51380 29986
rect 51212 29876 51268 29886
rect 51324 29876 51380 29934
rect 51268 29820 51380 29876
rect 51212 29810 51268 29820
rect 51436 29764 51492 30268
rect 51660 29988 51716 29998
rect 51324 29708 51492 29764
rect 51548 29986 51716 29988
rect 51548 29934 51662 29986
rect 51714 29934 51716 29986
rect 51548 29932 51716 29934
rect 51100 29474 51156 29484
rect 51212 29652 51268 29662
rect 51212 29538 51268 29596
rect 51212 29486 51214 29538
rect 51266 29486 51268 29538
rect 51212 28868 51268 29486
rect 51324 29314 51380 29708
rect 51324 29262 51326 29314
rect 51378 29262 51380 29314
rect 51324 29092 51380 29262
rect 51324 29026 51380 29036
rect 51436 29426 51492 29438
rect 51436 29374 51438 29426
rect 51490 29374 51492 29426
rect 51212 28802 51268 28812
rect 51436 28532 51492 29374
rect 51548 29316 51604 29932
rect 51660 29922 51716 29932
rect 52220 29986 52276 29998
rect 52220 29934 52222 29986
rect 52274 29934 52276 29986
rect 51548 29250 51604 29260
rect 51772 29876 51828 29886
rect 51772 29426 51828 29820
rect 51772 29374 51774 29426
rect 51826 29374 51828 29426
rect 51772 29316 51828 29374
rect 51772 29250 51828 29260
rect 51884 29540 51940 29550
rect 51884 28644 51940 29484
rect 52108 29314 52164 29326
rect 52108 29262 52110 29314
rect 52162 29262 52164 29314
rect 52108 29204 52164 29262
rect 52108 29138 52164 29148
rect 51660 28532 51716 28542
rect 51436 28476 51660 28532
rect 51660 28438 51716 28476
rect 51324 28420 51380 28430
rect 51324 28418 51604 28420
rect 51324 28366 51326 28418
rect 51378 28366 51604 28418
rect 51324 28364 51604 28366
rect 51324 28354 51380 28364
rect 50428 26870 50484 26908
rect 50204 26850 50260 26862
rect 50204 26798 50206 26850
rect 50258 26798 50260 26850
rect 50204 26180 50260 26798
rect 50876 26852 51044 26908
rect 51212 28084 51268 28094
rect 51212 27076 51268 28028
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50764 26292 50820 26302
rect 50876 26292 50932 26852
rect 50764 26290 50932 26292
rect 50764 26238 50766 26290
rect 50818 26238 50932 26290
rect 50764 26236 50932 26238
rect 50764 26226 50820 26236
rect 50204 26114 50260 26124
rect 50428 26066 50484 26078
rect 50428 26014 50430 26066
rect 50482 26014 50484 26066
rect 50428 25394 50484 26014
rect 50876 25730 50932 26236
rect 50988 26180 51044 26190
rect 50988 26086 51044 26124
rect 50876 25678 50878 25730
rect 50930 25678 50932 25730
rect 50876 25666 50932 25678
rect 50428 25342 50430 25394
rect 50482 25342 50484 25394
rect 50092 25284 50148 25294
rect 50092 25190 50148 25228
rect 49980 25004 50148 25060
rect 49980 24836 50036 24846
rect 49980 24742 50036 24780
rect 49644 24670 49646 24722
rect 49698 24670 49700 24722
rect 49644 24658 49700 24670
rect 49756 24722 49812 24734
rect 49756 24670 49758 24722
rect 49810 24670 49812 24722
rect 49644 24500 49700 24510
rect 49644 24406 49700 24444
rect 49756 24164 49812 24670
rect 49756 24098 49812 24108
rect 49868 24052 49924 24062
rect 49868 23938 49924 23996
rect 49868 23886 49870 23938
rect 49922 23886 49924 23938
rect 49868 23874 49924 23886
rect 49532 23716 49588 23726
rect 49532 23714 49700 23716
rect 49532 23662 49534 23714
rect 49586 23662 49700 23714
rect 49532 23660 49700 23662
rect 49532 23650 49588 23660
rect 49644 23604 49700 23660
rect 49644 23548 49924 23604
rect 49532 23492 49588 23502
rect 49532 23154 49588 23436
rect 49532 23102 49534 23154
rect 49586 23102 49588 23154
rect 49532 22596 49588 23102
rect 49756 23154 49812 23166
rect 49756 23102 49758 23154
rect 49810 23102 49812 23154
rect 49532 22530 49588 22540
rect 49644 23042 49700 23054
rect 49644 22990 49646 23042
rect 49698 22990 49700 23042
rect 49420 22306 49476 22316
rect 49084 22206 49086 22258
rect 49138 22206 49140 22258
rect 49084 22194 49140 22206
rect 49532 22148 49588 22158
rect 49532 22054 49588 22092
rect 49644 22036 49700 22990
rect 49756 22932 49812 23102
rect 49756 22866 49812 22876
rect 49868 23044 49924 23548
rect 50092 23380 50148 25004
rect 50204 24724 50260 24734
rect 50316 24724 50372 24734
rect 50204 24722 50316 24724
rect 50204 24670 50206 24722
rect 50258 24670 50316 24722
rect 50204 24668 50316 24670
rect 50204 24658 50260 24668
rect 49868 22484 49924 22988
rect 49868 22418 49924 22428
rect 49980 23324 50148 23380
rect 50204 24500 50260 24510
rect 49980 22372 50036 23324
rect 50092 23154 50148 23166
rect 50092 23102 50094 23154
rect 50146 23102 50148 23154
rect 50092 23044 50148 23102
rect 50092 22978 50148 22988
rect 49980 22316 50148 22372
rect 49980 22148 50036 22158
rect 49980 22054 50036 22092
rect 49756 22036 49812 22046
rect 49644 21980 49756 22036
rect 49756 21970 49812 21980
rect 48972 21812 49028 21822
rect 48860 21756 48972 21812
rect 48972 21746 49028 21756
rect 49420 21812 49476 21822
rect 49644 21812 49700 21822
rect 49476 21810 49700 21812
rect 49476 21758 49646 21810
rect 49698 21758 49700 21810
rect 49476 21756 49700 21758
rect 49420 21746 49476 21756
rect 49644 21746 49700 21756
rect 49756 21812 49812 21822
rect 50092 21812 50148 22316
rect 48748 21588 48804 21598
rect 48748 21494 48804 21532
rect 49532 21588 49588 21598
rect 49588 21532 49700 21588
rect 49532 21456 49588 21532
rect 48636 20962 48692 20972
rect 49532 21028 49588 21038
rect 49532 20934 49588 20972
rect 49196 20804 49252 20814
rect 48636 20690 48692 20702
rect 48636 20638 48638 20690
rect 48690 20638 48692 20690
rect 48636 20244 48692 20638
rect 48860 20690 48916 20702
rect 48860 20638 48862 20690
rect 48914 20638 48916 20690
rect 48636 20178 48692 20188
rect 48748 20578 48804 20590
rect 48748 20526 48750 20578
rect 48802 20526 48804 20578
rect 48636 20020 48692 20030
rect 48636 19926 48692 19964
rect 48524 19506 48580 19516
rect 48524 19348 48580 19358
rect 48412 19346 48580 19348
rect 48412 19294 48526 19346
rect 48578 19294 48580 19346
rect 48412 19292 48580 19294
rect 48524 19282 48580 19292
rect 48188 18788 48244 18798
rect 48188 18674 48244 18732
rect 48188 18622 48190 18674
rect 48242 18622 48244 18674
rect 48188 18610 48244 18622
rect 48412 18676 48468 18686
rect 48412 18582 48468 18620
rect 48300 18564 48356 18574
rect 48300 18470 48356 18508
rect 48300 18228 48356 18238
rect 48300 17778 48356 18172
rect 48300 17726 48302 17778
rect 48354 17726 48356 17778
rect 48300 17714 48356 17726
rect 48300 17332 48356 17342
rect 47852 17164 48244 17220
rect 48188 17106 48244 17164
rect 48188 17054 48190 17106
rect 48242 17054 48244 17106
rect 47852 16996 47908 17006
rect 47852 16210 47908 16940
rect 47852 16158 47854 16210
rect 47906 16158 47908 16210
rect 47852 15876 47908 16158
rect 47852 15810 47908 15820
rect 47964 16772 48020 16782
rect 47964 15652 48020 16716
rect 48188 16660 48244 17054
rect 48300 16772 48356 17276
rect 48748 17220 48804 20526
rect 48860 20468 48916 20638
rect 49084 20580 49140 20590
rect 49084 20486 49140 20524
rect 48860 19796 48916 20412
rect 48860 19730 48916 19740
rect 48972 19908 49028 19918
rect 48972 19346 49028 19852
rect 48972 19294 48974 19346
rect 49026 19294 49028 19346
rect 48972 19282 49028 19294
rect 49196 19012 49252 20748
rect 49420 20804 49476 20814
rect 49420 20710 49476 20748
rect 49644 20468 49700 21532
rect 49756 21586 49812 21756
rect 49756 21534 49758 21586
rect 49810 21534 49812 21586
rect 49756 21028 49812 21534
rect 49756 20962 49812 20972
rect 49980 21756 50148 21812
rect 49644 20402 49700 20412
rect 49420 19908 49476 19918
rect 49420 19906 49588 19908
rect 49420 19854 49422 19906
rect 49474 19854 49588 19906
rect 49420 19852 49588 19854
rect 49420 19842 49476 19852
rect 49420 19348 49476 19358
rect 49420 19254 49476 19292
rect 49196 18946 49252 18956
rect 48860 18450 48916 18462
rect 48860 18398 48862 18450
rect 48914 18398 48916 18450
rect 48860 18340 48916 18398
rect 48860 18274 48916 18284
rect 48972 18452 49028 18462
rect 48748 17154 48804 17164
rect 48860 17892 48916 17902
rect 48300 16706 48356 16716
rect 48748 16772 48804 16782
rect 48748 16678 48804 16716
rect 48188 16594 48244 16604
rect 48412 16324 48468 16334
rect 48300 16100 48356 16110
rect 47740 15026 47796 15036
rect 47852 15596 48020 15652
rect 48076 15652 48132 15662
rect 47404 13636 47460 13916
rect 47740 14530 47796 14542
rect 47740 14478 47742 14530
rect 47794 14478 47796 14530
rect 47740 14420 47796 14478
rect 47740 13972 47796 14364
rect 47740 13906 47796 13916
rect 47404 13570 47460 13580
rect 47292 12908 47684 12964
rect 47516 12738 47572 12750
rect 47516 12686 47518 12738
rect 47570 12686 47572 12738
rect 47516 12516 47572 12686
rect 47516 12450 47572 12460
rect 47180 12350 47182 12402
rect 47234 12350 47236 12402
rect 47180 12338 47236 12350
rect 47068 12226 47124 12236
rect 47404 12178 47460 12190
rect 47404 12126 47406 12178
rect 47458 12126 47460 12178
rect 47292 12068 47348 12078
rect 46844 12066 47348 12068
rect 46844 12014 47294 12066
rect 47346 12014 47348 12066
rect 46844 12012 47348 12014
rect 46844 11732 46900 12012
rect 47292 12002 47348 12012
rect 47404 11844 47460 12126
rect 46844 11666 46900 11676
rect 46956 11788 47460 11844
rect 47516 12068 47572 12078
rect 46956 11618 47012 11788
rect 46956 11566 46958 11618
rect 47010 11566 47012 11618
rect 46956 11554 47012 11566
rect 47404 11618 47460 11630
rect 47404 11566 47406 11618
rect 47458 11566 47460 11618
rect 46620 10882 46676 10892
rect 46732 11394 46788 11406
rect 46732 11342 46734 11394
rect 46786 11342 46788 11394
rect 46508 9808 46564 9884
rect 46732 10498 46788 11342
rect 47180 11396 47236 11406
rect 46732 10446 46734 10498
rect 46786 10446 46788 10498
rect 46284 9324 46564 9380
rect 46060 9268 46116 9278
rect 45948 9266 46116 9268
rect 45948 9214 46062 9266
rect 46114 9214 46116 9266
rect 45948 9212 46116 9214
rect 46060 9202 46116 9212
rect 46508 9266 46564 9324
rect 46508 9214 46510 9266
rect 46562 9214 46564 9266
rect 45836 8206 45838 8258
rect 45890 8206 45892 8258
rect 45836 8194 45892 8206
rect 45724 7980 45892 8036
rect 45724 7588 45780 7598
rect 45724 7494 45780 7532
rect 45612 7074 45668 7084
rect 45836 6244 45892 7980
rect 46396 7924 46452 7934
rect 46172 7474 46228 7486
rect 46172 7422 46174 7474
rect 46226 7422 46228 7474
rect 45948 7362 46004 7374
rect 45948 7310 45950 7362
rect 46002 7310 46004 7362
rect 45948 7028 46004 7310
rect 46172 7364 46228 7422
rect 46172 7298 46228 7308
rect 45948 6972 46228 7028
rect 46172 6690 46228 6972
rect 46172 6638 46174 6690
rect 46226 6638 46228 6690
rect 46172 6626 46228 6638
rect 46060 6580 46116 6590
rect 46060 6486 46116 6524
rect 45948 6244 46004 6254
rect 45836 6188 45948 6244
rect 45948 6130 46004 6188
rect 45948 6078 45950 6130
rect 46002 6078 46004 6130
rect 45948 6066 46004 6078
rect 45500 5966 45502 6018
rect 45554 5966 45556 6018
rect 45500 5954 45556 5966
rect 45388 5236 45444 5246
rect 45276 5234 45444 5236
rect 45276 5182 45390 5234
rect 45442 5182 45444 5234
rect 45276 5180 45444 5182
rect 43820 5170 43876 5180
rect 45388 5170 45444 5180
rect 46396 5234 46452 7868
rect 46508 6130 46564 9214
rect 46732 9044 46788 10446
rect 46732 8978 46788 8988
rect 46844 11282 46900 11294
rect 46844 11230 46846 11282
rect 46898 11230 46900 11282
rect 46844 11172 46900 11230
rect 46844 8484 46900 11116
rect 47180 10834 47236 11340
rect 47180 10782 47182 10834
rect 47234 10782 47236 10834
rect 47180 10770 47236 10782
rect 47404 11170 47460 11566
rect 47404 11118 47406 11170
rect 47458 11118 47460 11170
rect 47292 9604 47348 9614
rect 46844 8418 46900 8428
rect 47068 9602 47348 9604
rect 47068 9550 47294 9602
rect 47346 9550 47348 9602
rect 47068 9548 47348 9550
rect 47068 8372 47124 9548
rect 47292 9538 47348 9548
rect 47404 9604 47460 11118
rect 47404 9538 47460 9548
rect 47516 9826 47572 12012
rect 47628 10836 47684 12908
rect 47852 12178 47908 15596
rect 47964 15202 48020 15214
rect 47964 15150 47966 15202
rect 48018 15150 48020 15202
rect 47964 14756 48020 15150
rect 47964 14306 48020 14700
rect 47964 14254 47966 14306
rect 48018 14254 48020 14306
rect 47964 14196 48020 14254
rect 47964 14130 48020 14140
rect 48076 13188 48132 15596
rect 48300 14644 48356 16044
rect 48412 16098 48468 16268
rect 48524 16324 48580 16334
rect 48524 16322 48692 16324
rect 48524 16270 48526 16322
rect 48578 16270 48692 16322
rect 48524 16268 48692 16270
rect 48524 16258 48580 16268
rect 48412 16046 48414 16098
rect 48466 16046 48468 16098
rect 48412 15764 48468 16046
rect 48524 15988 48580 15998
rect 48524 15894 48580 15932
rect 48412 15708 48580 15764
rect 48412 15428 48468 15438
rect 48412 15334 48468 15372
rect 48412 14644 48468 14654
rect 48300 14642 48468 14644
rect 48300 14590 48414 14642
rect 48466 14590 48468 14642
rect 48300 14588 48468 14590
rect 48412 14578 48468 14588
rect 48188 14308 48244 14318
rect 48188 13970 48244 14252
rect 48188 13918 48190 13970
rect 48242 13918 48244 13970
rect 48188 13906 48244 13918
rect 48412 13748 48468 13758
rect 48412 13654 48468 13692
rect 47852 12126 47854 12178
rect 47906 12126 47908 12178
rect 47852 11396 47908 12126
rect 47852 11330 47908 11340
rect 47964 13132 48132 13188
rect 48188 13636 48244 13646
rect 47852 11170 47908 11182
rect 47852 11118 47854 11170
rect 47906 11118 47908 11170
rect 47740 10836 47796 10846
rect 47628 10834 47796 10836
rect 47628 10782 47742 10834
rect 47794 10782 47796 10834
rect 47628 10780 47796 10782
rect 47740 10770 47796 10780
rect 47852 10052 47908 11118
rect 47964 10836 48020 13132
rect 48076 12964 48132 12974
rect 48076 11060 48132 12908
rect 48188 12852 48244 13580
rect 48300 13634 48356 13646
rect 48300 13582 48302 13634
rect 48354 13582 48356 13634
rect 48300 13524 48356 13582
rect 48300 12964 48356 13468
rect 48300 12908 48468 12964
rect 48188 12796 48356 12852
rect 48188 12068 48244 12078
rect 48188 11974 48244 12012
rect 48300 11844 48356 12796
rect 48188 11788 48356 11844
rect 48188 11618 48244 11788
rect 48188 11566 48190 11618
rect 48242 11566 48244 11618
rect 48188 11554 48244 11566
rect 48300 11508 48356 11518
rect 48300 11414 48356 11452
rect 48412 11284 48468 12908
rect 48300 11228 48468 11284
rect 48076 11004 48244 11060
rect 48076 10836 48132 10846
rect 47964 10834 48132 10836
rect 47964 10782 48078 10834
rect 48130 10782 48132 10834
rect 47964 10780 48132 10782
rect 47852 9986 47908 9996
rect 48076 10050 48132 10780
rect 48076 9998 48078 10050
rect 48130 9998 48132 10050
rect 48076 9986 48132 9998
rect 48188 9828 48244 11004
rect 47516 9774 47518 9826
rect 47570 9774 47572 9826
rect 47292 9268 47348 9278
rect 47292 9174 47348 9212
rect 47516 8932 47572 9774
rect 47740 9772 48244 9828
rect 48300 9828 48356 11228
rect 48524 10836 48580 15708
rect 48636 12962 48692 16268
rect 48636 12910 48638 12962
rect 48690 12910 48692 12962
rect 48636 12898 48692 12910
rect 48748 15652 48804 15662
rect 48748 12402 48804 15596
rect 48860 14756 48916 17836
rect 48972 17220 49028 18396
rect 48972 16100 49028 17164
rect 49420 17108 49476 17118
rect 49084 16100 49140 16110
rect 48972 16098 49140 16100
rect 48972 16046 49086 16098
rect 49138 16046 49140 16098
rect 48972 16044 49140 16046
rect 49084 16034 49140 16044
rect 49084 15652 49140 15662
rect 48860 14642 48916 14700
rect 48860 14590 48862 14642
rect 48914 14590 48916 14642
rect 48860 14578 48916 14590
rect 48972 14980 49028 14990
rect 48972 14644 49028 14924
rect 48972 14578 49028 14588
rect 48972 14196 49028 14206
rect 48748 12350 48750 12402
rect 48802 12350 48804 12402
rect 48748 11508 48804 12350
rect 48748 11442 48804 11452
rect 48860 13860 48916 13870
rect 48860 12850 48916 13804
rect 48860 12798 48862 12850
rect 48914 12798 48916 12850
rect 48748 11284 48804 11294
rect 48748 11190 48804 11228
rect 48636 10836 48692 10846
rect 48524 10834 48692 10836
rect 48524 10782 48638 10834
rect 48690 10782 48692 10834
rect 48524 10780 48692 10782
rect 48636 10770 48692 10780
rect 48636 10164 48692 10174
rect 48524 10050 48580 10062
rect 48524 9998 48526 10050
rect 48578 9998 48580 10050
rect 48524 9938 48580 9998
rect 48524 9886 48526 9938
rect 48578 9886 48580 9938
rect 48524 9874 48580 9886
rect 48300 9772 48468 9828
rect 47740 9156 47796 9772
rect 48188 9604 48244 9614
rect 48188 9510 48244 9548
rect 47516 8866 47572 8876
rect 47628 9154 47796 9156
rect 47628 9102 47742 9154
rect 47794 9102 47796 9154
rect 47628 9100 47796 9102
rect 47068 8306 47124 8316
rect 47292 8484 47348 8494
rect 46844 8260 46900 8270
rect 46732 8148 46788 8158
rect 46620 7812 46676 7822
rect 46620 7474 46676 7756
rect 46620 7422 46622 7474
rect 46674 7422 46676 7474
rect 46620 7410 46676 7422
rect 46732 7364 46788 8092
rect 46844 7588 46900 8204
rect 46956 8034 47012 8046
rect 46956 7982 46958 8034
rect 47010 7982 47012 8034
rect 46956 7924 47012 7982
rect 46956 7858 47012 7868
rect 47068 8034 47124 8046
rect 47068 7982 47070 8034
rect 47122 7982 47124 8034
rect 46844 7474 46900 7532
rect 47068 7588 47124 7982
rect 47180 8036 47236 8046
rect 47180 7942 47236 7980
rect 47068 7522 47124 7532
rect 46844 7422 46846 7474
rect 46898 7422 46900 7474
rect 46844 7410 46900 7422
rect 46732 7252 46788 7308
rect 47068 7362 47124 7374
rect 47068 7310 47070 7362
rect 47122 7310 47124 7362
rect 47068 7252 47124 7310
rect 46732 7196 47124 7252
rect 46620 6692 46676 6702
rect 46620 6598 46676 6636
rect 46508 6078 46510 6130
rect 46562 6078 46564 6130
rect 46508 6066 46564 6078
rect 46396 5182 46398 5234
rect 46450 5182 46452 5234
rect 46396 5170 46452 5182
rect 46732 5236 46788 7196
rect 47180 6132 47236 6142
rect 47292 6132 47348 8428
rect 47516 7700 47572 7710
rect 47516 7606 47572 7644
rect 47516 7028 47572 7038
rect 47180 6130 47348 6132
rect 47180 6078 47182 6130
rect 47234 6078 47348 6130
rect 47180 6076 47348 6078
rect 47404 6580 47460 6590
rect 47180 6066 47236 6076
rect 47404 5796 47460 6524
rect 46732 5104 46788 5180
rect 46844 5460 46900 5470
rect 43596 4946 43652 4956
rect 46844 4562 46900 5404
rect 46844 4510 46846 4562
rect 46898 4510 46900 4562
rect 46844 4498 46900 4510
rect 47292 4564 47348 4574
rect 47404 4564 47460 5740
rect 47516 5010 47572 6972
rect 47628 6692 47684 9100
rect 47740 9090 47796 9100
rect 47852 9042 47908 9054
rect 47852 8990 47854 9042
rect 47906 8990 47908 9042
rect 47740 8260 47796 8270
rect 47740 8166 47796 8204
rect 47852 8148 47908 8990
rect 47964 9042 48020 9054
rect 47964 8990 47966 9042
rect 48018 8990 48020 9042
rect 47964 8932 48020 8990
rect 48020 8876 48356 8932
rect 47964 8866 48020 8876
rect 48076 8370 48132 8382
rect 48076 8318 48078 8370
rect 48130 8318 48132 8370
rect 48076 8260 48132 8318
rect 48076 8194 48132 8204
rect 47852 8082 47908 8092
rect 47964 8036 48020 8046
rect 47964 8034 48132 8036
rect 47964 7982 47966 8034
rect 48018 7982 48132 8034
rect 47964 7980 48132 7982
rect 47964 7970 48020 7980
rect 47852 7588 47908 7598
rect 47852 7474 47908 7532
rect 47852 7422 47854 7474
rect 47906 7422 47908 7474
rect 47852 7410 47908 7422
rect 47628 5460 47684 6636
rect 47964 7252 48020 7262
rect 47964 6690 48020 7196
rect 48076 7028 48132 7980
rect 48188 7700 48244 7710
rect 48188 7606 48244 7644
rect 48076 6962 48132 6972
rect 47964 6638 47966 6690
rect 48018 6638 48020 6690
rect 47964 6626 48020 6638
rect 48188 6692 48244 6702
rect 48076 6468 48132 6478
rect 47628 5394 47684 5404
rect 47964 6466 48132 6468
rect 47964 6414 48078 6466
rect 48130 6414 48132 6466
rect 47964 6412 48132 6414
rect 47516 4958 47518 5010
rect 47570 4958 47572 5010
rect 47516 4946 47572 4958
rect 47852 5346 47908 5358
rect 47852 5294 47854 5346
rect 47906 5294 47908 5346
rect 47852 5236 47908 5294
rect 47964 5348 48020 6412
rect 48076 6402 48132 6412
rect 48076 6244 48132 6254
rect 48076 6130 48132 6188
rect 48076 6078 48078 6130
rect 48130 6078 48132 6130
rect 48076 6066 48132 6078
rect 48188 6132 48244 6636
rect 48300 6132 48356 8876
rect 48412 8372 48468 9772
rect 48412 8306 48468 8316
rect 48524 9716 48580 9726
rect 48524 8370 48580 9660
rect 48636 9266 48692 10108
rect 48636 9214 48638 9266
rect 48690 9214 48692 9266
rect 48636 9202 48692 9214
rect 48524 8318 48526 8370
rect 48578 8318 48580 8370
rect 48524 8306 48580 8318
rect 48636 8484 48692 8494
rect 48412 7586 48468 7598
rect 48412 7534 48414 7586
rect 48466 7534 48468 7586
rect 48412 6580 48468 7534
rect 48524 7250 48580 7262
rect 48524 7198 48526 7250
rect 48578 7198 48580 7250
rect 48524 6804 48580 7198
rect 48524 6738 48580 6748
rect 48412 6514 48468 6524
rect 48524 6578 48580 6590
rect 48524 6526 48526 6578
rect 48578 6526 48580 6578
rect 48412 6132 48468 6142
rect 48300 6130 48468 6132
rect 48300 6078 48414 6130
rect 48466 6078 48468 6130
rect 48300 6076 48468 6078
rect 48188 6066 48244 6076
rect 47964 5282 48020 5292
rect 48300 5460 48356 5470
rect 47292 4562 47460 4564
rect 47292 4510 47294 4562
rect 47346 4510 47460 4562
rect 47292 4508 47460 4510
rect 47740 4564 47796 4574
rect 47852 4564 47908 5180
rect 48300 5234 48356 5404
rect 48300 5182 48302 5234
rect 48354 5182 48356 5234
rect 48300 5170 48356 5182
rect 48412 5236 48468 6076
rect 48524 6132 48580 6526
rect 48636 6580 48692 8428
rect 48860 7364 48916 12798
rect 48972 8370 49028 14140
rect 49084 10948 49140 15596
rect 49420 15538 49476 17052
rect 49532 16212 49588 19852
rect 49868 19906 49924 19918
rect 49868 19854 49870 19906
rect 49922 19854 49924 19906
rect 49868 19796 49924 19854
rect 49868 19730 49924 19740
rect 49868 19348 49924 19358
rect 49868 19254 49924 19292
rect 49980 19124 50036 21756
rect 50092 21588 50148 21598
rect 50092 21494 50148 21532
rect 50092 20690 50148 20702
rect 50092 20638 50094 20690
rect 50146 20638 50148 20690
rect 50092 20580 50148 20638
rect 50092 20514 50148 20524
rect 49980 18676 50036 19068
rect 49980 18610 50036 18620
rect 49644 18452 49700 18462
rect 49644 18358 49700 18396
rect 49980 18450 50036 18462
rect 49980 18398 49982 18450
rect 50034 18398 50036 18450
rect 49756 18228 49812 18238
rect 49980 18228 50036 18398
rect 49756 18226 49924 18228
rect 49756 18174 49758 18226
rect 49810 18174 49924 18226
rect 49756 18172 49924 18174
rect 49756 18162 49812 18172
rect 49644 18004 49700 18014
rect 49644 17668 49700 17948
rect 49644 17536 49700 17612
rect 49756 17556 49812 17566
rect 49756 17462 49812 17500
rect 49868 16882 49924 18172
rect 49980 18162 50036 18172
rect 50204 16994 50260 24444
rect 50316 21140 50372 24668
rect 50428 23940 50484 25342
rect 50876 25396 50932 25406
rect 50876 25302 50932 25340
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 51212 24948 51268 27020
rect 51548 26908 51604 28364
rect 51772 28084 51828 28094
rect 51772 27990 51828 28028
rect 51324 26850 51380 26862
rect 51324 26798 51326 26850
rect 51378 26798 51380 26850
rect 51324 26404 51380 26798
rect 51436 26852 51604 26908
rect 51660 27858 51716 27870
rect 51660 27806 51662 27858
rect 51714 27806 51716 27858
rect 51660 27074 51716 27806
rect 51884 27858 51940 28588
rect 51884 27806 51886 27858
rect 51938 27806 51940 27858
rect 51884 27794 51940 27806
rect 51996 29092 52052 29102
rect 51660 27022 51662 27074
rect 51714 27022 51716 27074
rect 51660 26908 51716 27022
rect 51884 27188 51940 27198
rect 51660 26852 51828 26908
rect 51436 26404 51492 26852
rect 51772 26404 51828 26852
rect 51436 26348 51716 26404
rect 51324 26338 51380 26348
rect 51548 26180 51604 26190
rect 51436 26178 51604 26180
rect 51436 26126 51550 26178
rect 51602 26126 51604 26178
rect 51436 26124 51604 26126
rect 51324 25844 51380 25854
rect 51324 25618 51380 25788
rect 51436 25730 51492 26124
rect 51548 26114 51604 26124
rect 51436 25678 51438 25730
rect 51490 25678 51492 25730
rect 51436 25666 51492 25678
rect 51548 25844 51604 25854
rect 51324 25566 51326 25618
rect 51378 25566 51380 25618
rect 51324 25554 51380 25566
rect 51548 25508 51604 25788
rect 51548 25442 51604 25452
rect 51660 25396 51716 26348
rect 51772 26338 51828 26348
rect 51772 26068 51828 26078
rect 51772 25974 51828 26012
rect 51772 25620 51828 25630
rect 51884 25620 51940 27132
rect 51772 25618 51940 25620
rect 51772 25566 51774 25618
rect 51826 25566 51940 25618
rect 51772 25564 51940 25566
rect 51772 25554 51828 25564
rect 51772 25396 51828 25406
rect 51660 25340 51772 25396
rect 51660 24948 51716 24958
rect 51212 24892 51604 24948
rect 51100 24836 51156 24846
rect 51100 24834 51268 24836
rect 51100 24782 51102 24834
rect 51154 24782 51268 24834
rect 51100 24780 51268 24782
rect 51100 24770 51156 24780
rect 50876 24724 50932 24734
rect 50876 24722 51044 24724
rect 50876 24670 50878 24722
rect 50930 24670 51044 24722
rect 50876 24668 51044 24670
rect 50876 24658 50932 24668
rect 50764 24052 50820 24062
rect 50764 23958 50820 23996
rect 50988 23940 51044 24668
rect 50428 23884 50596 23940
rect 50428 23716 50484 23726
rect 50540 23716 50596 23884
rect 50988 23846 51044 23884
rect 50540 23660 51156 23716
rect 50428 23622 50484 23660
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50428 23380 50484 23390
rect 50428 22482 50484 23324
rect 50652 23380 50708 23390
rect 50540 23044 50596 23054
rect 50540 22950 50596 22988
rect 50428 22430 50430 22482
rect 50482 22430 50484 22482
rect 50428 22418 50484 22430
rect 50652 22148 50708 23324
rect 50988 23156 51044 23166
rect 50988 23062 51044 23100
rect 50316 21074 50372 21084
rect 50428 22092 50708 22148
rect 50876 22148 50932 22158
rect 50876 22146 51044 22148
rect 50876 22094 50878 22146
rect 50930 22094 51044 22146
rect 50876 22092 51044 22094
rect 50428 21028 50484 22092
rect 50876 22082 50932 22092
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50988 21924 51044 22092
rect 50988 21858 51044 21868
rect 50652 21812 50708 21822
rect 50652 21698 50708 21756
rect 50652 21646 50654 21698
rect 50706 21646 50708 21698
rect 50540 21140 50596 21150
rect 50540 21028 50596 21084
rect 50428 21026 50596 21028
rect 50428 20974 50542 21026
rect 50594 20974 50596 21026
rect 50428 20972 50596 20974
rect 50540 20962 50596 20972
rect 50652 20804 50708 21646
rect 50988 21588 51044 21598
rect 50988 21494 51044 21532
rect 50876 20804 50932 20814
rect 50652 20802 51044 20804
rect 50652 20750 50878 20802
rect 50930 20750 51044 20802
rect 50652 20748 51044 20750
rect 50876 20738 50932 20748
rect 50316 20692 50372 20702
rect 50316 20598 50372 20636
rect 50876 20580 50932 20590
rect 50876 20486 50932 20524
rect 50988 20468 51044 20748
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50988 20402 51044 20412
rect 50556 20346 50820 20356
rect 50764 20132 50820 20142
rect 50764 20038 50820 20076
rect 50876 20132 50932 20142
rect 51100 20132 51156 23660
rect 51212 21588 51268 24780
rect 51548 23044 51604 24892
rect 51660 24052 51716 24892
rect 51772 24946 51828 25340
rect 51772 24894 51774 24946
rect 51826 24894 51828 24946
rect 51772 24882 51828 24894
rect 51996 24948 52052 29036
rect 52108 28644 52164 28654
rect 52108 28550 52164 28588
rect 52220 28532 52276 29934
rect 52220 28466 52276 28476
rect 52332 27748 52388 27758
rect 52332 27654 52388 27692
rect 52332 26850 52388 26862
rect 52332 26798 52334 26850
rect 52386 26798 52388 26850
rect 51996 24882 52052 24892
rect 52108 26066 52164 26078
rect 52108 26014 52110 26066
rect 52162 26014 52164 26066
rect 52108 25396 52164 26014
rect 52332 26068 52388 26798
rect 52332 26002 52388 26012
rect 52332 25620 52388 25630
rect 52332 25526 52388 25564
rect 51884 24724 51940 24734
rect 52108 24724 52164 25340
rect 52332 25284 52388 25294
rect 52332 24946 52388 25228
rect 52332 24894 52334 24946
rect 52386 24894 52388 24946
rect 52332 24882 52388 24894
rect 51884 24722 52052 24724
rect 51884 24670 51886 24722
rect 51938 24670 52052 24722
rect 51884 24668 52052 24670
rect 51884 24658 51940 24668
rect 51772 24500 51828 24510
rect 51772 24406 51828 24444
rect 51660 23986 51716 23996
rect 51772 23828 51828 23838
rect 51660 23156 51716 23166
rect 51660 23062 51716 23100
rect 51324 22148 51380 22158
rect 51324 22146 51492 22148
rect 51324 22094 51326 22146
rect 51378 22094 51492 22146
rect 51324 22092 51492 22094
rect 51324 22082 51380 22092
rect 51436 21700 51492 22092
rect 51436 21634 51492 21644
rect 51212 21532 51380 21588
rect 50876 20130 51156 20132
rect 50876 20078 50878 20130
rect 50930 20078 51156 20130
rect 50876 20076 51156 20078
rect 51324 20132 51380 21532
rect 51436 21476 51492 21486
rect 51436 21382 51492 21420
rect 51436 21026 51492 21038
rect 51436 20974 51438 21026
rect 51490 20974 51492 21026
rect 51436 20914 51492 20974
rect 51436 20862 51438 20914
rect 51490 20862 51492 20914
rect 51436 20850 51492 20862
rect 50876 20066 50932 20076
rect 51324 20066 51380 20076
rect 50540 20018 50596 20030
rect 50540 19966 50542 20018
rect 50594 19966 50596 20018
rect 50540 19684 50596 19966
rect 50540 19618 50596 19628
rect 51212 20018 51268 20030
rect 51212 19966 51214 20018
rect 51266 19966 51268 20018
rect 50540 19460 50596 19470
rect 50540 19234 50596 19404
rect 50540 19182 50542 19234
rect 50594 19182 50596 19234
rect 50540 19170 50596 19182
rect 50876 19460 50932 19470
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50764 18452 50820 18462
rect 50764 18358 50820 18396
rect 50876 17780 50932 19404
rect 51100 19460 51156 19470
rect 51212 19460 51268 19966
rect 51548 20020 51604 22988
rect 51772 23042 51828 23772
rect 51884 23826 51940 23838
rect 51884 23774 51886 23826
rect 51938 23774 51940 23826
rect 51884 23716 51940 23774
rect 51884 23650 51940 23660
rect 51884 23380 51940 23390
rect 51996 23380 52052 24668
rect 52108 24658 52164 24668
rect 52108 24498 52164 24510
rect 52108 24446 52110 24498
rect 52162 24446 52164 24498
rect 52108 23940 52164 24446
rect 52444 24164 52500 31500
rect 52668 30884 52724 32620
rect 52556 30882 52724 30884
rect 52556 30830 52670 30882
rect 52722 30830 52724 30882
rect 52556 30828 52724 30830
rect 52556 30210 52612 30828
rect 52668 30818 52724 30828
rect 52556 30158 52558 30210
rect 52610 30158 52612 30210
rect 52556 30146 52612 30158
rect 52556 29428 52612 29438
rect 52556 29314 52612 29372
rect 52780 29428 52836 35756
rect 52892 34692 52948 52780
rect 52892 34626 52948 34636
rect 53900 32564 53956 32574
rect 53228 32452 53284 32462
rect 53676 32452 53732 32462
rect 53228 32450 53732 32452
rect 53228 32398 53230 32450
rect 53282 32398 53678 32450
rect 53730 32398 53732 32450
rect 53228 32396 53732 32398
rect 53228 32386 53284 32396
rect 53340 31554 53396 32396
rect 53676 32386 53732 32396
rect 53900 32004 53956 32508
rect 54236 32116 54292 55020
rect 54348 55010 54404 55020
rect 54908 52164 54964 52174
rect 54908 52070 54964 52108
rect 56028 52162 56084 52174
rect 56028 52110 56030 52162
rect 56082 52110 56084 52162
rect 56028 51828 56084 52110
rect 56028 51762 56084 51772
rect 58156 48916 58212 48926
rect 56140 46674 56196 46686
rect 56140 46622 56142 46674
rect 56194 46622 56196 46674
rect 55356 46562 55412 46574
rect 55356 46510 55358 46562
rect 55410 46510 55412 46562
rect 55356 46452 55412 46510
rect 55356 46386 55412 46396
rect 56140 45780 56196 46622
rect 56140 45714 56196 45724
rect 56700 45892 56756 45902
rect 56700 45668 56756 45836
rect 57372 45892 57428 45902
rect 57372 45798 57428 45836
rect 57148 45780 57204 45790
rect 57148 45686 57204 45724
rect 56588 45666 56756 45668
rect 56588 45614 56702 45666
rect 56754 45614 56756 45666
rect 56588 45612 56756 45614
rect 55356 41298 55412 41310
rect 55356 41246 55358 41298
rect 55410 41246 55412 41298
rect 55356 40404 55412 41246
rect 55356 40338 55412 40348
rect 56140 41186 56196 41198
rect 56140 41134 56142 41186
rect 56194 41134 56196 41186
rect 56140 39508 56196 41134
rect 56140 39442 56196 39452
rect 54348 35924 54404 35934
rect 54348 35830 54404 35868
rect 54908 35924 54964 35934
rect 54908 35698 54964 35868
rect 54908 35646 54910 35698
rect 54962 35646 54964 35698
rect 54908 35634 54964 35646
rect 56028 35586 56084 35598
rect 56028 35534 56030 35586
rect 56082 35534 56084 35586
rect 56028 35028 56084 35534
rect 56028 34962 56084 34972
rect 56588 32788 56644 45612
rect 56700 45602 56756 45612
rect 56588 32722 56644 32732
rect 56700 39620 56756 39630
rect 56700 39394 56756 39564
rect 57372 39620 57428 39630
rect 57372 39526 57428 39564
rect 57148 39508 57204 39518
rect 57148 39414 57204 39452
rect 56700 39342 56702 39394
rect 56754 39342 56756 39394
rect 54236 32050 54292 32060
rect 55020 32450 55076 32462
rect 55916 32452 55972 32462
rect 55020 32398 55022 32450
rect 55074 32398 55076 32450
rect 53900 31890 53956 31948
rect 53900 31838 53902 31890
rect 53954 31838 53956 31890
rect 53900 31826 53956 31838
rect 54684 32004 54740 32014
rect 54684 31778 54740 31948
rect 55020 32004 55076 32398
rect 55804 32450 55972 32452
rect 55804 32398 55918 32450
rect 55970 32398 55972 32450
rect 55804 32396 55972 32398
rect 55020 31938 55076 31948
rect 55356 32004 55412 32014
rect 54684 31726 54686 31778
rect 54738 31726 54740 31778
rect 54684 31714 54740 31726
rect 55356 31778 55412 31948
rect 55356 31726 55358 31778
rect 55410 31726 55412 31778
rect 55356 31714 55412 31726
rect 53340 31502 53342 31554
rect 53394 31502 53396 31554
rect 53116 30994 53172 31006
rect 53116 30942 53118 30994
rect 53170 30942 53172 30994
rect 52780 29362 52836 29372
rect 52892 30884 52948 30894
rect 52556 29262 52558 29314
rect 52610 29262 52612 29314
rect 52556 29202 52612 29262
rect 52556 29150 52558 29202
rect 52610 29150 52612 29202
rect 52556 29138 52612 29150
rect 52668 29316 52724 29326
rect 52556 28756 52612 28766
rect 52668 28756 52724 29260
rect 52556 28754 52724 28756
rect 52556 28702 52558 28754
rect 52610 28702 52724 28754
rect 52556 28700 52724 28702
rect 52556 28690 52612 28700
rect 52668 27076 52724 27086
rect 52668 26982 52724 27020
rect 52892 26908 52948 30828
rect 53116 30324 53172 30942
rect 53340 30884 53396 31502
rect 54460 31554 54516 31566
rect 54460 31502 54462 31554
rect 54514 31502 54516 31554
rect 53340 30818 53396 30828
rect 53788 30884 53844 30894
rect 54348 30884 54404 30894
rect 53788 30790 53844 30828
rect 54012 30882 54404 30884
rect 54012 30830 54350 30882
rect 54402 30830 54404 30882
rect 54012 30828 54404 30830
rect 53900 30770 53956 30782
rect 53900 30718 53902 30770
rect 53954 30718 53956 30770
rect 53116 30258 53172 30268
rect 53788 30324 53844 30334
rect 53788 30210 53844 30268
rect 53788 30158 53790 30210
rect 53842 30158 53844 30210
rect 53788 30146 53844 30158
rect 53452 29986 53508 29998
rect 53452 29934 53454 29986
rect 53506 29934 53508 29986
rect 53452 29652 53508 29934
rect 53508 29596 53732 29652
rect 53452 29586 53508 29596
rect 53564 29428 53620 29438
rect 53564 29334 53620 29372
rect 53004 29316 53060 29326
rect 53004 29222 53060 29260
rect 53676 28642 53732 29596
rect 53900 29204 53956 30718
rect 53676 28590 53678 28642
rect 53730 28590 53732 28642
rect 53676 28578 53732 28590
rect 53788 29202 53956 29204
rect 53788 29150 53902 29202
rect 53954 29150 53956 29202
rect 53788 29148 53956 29150
rect 53452 28532 53508 28542
rect 53452 28438 53508 28476
rect 53564 28418 53620 28430
rect 53564 28366 53566 28418
rect 53618 28366 53620 28418
rect 53004 27970 53060 27982
rect 53004 27918 53006 27970
rect 53058 27918 53060 27970
rect 53004 27636 53060 27918
rect 53004 27570 53060 27580
rect 53228 27858 53284 27870
rect 53228 27806 53230 27858
rect 53282 27806 53284 27858
rect 53228 27076 53284 27806
rect 53564 27636 53620 28366
rect 53676 27972 53732 27982
rect 53676 27748 53732 27916
rect 53788 27860 53844 29148
rect 53900 29138 53956 29148
rect 54012 28530 54068 30828
rect 54348 30818 54404 30828
rect 54236 30324 54292 30334
rect 54236 29650 54292 30268
rect 54460 30324 54516 31502
rect 55692 31556 55748 31566
rect 55804 31556 55860 32396
rect 55916 32386 55972 32396
rect 56364 32450 56420 32462
rect 56364 32398 56366 32450
rect 56418 32398 56420 32450
rect 56252 31556 56308 31566
rect 55692 31554 55860 31556
rect 55692 31502 55694 31554
rect 55746 31502 55860 31554
rect 55692 31500 55860 31502
rect 55916 31554 56308 31556
rect 55916 31502 56254 31554
rect 56306 31502 56308 31554
rect 55916 31500 56308 31502
rect 54908 31108 54964 31118
rect 54684 31106 54964 31108
rect 54684 31054 54910 31106
rect 54962 31054 54964 31106
rect 54684 31052 54964 31054
rect 54684 30770 54740 31052
rect 54908 31042 54964 31052
rect 55244 30994 55300 31006
rect 55244 30942 55246 30994
rect 55298 30942 55300 30994
rect 55244 30884 55300 30942
rect 55244 30818 55300 30828
rect 55692 30884 55748 31500
rect 55692 30790 55748 30828
rect 54684 30718 54686 30770
rect 54738 30718 54740 30770
rect 54684 30706 54740 30718
rect 55804 30770 55860 30782
rect 55804 30718 55806 30770
rect 55858 30718 55860 30770
rect 54460 30258 54516 30268
rect 54572 30436 54628 30446
rect 54572 29986 54628 30380
rect 55356 30324 55412 30334
rect 54572 29934 54574 29986
rect 54626 29934 54628 29986
rect 54572 29876 54628 29934
rect 54908 29988 54964 29998
rect 54908 29894 54964 29932
rect 54572 29810 54628 29820
rect 54236 29598 54238 29650
rect 54290 29598 54292 29650
rect 54236 29586 54292 29598
rect 54348 29540 54404 29550
rect 54348 29446 54404 29484
rect 54908 29428 54964 29438
rect 54908 29334 54964 29372
rect 54236 29204 54292 29214
rect 54012 28478 54014 28530
rect 54066 28478 54068 28530
rect 54012 28420 54068 28478
rect 54012 28354 54068 28364
rect 54124 29202 54292 29204
rect 54124 29150 54238 29202
rect 54290 29150 54292 29202
rect 54124 29148 54292 29150
rect 53900 28084 53956 28094
rect 53900 27990 53956 28028
rect 53788 27804 54068 27860
rect 53676 27692 53956 27748
rect 53228 27010 53284 27020
rect 53452 27580 53620 27636
rect 53900 27636 53956 27692
rect 52892 26852 53060 26908
rect 52332 24108 52500 24164
rect 52556 26404 52612 26414
rect 52556 25172 52612 26348
rect 52668 26292 52724 26302
rect 52668 26198 52724 26236
rect 52892 25844 52948 25854
rect 52668 25732 52724 25742
rect 52668 25618 52724 25676
rect 52668 25566 52670 25618
rect 52722 25566 52724 25618
rect 52668 25284 52724 25566
rect 52668 25218 52724 25228
rect 52108 23938 52276 23940
rect 52108 23886 52110 23938
rect 52162 23886 52276 23938
rect 52108 23884 52276 23886
rect 52108 23874 52164 23884
rect 52108 23380 52164 23390
rect 51996 23378 52164 23380
rect 51996 23326 52110 23378
rect 52162 23326 52164 23378
rect 51996 23324 52164 23326
rect 51884 23286 51940 23324
rect 52108 23268 52164 23324
rect 52220 23380 52276 23884
rect 52220 23314 52276 23324
rect 52108 23202 52164 23212
rect 51772 22990 51774 23042
rect 51826 22990 51828 23042
rect 51772 22596 51828 22990
rect 51660 22540 51828 22596
rect 51884 23044 51940 23054
rect 51884 22820 51940 22988
rect 51660 21700 51716 22540
rect 51772 22148 51828 22158
rect 51884 22148 51940 22764
rect 51772 22146 51940 22148
rect 51772 22094 51774 22146
rect 51826 22094 51940 22146
rect 51772 22092 51940 22094
rect 51996 22708 52052 22718
rect 51772 22036 51828 22092
rect 51772 21970 51828 21980
rect 51660 21634 51716 21644
rect 51884 21588 51940 21598
rect 51884 21140 51940 21532
rect 51884 21074 51940 21084
rect 51996 21026 52052 22652
rect 51996 20974 51998 21026
rect 52050 20974 52052 21026
rect 51996 20962 52052 20974
rect 52108 22036 52164 22046
rect 52108 20804 52164 21980
rect 52332 21700 52388 24108
rect 52220 21644 52388 21700
rect 52444 23714 52500 23726
rect 52444 23662 52446 23714
rect 52498 23662 52500 23714
rect 52220 20914 52276 21644
rect 52332 21474 52388 21486
rect 52332 21422 52334 21474
rect 52386 21422 52388 21474
rect 52332 21362 52388 21422
rect 52332 21310 52334 21362
rect 52386 21310 52388 21362
rect 52332 21298 52388 21310
rect 52220 20862 52222 20914
rect 52274 20862 52276 20914
rect 52220 20850 52276 20862
rect 52332 21026 52388 21038
rect 52332 20974 52334 21026
rect 52386 20974 52388 21026
rect 51996 20748 52164 20804
rect 51772 20578 51828 20590
rect 51772 20526 51774 20578
rect 51826 20526 51828 20578
rect 51772 20468 51828 20526
rect 51772 20402 51828 20412
rect 51996 20244 52052 20748
rect 51548 19954 51604 19964
rect 51772 20188 52052 20244
rect 52108 20580 52164 20590
rect 51324 19908 51380 19918
rect 51324 19814 51380 19852
rect 51772 19684 51828 20188
rect 52108 20130 52164 20524
rect 52332 20242 52388 20974
rect 52332 20190 52334 20242
rect 52386 20190 52388 20242
rect 52332 20178 52388 20190
rect 52108 20078 52110 20130
rect 52162 20078 52164 20130
rect 52108 20066 52164 20078
rect 51772 19618 51828 19628
rect 51884 20018 51940 20030
rect 51884 19966 51886 20018
rect 51938 19966 51940 20018
rect 51100 19458 51268 19460
rect 51100 19406 51102 19458
rect 51154 19406 51268 19458
rect 51100 19404 51268 19406
rect 51324 19460 51380 19470
rect 50988 19236 51044 19246
rect 50988 19142 51044 19180
rect 50988 18788 51044 18798
rect 50988 18564 51044 18732
rect 50988 18498 51044 18508
rect 50988 18116 51044 18126
rect 50988 17890 51044 18060
rect 50988 17838 50990 17890
rect 51042 17838 51044 17890
rect 50988 17826 51044 17838
rect 50876 17714 50932 17724
rect 50876 17556 50932 17566
rect 50428 17554 50932 17556
rect 50428 17502 50878 17554
rect 50930 17502 50932 17554
rect 50428 17500 50932 17502
rect 50316 17444 50372 17454
rect 50316 17350 50372 17388
rect 50204 16942 50206 16994
rect 50258 16942 50260 16994
rect 50204 16930 50260 16942
rect 49868 16830 49870 16882
rect 49922 16830 49924 16882
rect 49868 16818 49924 16830
rect 49756 16772 49812 16782
rect 49532 16146 49588 16156
rect 49644 16770 49812 16772
rect 49644 16718 49758 16770
rect 49810 16718 49812 16770
rect 49644 16716 49812 16718
rect 49420 15486 49422 15538
rect 49474 15486 49476 15538
rect 49420 15474 49476 15486
rect 49308 14420 49364 14430
rect 49308 14326 49364 14364
rect 49420 13748 49476 13758
rect 49420 13654 49476 13692
rect 49644 12964 49700 16716
rect 49756 16706 49812 16716
rect 49980 16772 50036 16782
rect 49868 16100 49924 16110
rect 49868 16006 49924 16044
rect 49756 15988 49812 15998
rect 49756 15894 49812 15932
rect 49980 13860 50036 16716
rect 50092 16324 50148 16334
rect 50148 16268 50260 16324
rect 50092 16258 50148 16268
rect 50092 15986 50148 15998
rect 50092 15934 50094 15986
rect 50146 15934 50148 15986
rect 50092 15316 50148 15934
rect 50204 15988 50260 16268
rect 50204 15922 50260 15932
rect 50316 16098 50372 16110
rect 50316 16046 50318 16098
rect 50370 16046 50372 16098
rect 50204 15316 50260 15326
rect 50092 15314 50260 15316
rect 50092 15262 50206 15314
rect 50258 15262 50260 15314
rect 50092 15260 50260 15262
rect 50204 15250 50260 15260
rect 50316 14980 50372 16046
rect 50428 15428 50484 17500
rect 50876 17490 50932 17500
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50876 16882 50932 16894
rect 50876 16830 50878 16882
rect 50930 16830 50932 16882
rect 50764 16772 50820 16782
rect 50764 16678 50820 16716
rect 50540 16324 50596 16334
rect 50540 16230 50596 16268
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50428 15372 50596 15428
rect 50540 15314 50596 15372
rect 50540 15262 50542 15314
rect 50594 15262 50596 15314
rect 50540 15250 50596 15262
rect 50876 15204 50932 16830
rect 51100 16324 51156 19404
rect 51324 19236 51380 19404
rect 51884 19236 51940 19966
rect 51996 19906 52052 19918
rect 51996 19854 51998 19906
rect 52050 19854 52052 19906
rect 51996 19460 52052 19854
rect 51996 19394 52052 19404
rect 51324 19234 51492 19236
rect 51324 19182 51326 19234
rect 51378 19182 51492 19234
rect 51324 19180 51492 19182
rect 51324 19170 51380 19180
rect 51324 18452 51380 18462
rect 51324 18358 51380 18396
rect 51436 18340 51492 19180
rect 51660 19180 51940 19236
rect 52444 19236 52500 23662
rect 52556 23716 52612 25116
rect 52780 25060 52836 25070
rect 52780 24946 52836 25004
rect 52780 24894 52782 24946
rect 52834 24894 52836 24946
rect 52780 24276 52836 24894
rect 52780 24210 52836 24220
rect 52892 24052 52948 25788
rect 53004 24498 53060 26852
rect 53452 26628 53508 27580
rect 53340 26572 53508 26628
rect 53564 27074 53620 27086
rect 53564 27022 53566 27074
rect 53618 27022 53620 27074
rect 53564 26628 53620 27022
rect 53004 24446 53006 24498
rect 53058 24446 53060 24498
rect 53004 24434 53060 24446
rect 53116 26178 53172 26190
rect 53116 26126 53118 26178
rect 53170 26126 53172 26178
rect 52780 23996 52948 24052
rect 52556 23650 52612 23660
rect 52668 23940 52724 23950
rect 52668 23604 52724 23884
rect 52668 23538 52724 23548
rect 52556 22596 52612 22606
rect 52556 22502 52612 22540
rect 52556 22372 52612 22382
rect 52556 22258 52612 22316
rect 52556 22206 52558 22258
rect 52610 22206 52612 22258
rect 52556 22194 52612 22206
rect 52668 22258 52724 22270
rect 52668 22206 52670 22258
rect 52722 22206 52724 22258
rect 52668 21924 52724 22206
rect 52668 21858 52724 21868
rect 52668 21476 52724 21486
rect 52668 20578 52724 21420
rect 52668 20526 52670 20578
rect 52722 20526 52724 20578
rect 52444 19180 52612 19236
rect 51548 19124 51604 19134
rect 51548 19030 51604 19068
rect 51660 19010 51716 19180
rect 51660 18958 51662 19010
rect 51714 18958 51716 19010
rect 51660 18946 51716 18958
rect 51996 19010 52052 19022
rect 52444 19012 52500 19022
rect 51996 18958 51998 19010
rect 52050 18958 52052 19010
rect 51996 18900 52052 18958
rect 51996 18834 52052 18844
rect 52220 19010 52500 19012
rect 52220 18958 52446 19010
rect 52498 18958 52500 19010
rect 52220 18956 52500 18958
rect 51660 18676 51716 18686
rect 51660 18562 51716 18620
rect 51660 18510 51662 18562
rect 51714 18510 51716 18562
rect 51660 18498 51716 18510
rect 51884 18452 51940 18462
rect 51436 18284 51716 18340
rect 51324 18004 51380 18014
rect 51324 17890 51380 17948
rect 51324 17838 51326 17890
rect 51378 17838 51380 17890
rect 51324 17826 51380 17838
rect 51212 17668 51268 17678
rect 51212 17574 51268 17612
rect 51100 16268 51268 16324
rect 51100 15988 51156 15998
rect 51100 15894 51156 15932
rect 50764 15092 50932 15204
rect 50316 14914 50372 14924
rect 50204 14644 50260 14654
rect 50204 14550 50260 14588
rect 50540 14532 50596 14542
rect 50428 14476 50540 14532
rect 50316 14306 50372 14318
rect 50316 14254 50318 14306
rect 50370 14254 50372 14306
rect 50316 13972 50372 14254
rect 50428 13972 50484 14476
rect 50540 14438 50596 14476
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50540 13972 50596 13982
rect 50428 13970 50596 13972
rect 50428 13918 50542 13970
rect 50594 13918 50596 13970
rect 50428 13916 50596 13918
rect 50316 13906 50372 13916
rect 50540 13906 50596 13916
rect 49980 13794 50036 13804
rect 50876 13858 50932 15092
rect 50876 13806 50878 13858
rect 50930 13806 50932 13858
rect 49644 12898 49700 12908
rect 49756 13746 49812 13758
rect 49756 13694 49758 13746
rect 49810 13694 49812 13746
rect 49644 12740 49700 12750
rect 49420 12738 49700 12740
rect 49420 12686 49646 12738
rect 49698 12686 49700 12738
rect 49420 12684 49700 12686
rect 49196 11508 49252 11518
rect 49196 11414 49252 11452
rect 49084 10882 49140 10892
rect 49084 10612 49140 10622
rect 49084 9938 49140 10556
rect 49084 9886 49086 9938
rect 49138 9886 49140 9938
rect 49084 9874 49140 9886
rect 48972 8318 48974 8370
rect 49026 8318 49028 8370
rect 48972 8306 49028 8318
rect 49420 8148 49476 12684
rect 49644 12674 49700 12684
rect 49532 12516 49588 12526
rect 49532 12402 49588 12460
rect 49532 12350 49534 12402
rect 49586 12350 49588 12402
rect 49532 12338 49588 12350
rect 49644 11172 49700 11182
rect 49644 11078 49700 11116
rect 49532 10836 49588 10846
rect 49532 10742 49588 10780
rect 49756 10500 49812 13694
rect 49980 13634 50036 13646
rect 49980 13582 49982 13634
rect 50034 13582 50036 13634
rect 49756 10434 49812 10444
rect 49868 12964 49924 12974
rect 49868 12292 49924 12908
rect 49868 12178 49924 12236
rect 49868 12126 49870 12178
rect 49922 12126 49924 12178
rect 49644 9938 49700 9950
rect 49644 9886 49646 9938
rect 49698 9886 49700 9938
rect 49532 8372 49588 8382
rect 49532 8278 49588 8316
rect 49420 8082 49476 8092
rect 48860 7298 48916 7308
rect 49084 8036 49140 8046
rect 48636 6514 48692 6524
rect 48524 6066 48580 6076
rect 48748 5236 48804 5246
rect 48412 5234 48804 5236
rect 48412 5182 48750 5234
rect 48802 5182 48804 5234
rect 48412 5180 48804 5182
rect 48748 5170 48804 5180
rect 47740 4562 47908 4564
rect 47740 4510 47742 4562
rect 47794 4510 47908 4562
rect 47740 4508 47908 4510
rect 47292 4498 47348 4508
rect 47740 4498 47796 4508
rect 48524 4452 48580 4462
rect 48524 4358 48580 4396
rect 48300 4338 48356 4350
rect 48300 4286 48302 4338
rect 48354 4286 48356 4338
rect 47964 4228 48020 4238
rect 47964 3666 48020 4172
rect 48300 4228 48356 4286
rect 48300 4162 48356 4172
rect 47964 3614 47966 3666
rect 48018 3614 48020 3666
rect 47964 3602 48020 3614
rect 44268 3556 44324 3566
rect 44268 3388 44324 3500
rect 45164 3556 45220 3566
rect 45164 3462 45220 3500
rect 44268 3332 44436 3388
rect 39004 800 39060 3332
rect 41804 3266 41860 3276
rect 44380 800 44436 3332
rect 44940 3332 44996 3342
rect 44940 3238 44996 3276
rect 49084 2884 49140 7980
rect 49644 7812 49700 9886
rect 49868 9156 49924 12126
rect 49980 11394 50036 13582
rect 50428 13524 50484 13534
rect 50316 13300 50372 13310
rect 50316 12962 50372 13244
rect 50316 12910 50318 12962
rect 50370 12910 50372 12962
rect 50316 12898 50372 12910
rect 50092 12292 50148 12302
rect 50092 12178 50148 12236
rect 50092 12126 50094 12178
rect 50146 12126 50148 12178
rect 50092 12114 50148 12126
rect 49980 11342 49982 11394
rect 50034 11342 50036 11394
rect 49980 10724 50036 11342
rect 49980 10658 50036 10668
rect 50204 11396 50260 11406
rect 50204 10722 50260 11340
rect 50428 11394 50484 13468
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50764 12404 50820 12414
rect 50764 12178 50820 12348
rect 50764 12126 50766 12178
rect 50818 12126 50820 12178
rect 50764 12068 50820 12126
rect 50764 12002 50820 12012
rect 50876 11508 50932 13806
rect 50988 15426 51044 15438
rect 50988 15374 50990 15426
rect 51042 15374 51044 15426
rect 50988 13524 51044 15374
rect 51212 14532 51268 16268
rect 51548 15876 51604 15886
rect 51548 15782 51604 15820
rect 51212 14466 51268 14476
rect 51324 15764 51380 15774
rect 51100 14306 51156 14318
rect 51100 14254 51102 14306
rect 51154 14254 51156 14306
rect 51100 13972 51156 14254
rect 51100 13906 51156 13916
rect 50988 13458 51044 13468
rect 51100 13188 51156 13198
rect 50988 12292 51044 12302
rect 50988 12198 51044 12236
rect 51100 11844 51156 13132
rect 51324 12740 51380 15708
rect 51436 15426 51492 15438
rect 51436 15374 51438 15426
rect 51490 15374 51492 15426
rect 51436 15204 51492 15374
rect 51436 15138 51492 15148
rect 51436 14644 51492 14654
rect 51436 14418 51492 14588
rect 51436 14366 51438 14418
rect 51490 14366 51492 14418
rect 51436 14196 51492 14366
rect 51436 14130 51492 14140
rect 51548 14532 51604 14542
rect 51436 13972 51492 13982
rect 51548 13972 51604 14476
rect 51436 13970 51604 13972
rect 51436 13918 51438 13970
rect 51490 13918 51604 13970
rect 51436 13916 51604 13918
rect 51436 13906 51492 13916
rect 51100 11778 51156 11788
rect 51212 12684 51380 12740
rect 51436 12850 51492 12862
rect 51436 12798 51438 12850
rect 51490 12798 51492 12850
rect 50764 11452 50932 11508
rect 51100 11508 51156 11518
rect 50428 11342 50430 11394
rect 50482 11342 50484 11394
rect 50316 11284 50372 11294
rect 50316 11190 50372 11228
rect 50204 10670 50206 10722
rect 50258 10670 50260 10722
rect 50204 10658 50260 10670
rect 50316 10834 50372 10846
rect 50316 10782 50318 10834
rect 50370 10782 50372 10834
rect 50092 10610 50148 10622
rect 50092 10558 50094 10610
rect 50146 10558 50148 10610
rect 49980 10500 50036 10510
rect 49980 9492 50036 10444
rect 50092 9716 50148 10558
rect 50316 10388 50372 10782
rect 50428 10724 50484 11342
rect 50652 11396 50708 11406
rect 50652 11302 50708 11340
rect 50764 11172 50820 11452
rect 51100 11414 51156 11452
rect 50764 11106 50820 11116
rect 50876 11284 50932 11294
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50540 10724 50596 10734
rect 50428 10722 50596 10724
rect 50428 10670 50542 10722
rect 50594 10670 50596 10722
rect 50428 10668 50596 10670
rect 50204 10332 50372 10388
rect 50204 9826 50260 10332
rect 50316 9940 50372 9950
rect 50316 9846 50372 9884
rect 50204 9774 50206 9826
rect 50258 9774 50260 9826
rect 50204 9762 50260 9774
rect 50092 9650 50148 9660
rect 50428 9716 50484 9726
rect 50316 9604 50372 9614
rect 49980 9436 50148 9492
rect 49868 9100 50036 9156
rect 49868 8932 49924 8942
rect 49420 7756 49700 7812
rect 49756 8930 49924 8932
rect 49756 8878 49870 8930
rect 49922 8878 49924 8930
rect 49756 8876 49924 8878
rect 49196 6804 49252 6814
rect 49196 6710 49252 6748
rect 49308 6692 49364 6702
rect 49308 6598 49364 6636
rect 49420 5908 49476 7756
rect 49644 7588 49700 7598
rect 49420 5842 49476 5852
rect 49532 7586 49700 7588
rect 49532 7534 49646 7586
rect 49698 7534 49700 7586
rect 49532 7532 49700 7534
rect 49532 6804 49588 7532
rect 49644 7522 49700 7532
rect 49756 7588 49812 8876
rect 49868 8866 49924 8876
rect 49868 8372 49924 8382
rect 49980 8372 50036 9100
rect 49868 8370 50036 8372
rect 49868 8318 49870 8370
rect 49922 8318 50036 8370
rect 49868 8316 50036 8318
rect 49868 8306 49924 8316
rect 49980 8036 50036 8316
rect 49980 7970 50036 7980
rect 50092 7700 50148 9436
rect 50316 9042 50372 9548
rect 50316 8990 50318 9042
rect 50370 8990 50372 9042
rect 50316 8978 50372 8990
rect 50092 7634 50148 7644
rect 50316 8034 50372 8046
rect 50316 7982 50318 8034
rect 50370 7982 50372 8034
rect 49756 7586 49924 7588
rect 49756 7534 49758 7586
rect 49810 7534 49924 7586
rect 49756 7532 49924 7534
rect 49756 7522 49812 7532
rect 49644 7252 49700 7262
rect 49644 7158 49700 7196
rect 49532 5906 49588 6748
rect 49868 6692 49924 7532
rect 50204 7364 50260 7374
rect 50204 7270 50260 7308
rect 50316 7252 50372 7982
rect 50316 7186 50372 7196
rect 49756 6132 49812 6142
rect 49756 6038 49812 6076
rect 49868 6018 49924 6636
rect 49868 5966 49870 6018
rect 49922 5966 49924 6018
rect 49868 5954 49924 5966
rect 49980 6468 50036 6478
rect 49532 5854 49534 5906
rect 49586 5854 49588 5906
rect 49532 5842 49588 5854
rect 49196 5346 49252 5358
rect 49196 5294 49198 5346
rect 49250 5294 49252 5346
rect 49196 5234 49252 5294
rect 49196 5182 49198 5234
rect 49250 5182 49252 5234
rect 49196 5170 49252 5182
rect 49644 5122 49700 5134
rect 49644 5070 49646 5122
rect 49698 5070 49700 5122
rect 49644 5012 49700 5070
rect 49644 3668 49700 4956
rect 49644 3602 49700 3612
rect 49980 3388 50036 6412
rect 50316 5796 50372 5806
rect 50316 5702 50372 5740
rect 50428 5234 50484 9660
rect 50540 9604 50596 10668
rect 50540 9538 50596 9548
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50764 9156 50820 9166
rect 50764 9042 50820 9100
rect 50764 8990 50766 9042
rect 50818 8990 50820 9042
rect 50764 8978 50820 8990
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50652 7700 50708 7710
rect 50652 7606 50708 7644
rect 50652 6692 50708 6702
rect 50652 6598 50708 6636
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 50876 6020 50932 11228
rect 51212 11284 51268 12684
rect 51436 12628 51492 12798
rect 51436 12562 51492 12572
rect 51660 12628 51716 18284
rect 51884 17444 51940 18396
rect 51884 17378 51940 17388
rect 52108 18116 52164 18126
rect 51772 17332 51828 17342
rect 51772 17106 51828 17276
rect 51772 17054 51774 17106
rect 51826 17054 51828 17106
rect 51772 17042 51828 17054
rect 51996 17220 52052 17230
rect 51996 17106 52052 17164
rect 51996 17054 51998 17106
rect 52050 17054 52052 17106
rect 51996 17042 52052 17054
rect 51884 16770 51940 16782
rect 51884 16718 51886 16770
rect 51938 16718 51940 16770
rect 51772 15316 51828 15326
rect 51772 15222 51828 15260
rect 51772 13746 51828 13758
rect 51772 13694 51774 13746
rect 51826 13694 51828 13746
rect 51772 13524 51828 13694
rect 51772 13458 51828 13468
rect 51884 13188 51940 16718
rect 51996 16324 52052 16334
rect 51996 16210 52052 16268
rect 51996 16158 51998 16210
rect 52050 16158 52052 16210
rect 51996 16146 52052 16158
rect 52108 15148 52164 18060
rect 52220 16548 52276 18956
rect 52444 18946 52500 18956
rect 52444 18116 52500 18126
rect 52332 17442 52388 17454
rect 52332 17390 52334 17442
rect 52386 17390 52388 17442
rect 52332 17108 52388 17390
rect 52332 17042 52388 17052
rect 52444 16882 52500 18060
rect 52556 18004 52612 19180
rect 52668 18564 52724 20526
rect 52780 21026 52836 23996
rect 53004 23940 53060 23950
rect 52892 23884 53004 23940
rect 52892 21810 52948 23884
rect 53004 23874 53060 23884
rect 53004 23716 53060 23726
rect 53004 22372 53060 23660
rect 53116 22820 53172 26126
rect 53228 24612 53284 24622
rect 53228 24518 53284 24556
rect 53340 23492 53396 26572
rect 53564 26562 53620 26572
rect 53788 27076 53844 27086
rect 53788 26850 53844 27020
rect 53788 26798 53790 26850
rect 53842 26798 53844 26850
rect 53452 26404 53508 26414
rect 53452 26290 53508 26348
rect 53452 26238 53454 26290
rect 53506 26238 53508 26290
rect 53452 26180 53508 26238
rect 53452 26114 53508 26124
rect 53676 26290 53732 26302
rect 53676 26238 53678 26290
rect 53730 26238 53732 26290
rect 53676 26068 53732 26238
rect 53452 25284 53508 25294
rect 53676 25284 53732 26012
rect 53788 25506 53844 26798
rect 53900 26516 53956 27580
rect 53900 26450 53956 26460
rect 54012 26404 54068 27804
rect 54012 26338 54068 26348
rect 53788 25454 53790 25506
rect 53842 25454 53844 25506
rect 53788 25442 53844 25454
rect 53452 25282 53620 25284
rect 53452 25230 53454 25282
rect 53506 25230 53620 25282
rect 53452 25228 53620 25230
rect 53676 25228 54068 25284
rect 53452 25218 53508 25228
rect 53452 23940 53508 23950
rect 53452 23846 53508 23884
rect 53564 23604 53620 25228
rect 53900 24836 53956 24846
rect 53788 24834 53956 24836
rect 53788 24782 53902 24834
rect 53954 24782 53956 24834
rect 53788 24780 53956 24782
rect 53564 23538 53620 23548
rect 53676 24498 53732 24510
rect 53676 24446 53678 24498
rect 53730 24446 53732 24498
rect 53676 23938 53732 24446
rect 53676 23886 53678 23938
rect 53730 23886 53732 23938
rect 53116 22754 53172 22764
rect 53228 23436 53396 23492
rect 53004 22306 53060 22316
rect 52892 21758 52894 21810
rect 52946 21758 52948 21810
rect 52892 21746 52948 21758
rect 53228 21700 53284 23436
rect 53676 23380 53732 23886
rect 53340 23324 53732 23380
rect 53340 23154 53396 23324
rect 53340 23102 53342 23154
rect 53394 23102 53396 23154
rect 53340 23090 53396 23102
rect 53788 23268 53844 24780
rect 53900 24770 53956 24780
rect 54012 24500 54068 25228
rect 54124 24836 54180 29148
rect 54236 29138 54292 29148
rect 54572 28642 54628 28654
rect 54572 28590 54574 28642
rect 54626 28590 54628 28642
rect 54572 27972 54628 28590
rect 54684 28644 54740 28654
rect 54684 28082 54740 28588
rect 54684 28030 54686 28082
rect 54738 28030 54740 28082
rect 54684 28018 54740 28030
rect 55020 28644 55076 28654
rect 54236 27748 54292 27786
rect 54236 27682 54292 27692
rect 54236 27524 54292 27534
rect 54236 25620 54292 27468
rect 54348 27076 54404 27086
rect 54348 26982 54404 27020
rect 54572 26908 54628 27916
rect 54460 26852 54628 26908
rect 54684 27412 54740 27422
rect 54460 26178 54516 26852
rect 54684 26850 54740 27356
rect 54684 26798 54686 26850
rect 54738 26798 54740 26850
rect 54684 26786 54740 26798
rect 54908 26404 54964 26414
rect 54908 26310 54964 26348
rect 54460 26126 54462 26178
rect 54514 26126 54516 26178
rect 54236 25564 54404 25620
rect 54236 25396 54292 25406
rect 54236 25302 54292 25340
rect 54124 24722 54180 24780
rect 54124 24670 54126 24722
rect 54178 24670 54180 24722
rect 54124 24658 54180 24670
rect 54012 24444 54180 24500
rect 54012 23828 54068 23866
rect 54012 23762 54068 23772
rect 53900 23716 53956 23726
rect 53900 23622 53956 23660
rect 54012 23604 54068 23614
rect 53452 23042 53508 23054
rect 53452 22990 53454 23042
rect 53506 22990 53508 23042
rect 53228 21634 53284 21644
rect 53340 22930 53396 22942
rect 53340 22878 53342 22930
rect 53394 22878 53396 22930
rect 53228 21476 53284 21486
rect 53228 21382 53284 21420
rect 52780 20974 52782 21026
rect 52834 20974 52836 21026
rect 52780 20244 52836 20974
rect 52780 20178 52836 20188
rect 52892 21362 52948 21374
rect 52892 21310 52894 21362
rect 52946 21310 52948 21362
rect 52892 20020 52948 21310
rect 52892 19572 52948 19964
rect 52892 19506 52948 19516
rect 53004 20580 53060 20590
rect 53340 20580 53396 22878
rect 53452 22820 53508 22990
rect 53452 22754 53508 22764
rect 53788 22372 53844 23212
rect 53900 23380 53956 23390
rect 53900 22708 53956 23324
rect 54012 23154 54068 23548
rect 54012 23102 54014 23154
rect 54066 23102 54068 23154
rect 54012 23090 54068 23102
rect 53900 22642 53956 22652
rect 54012 22596 54068 22606
rect 54124 22596 54180 24444
rect 54068 22540 54180 22596
rect 53900 22372 53956 22382
rect 53788 22370 53956 22372
rect 53788 22318 53902 22370
rect 53954 22318 53956 22370
rect 53788 22316 53956 22318
rect 53900 22306 53956 22316
rect 54012 22370 54068 22540
rect 54012 22318 54014 22370
rect 54066 22318 54068 22370
rect 54012 22306 54068 22318
rect 54236 22370 54292 22382
rect 54236 22318 54238 22370
rect 54290 22318 54292 22370
rect 53676 22260 53732 22270
rect 53452 22146 53508 22158
rect 53452 22094 53454 22146
rect 53506 22094 53508 22146
rect 53452 22036 53508 22094
rect 53452 21970 53508 21980
rect 53676 21810 53732 22204
rect 53676 21758 53678 21810
rect 53730 21758 53732 21810
rect 53676 21746 53732 21758
rect 53788 22036 53844 22046
rect 53004 20018 53060 20524
rect 53228 20524 53396 20580
rect 53452 20802 53508 20814
rect 53452 20750 53454 20802
rect 53506 20750 53508 20802
rect 53452 20580 53508 20750
rect 53788 20804 53844 21980
rect 54236 21924 54292 22318
rect 54236 21858 54292 21868
rect 54236 21700 54292 21710
rect 54124 21588 54180 21598
rect 54124 21494 54180 21532
rect 54012 20916 54068 20926
rect 53788 20802 53956 20804
rect 53788 20750 53790 20802
rect 53842 20750 53956 20802
rect 53788 20748 53956 20750
rect 53788 20738 53844 20748
rect 53228 20244 53284 20524
rect 53452 20514 53508 20524
rect 53004 19966 53006 20018
rect 53058 19966 53060 20018
rect 52668 18498 52724 18508
rect 52780 18452 52836 18462
rect 52780 18116 52836 18396
rect 52780 18050 52836 18060
rect 52556 17938 52612 17948
rect 52444 16830 52446 16882
rect 52498 16830 52500 16882
rect 52444 16818 52500 16830
rect 52556 17668 52612 17678
rect 53004 17668 53060 19966
rect 52556 17666 53060 17668
rect 52556 17614 52558 17666
rect 52610 17614 53060 17666
rect 52556 17612 53060 17614
rect 53116 20188 53284 20244
rect 53340 20244 53396 20254
rect 52556 16660 52612 17612
rect 52220 16324 52276 16492
rect 52220 16258 52276 16268
rect 52332 16604 52612 16660
rect 52668 17108 52724 17118
rect 52108 15082 52164 15092
rect 52108 14980 52164 14990
rect 52332 14980 52388 16604
rect 52444 16212 52500 16222
rect 52668 16212 52724 17052
rect 53004 17108 53060 17118
rect 53004 17014 53060 17052
rect 52444 16210 52724 16212
rect 52444 16158 52446 16210
rect 52498 16158 52724 16210
rect 52444 16156 52724 16158
rect 52444 15092 52500 16156
rect 53116 15876 53172 20188
rect 53340 20020 53396 20188
rect 53228 19964 53396 20020
rect 53788 20020 53844 20030
rect 53228 17332 53284 19964
rect 53788 19926 53844 19964
rect 53340 19572 53396 19582
rect 53340 19346 53396 19516
rect 53340 19294 53342 19346
rect 53394 19294 53396 19346
rect 53340 19282 53396 19294
rect 53900 18900 53956 20748
rect 54012 20802 54068 20860
rect 54012 20750 54014 20802
rect 54066 20750 54068 20802
rect 54012 20738 54068 20750
rect 54124 20804 54180 20814
rect 54124 20710 54180 20748
rect 54236 20802 54292 21644
rect 54236 20750 54238 20802
rect 54290 20750 54292 20802
rect 54124 20468 54180 20478
rect 54012 19012 54068 19022
rect 54012 18918 54068 18956
rect 53900 18834 53956 18844
rect 53452 18564 53508 18574
rect 54124 18564 54180 20412
rect 53340 18562 53508 18564
rect 53340 18510 53454 18562
rect 53506 18510 53508 18562
rect 53340 18508 53508 18510
rect 53340 18340 53396 18508
rect 53452 18498 53508 18508
rect 54012 18508 54180 18564
rect 53676 18452 53732 18462
rect 53676 18358 53732 18396
rect 53900 18452 53956 18462
rect 53900 18358 53956 18396
rect 53340 17444 53396 18284
rect 53452 17668 53508 17678
rect 53452 17574 53508 17612
rect 53340 17378 53396 17388
rect 53788 17442 53844 17454
rect 53788 17390 53790 17442
rect 53842 17390 53844 17442
rect 53228 17266 53284 17276
rect 53788 17108 53844 17390
rect 53788 17042 53844 17052
rect 53452 16996 53508 17006
rect 53452 16902 53508 16940
rect 53228 16882 53284 16894
rect 53900 16884 53956 16894
rect 53228 16830 53230 16882
rect 53282 16830 53284 16882
rect 53228 16324 53284 16830
rect 53676 16882 53956 16884
rect 53676 16830 53902 16882
rect 53954 16830 53956 16882
rect 53676 16828 53956 16830
rect 53340 16772 53396 16782
rect 53340 16770 53508 16772
rect 53340 16718 53342 16770
rect 53394 16718 53508 16770
rect 53340 16716 53508 16718
rect 53340 16706 53396 16716
rect 53228 16258 53284 16268
rect 52892 15820 53172 15876
rect 53340 15876 53396 15886
rect 52892 15538 52948 15820
rect 53340 15782 53396 15820
rect 52892 15486 52894 15538
rect 52946 15486 52948 15538
rect 52668 15428 52724 15438
rect 52668 15334 52724 15372
rect 52556 15316 52612 15326
rect 52556 15222 52612 15260
rect 52780 15204 52836 15214
rect 52668 15092 52836 15148
rect 52444 15036 52612 15092
rect 52164 14924 52276 14980
rect 52108 14914 52164 14924
rect 52220 13748 52276 14924
rect 52332 14914 52388 14924
rect 52220 13654 52276 13692
rect 52332 14756 52388 14766
rect 52220 13412 52276 13422
rect 51884 13132 52052 13188
rect 51660 12562 51716 12572
rect 51772 13076 51828 13086
rect 51660 12404 51716 12414
rect 51772 12404 51828 13020
rect 51660 12402 51828 12404
rect 51660 12350 51662 12402
rect 51714 12350 51828 12402
rect 51660 12348 51828 12350
rect 51884 12962 51940 12974
rect 51884 12910 51886 12962
rect 51938 12910 51940 12962
rect 51884 12740 51940 12910
rect 51996 12852 52052 13132
rect 51996 12786 52052 12796
rect 51660 12292 51716 12348
rect 51324 12236 51604 12292
rect 51324 12180 51380 12236
rect 51324 12114 51380 12124
rect 51548 12178 51604 12236
rect 51660 12226 51716 12236
rect 51548 12126 51550 12178
rect 51602 12126 51604 12178
rect 51548 12114 51604 12126
rect 51772 12180 51828 12190
rect 51212 10834 51268 11228
rect 51212 10782 51214 10834
rect 51266 10782 51268 10834
rect 51212 10770 51268 10782
rect 51436 12068 51492 12078
rect 51100 10724 51156 10734
rect 51100 10630 51156 10668
rect 51212 10386 51268 10398
rect 51212 10334 51214 10386
rect 51266 10334 51268 10386
rect 51100 10164 51156 10174
rect 50988 8148 51044 8158
rect 50988 8054 51044 8092
rect 51100 7588 51156 10108
rect 51212 9940 51268 10334
rect 51212 9874 51268 9884
rect 51436 9828 51492 12012
rect 51660 11954 51716 11966
rect 51660 11902 51662 11954
rect 51714 11902 51716 11954
rect 51660 11844 51716 11902
rect 51660 11778 51716 11788
rect 51660 11620 51716 11630
rect 51660 11506 51716 11564
rect 51660 11454 51662 11506
rect 51714 11454 51716 11506
rect 51660 11442 51716 11454
rect 51548 11396 51604 11406
rect 51548 10050 51604 11340
rect 51772 10834 51828 12124
rect 51884 11620 51940 12684
rect 52220 12402 52276 13356
rect 52220 12350 52222 12402
rect 52274 12350 52276 12402
rect 52220 12338 52276 12350
rect 51884 11554 51940 11564
rect 51996 12292 52052 12302
rect 51772 10782 51774 10834
rect 51826 10782 51828 10834
rect 51772 10770 51828 10782
rect 51548 9998 51550 10050
rect 51602 9998 51604 10050
rect 51548 9986 51604 9998
rect 51660 10164 51716 10174
rect 51436 9772 51604 9828
rect 51324 9716 51380 9726
rect 51324 9622 51380 9660
rect 51436 9602 51492 9614
rect 51436 9550 51438 9602
rect 51490 9550 51492 9602
rect 51436 9268 51492 9550
rect 51324 9212 51492 9268
rect 51324 9156 51380 9212
rect 51324 9090 51380 9100
rect 51436 9044 51492 9054
rect 51548 9044 51604 9772
rect 51436 9042 51604 9044
rect 51436 8990 51438 9042
rect 51490 8990 51604 9042
rect 51436 8988 51604 8990
rect 51436 8978 51492 8988
rect 51660 8372 51716 10108
rect 51884 9604 51940 9614
rect 51884 9266 51940 9548
rect 51884 9214 51886 9266
rect 51938 9214 51940 9266
rect 51884 9044 51940 9214
rect 51884 8978 51940 8988
rect 51996 8820 52052 12236
rect 52220 11620 52276 11630
rect 52108 9940 52164 9950
rect 52108 9716 52164 9884
rect 52108 9622 52164 9660
rect 51548 8316 51716 8372
rect 51884 8764 52052 8820
rect 50988 7532 51156 7588
rect 51212 8036 51268 8046
rect 50988 6580 51044 7532
rect 51100 7362 51156 7374
rect 51100 7310 51102 7362
rect 51154 7310 51156 7362
rect 51100 7028 51156 7310
rect 51100 6962 51156 6972
rect 50988 6514 51044 6524
rect 51212 6132 51268 7980
rect 51548 7700 51604 8316
rect 51660 8148 51716 8158
rect 51660 8054 51716 8092
rect 51772 8036 51828 8046
rect 51772 7942 51828 7980
rect 51660 7700 51716 7710
rect 51548 7698 51716 7700
rect 51548 7646 51662 7698
rect 51714 7646 51716 7698
rect 51548 7644 51716 7646
rect 51660 7634 51716 7644
rect 51324 6916 51380 6926
rect 51324 6822 51380 6860
rect 51324 6132 51380 6142
rect 51212 6130 51380 6132
rect 51212 6078 51326 6130
rect 51378 6078 51380 6130
rect 51212 6076 51380 6078
rect 51324 6066 51380 6076
rect 50876 5964 51044 6020
rect 50876 5794 50932 5806
rect 50876 5742 50878 5794
rect 50930 5742 50932 5794
rect 50876 5682 50932 5742
rect 50876 5630 50878 5682
rect 50930 5630 50932 5682
rect 50876 5618 50932 5630
rect 50428 5182 50430 5234
rect 50482 5182 50484 5234
rect 50428 5124 50484 5182
rect 50988 5236 51044 5964
rect 51772 5796 51828 5806
rect 51884 5796 51940 8764
rect 51996 8372 52052 8382
rect 51996 8258 52052 8316
rect 51996 8206 51998 8258
rect 52050 8206 52052 8258
rect 51996 8194 52052 8206
rect 51996 7362 52052 7374
rect 51996 7310 51998 7362
rect 52050 7310 52052 7362
rect 51996 7252 52052 7310
rect 51996 7186 52052 7196
rect 52108 6580 52164 6590
rect 51996 6468 52052 6478
rect 51996 6374 52052 6412
rect 51772 5794 51940 5796
rect 51772 5742 51774 5794
rect 51826 5742 51940 5794
rect 51772 5740 51940 5742
rect 51772 5682 51828 5740
rect 51772 5630 51774 5682
rect 51826 5630 51828 5682
rect 51772 5618 51828 5630
rect 51660 5236 51716 5246
rect 50988 5234 51716 5236
rect 50988 5182 50990 5234
rect 51042 5182 51662 5234
rect 51714 5182 51716 5234
rect 50988 5180 51716 5182
rect 50988 5170 51044 5180
rect 51660 5170 51716 5180
rect 52108 5234 52164 6524
rect 52220 6132 52276 11564
rect 52332 9940 52388 14700
rect 52556 14532 52612 15036
rect 52668 14754 52724 15092
rect 52668 14702 52670 14754
rect 52722 14702 52724 14754
rect 52668 14690 52724 14702
rect 52556 14476 52836 14532
rect 52444 14306 52500 14318
rect 52444 14254 52446 14306
rect 52498 14254 52500 14306
rect 52444 14196 52500 14254
rect 52556 14308 52612 14318
rect 52556 14214 52612 14252
rect 52444 14130 52500 14140
rect 52444 13972 52500 13982
rect 52444 13878 52500 13916
rect 52556 13746 52612 13758
rect 52556 13694 52558 13746
rect 52610 13694 52612 13746
rect 52556 13524 52612 13694
rect 52556 13458 52612 13468
rect 52668 13076 52724 13086
rect 52668 12982 52724 13020
rect 52556 12740 52612 12750
rect 52332 9874 52388 9884
rect 52444 11732 52500 11742
rect 52444 11282 52500 11676
rect 52556 11396 52612 12684
rect 52668 12068 52724 12078
rect 52668 11974 52724 12012
rect 52556 11340 52724 11396
rect 52444 11230 52446 11282
rect 52498 11230 52500 11282
rect 52444 9716 52500 11230
rect 52556 11172 52612 11182
rect 52556 11078 52612 11116
rect 52556 9940 52612 9950
rect 52556 9846 52612 9884
rect 52332 9660 52500 9716
rect 52332 6468 52388 9660
rect 52668 9156 52724 11340
rect 52780 10948 52836 14476
rect 52892 14420 52948 15486
rect 53228 15316 53284 15326
rect 53228 15222 53284 15260
rect 53340 15204 53396 15214
rect 52892 14354 52948 14364
rect 53004 15092 53396 15148
rect 53004 12740 53060 15092
rect 53004 12674 53060 12684
rect 53116 14980 53172 14990
rect 53116 13858 53172 14924
rect 53452 14756 53508 16716
rect 53676 15540 53732 16828
rect 53900 16818 53956 16828
rect 53900 16212 53956 16222
rect 54012 16212 54068 18508
rect 53900 16210 54068 16212
rect 53900 16158 53902 16210
rect 53954 16158 54068 16210
rect 53900 16156 54068 16158
rect 54124 18004 54180 18014
rect 54124 16994 54180 17948
rect 54236 17668 54292 20750
rect 54348 20916 54404 25564
rect 54460 25172 54516 26126
rect 54796 25284 54852 25294
rect 54796 25282 54964 25284
rect 54796 25230 54798 25282
rect 54850 25230 54964 25282
rect 54796 25228 54964 25230
rect 54796 25218 54852 25228
rect 54460 25106 54516 25116
rect 54796 24836 54852 24846
rect 54796 24742 54852 24780
rect 54908 24612 54964 25228
rect 54908 24546 54964 24556
rect 55020 23938 55076 28588
rect 55356 28642 55412 30268
rect 55580 30098 55636 30110
rect 55580 30046 55582 30098
rect 55634 30046 55636 30098
rect 55468 29988 55524 29998
rect 55468 29894 55524 29932
rect 55580 29540 55636 30046
rect 55580 29474 55636 29484
rect 55356 28590 55358 28642
rect 55410 28590 55412 28642
rect 55356 28578 55412 28590
rect 55692 28418 55748 28430
rect 55692 28366 55694 28418
rect 55746 28366 55748 28418
rect 55468 27972 55524 27982
rect 55468 27878 55524 27916
rect 55692 27858 55748 28366
rect 55692 27806 55694 27858
rect 55746 27806 55748 27858
rect 55580 26962 55636 26974
rect 55580 26910 55582 26962
rect 55634 26910 55636 26962
rect 55244 26850 55300 26862
rect 55244 26798 55246 26850
rect 55298 26798 55300 26850
rect 55244 25620 55300 26798
rect 55244 25554 55300 25564
rect 55356 26628 55412 26638
rect 55356 26178 55412 26572
rect 55356 26126 55358 26178
rect 55410 26126 55412 26178
rect 55132 25508 55188 25518
rect 55132 25414 55188 25452
rect 55356 25172 55412 26126
rect 55356 25106 55412 25116
rect 55132 24836 55188 24846
rect 55132 24834 55300 24836
rect 55132 24782 55134 24834
rect 55186 24782 55300 24834
rect 55132 24780 55300 24782
rect 55132 24770 55188 24780
rect 55020 23886 55022 23938
rect 55074 23886 55076 23938
rect 55020 23874 55076 23886
rect 55132 24164 55188 24174
rect 55020 23380 55076 23390
rect 55132 23380 55188 24108
rect 55076 23324 55188 23380
rect 55244 23380 55300 24780
rect 55020 23248 55076 23324
rect 55244 23314 55300 23324
rect 55468 24500 55524 24510
rect 55468 23378 55524 24444
rect 55468 23326 55470 23378
rect 55522 23326 55524 23378
rect 55468 23314 55524 23326
rect 55580 23380 55636 26910
rect 55692 25508 55748 27806
rect 55804 27636 55860 30718
rect 55804 27570 55860 27580
rect 55692 25442 55748 25452
rect 55916 25172 55972 31500
rect 56252 31490 56308 31500
rect 56364 31556 56420 32398
rect 56700 31892 56756 39342
rect 56700 31826 56756 31836
rect 56812 32450 56868 32462
rect 56812 32398 56814 32450
rect 56866 32398 56868 32450
rect 56364 31490 56420 31500
rect 56140 30882 56196 30894
rect 56140 30830 56142 30882
rect 56194 30830 56196 30882
rect 56140 30770 56196 30830
rect 56140 30718 56142 30770
rect 56194 30718 56196 30770
rect 56140 30706 56196 30718
rect 56700 30882 56756 30894
rect 56700 30830 56702 30882
rect 56754 30830 56756 30882
rect 56700 30660 56756 30830
rect 56476 30098 56532 30110
rect 56476 30046 56478 30098
rect 56530 30046 56532 30098
rect 56140 29986 56196 29998
rect 56140 29934 56142 29986
rect 56194 29934 56196 29986
rect 56028 29314 56084 29326
rect 56028 29262 56030 29314
rect 56082 29262 56084 29314
rect 56028 28980 56084 29262
rect 56028 28914 56084 28924
rect 56140 28756 56196 29934
rect 56140 28690 56196 28700
rect 56364 29876 56420 29886
rect 56364 29316 56420 29820
rect 56364 28532 56420 29260
rect 56252 28530 56420 28532
rect 56252 28478 56366 28530
rect 56418 28478 56420 28530
rect 56252 28476 56420 28478
rect 56252 27636 56308 28476
rect 56364 28466 56420 28476
rect 56476 28532 56532 30046
rect 56700 29650 56756 30604
rect 56700 29598 56702 29650
rect 56754 29598 56756 29650
rect 56588 29540 56644 29550
rect 56588 28642 56644 29484
rect 56588 28590 56590 28642
rect 56642 28590 56644 28642
rect 56588 28578 56644 28590
rect 56700 28644 56756 29598
rect 56812 29652 56868 32398
rect 57372 32452 57428 32462
rect 57372 32358 57428 32396
rect 56924 31892 56980 31902
rect 57260 31892 57316 31902
rect 56924 31890 57316 31892
rect 56924 31838 56926 31890
rect 56978 31838 57262 31890
rect 57314 31838 57316 31890
rect 56924 31836 57316 31838
rect 56924 29876 56980 31836
rect 57260 31826 57316 31836
rect 57148 31556 57204 31566
rect 57036 30660 57092 30670
rect 57036 30210 57092 30604
rect 57036 30158 57038 30210
rect 57090 30158 57092 30210
rect 57036 30146 57092 30158
rect 56924 29810 56980 29820
rect 56812 29596 56980 29652
rect 56700 28578 56756 28588
rect 56476 28466 56532 28476
rect 56588 28420 56644 28430
rect 56364 27970 56420 27982
rect 56364 27918 56366 27970
rect 56418 27918 56420 27970
rect 56364 27860 56420 27918
rect 56364 27794 56420 27804
rect 56252 27580 56420 27636
rect 56252 27300 56308 27310
rect 56252 27206 56308 27244
rect 56028 26402 56084 26414
rect 56028 26350 56030 26402
rect 56082 26350 56084 26402
rect 56028 25732 56084 26350
rect 56028 25666 56084 25676
rect 56252 26292 56308 26302
rect 55916 24948 55972 25116
rect 56028 25394 56084 25406
rect 56028 25342 56030 25394
rect 56082 25342 56084 25394
rect 56028 25060 56084 25342
rect 56028 24994 56084 25004
rect 56140 25284 56196 25294
rect 55580 23314 55636 23324
rect 55692 24892 55972 24948
rect 55244 23154 55300 23166
rect 55244 23102 55246 23154
rect 55298 23102 55300 23154
rect 55132 23044 55188 23054
rect 55132 22950 55188 22988
rect 55244 22596 55300 23102
rect 55244 22530 55300 22540
rect 55692 22820 55748 24892
rect 56028 24836 56084 24846
rect 56140 24836 56196 25228
rect 56028 24834 56196 24836
rect 56028 24782 56030 24834
rect 56082 24782 56196 24834
rect 56028 24780 56196 24782
rect 56028 24770 56084 24780
rect 56252 24724 56308 26236
rect 56364 25618 56420 27580
rect 56364 25566 56366 25618
rect 56418 25566 56420 25618
rect 56364 25172 56420 25566
rect 56588 27298 56644 28364
rect 56700 27860 56756 27870
rect 56700 27858 56868 27860
rect 56700 27806 56702 27858
rect 56754 27806 56868 27858
rect 56700 27804 56868 27806
rect 56700 27794 56756 27804
rect 56588 27246 56590 27298
rect 56642 27246 56644 27298
rect 56588 25620 56644 27246
rect 56812 27186 56868 27804
rect 56812 27134 56814 27186
rect 56866 27134 56868 27186
rect 56812 26852 56868 27134
rect 56812 26292 56868 26796
rect 56812 26226 56868 26236
rect 56588 25564 56868 25620
rect 56476 25508 56532 25518
rect 56532 25452 56756 25508
rect 56476 25414 56532 25452
rect 56364 25116 56644 25172
rect 56364 24724 56420 24734
rect 56252 24722 56420 24724
rect 56252 24670 56366 24722
rect 56418 24670 56420 24722
rect 56252 24668 56420 24670
rect 56364 24658 56420 24668
rect 56588 24722 56644 25116
rect 56588 24670 56590 24722
rect 56642 24670 56644 24722
rect 56588 24658 56644 24670
rect 56140 24612 56196 24622
rect 56140 24518 56196 24556
rect 55804 24500 55860 24510
rect 55804 24406 55860 24444
rect 54348 20244 54404 20860
rect 54684 22484 54740 22494
rect 54684 20914 54740 22428
rect 54796 22260 54852 22270
rect 54796 22166 54852 22204
rect 55132 22148 55188 22158
rect 55132 22054 55188 22092
rect 55580 22148 55636 22158
rect 55580 22054 55636 22092
rect 55132 21924 55188 21934
rect 54684 20862 54686 20914
rect 54738 20862 54740 20914
rect 54348 20178 54404 20188
rect 54572 20692 54628 20702
rect 54460 20020 54516 20030
rect 54348 19124 54404 19134
rect 54348 19030 54404 19068
rect 54348 18788 54404 18798
rect 54348 18562 54404 18732
rect 54460 18676 54516 19964
rect 54460 18610 54516 18620
rect 54348 18510 54350 18562
rect 54402 18510 54404 18562
rect 54348 18498 54404 18510
rect 54460 18452 54516 18462
rect 54460 18358 54516 18396
rect 54292 17612 54404 17668
rect 54236 17602 54292 17612
rect 54236 17444 54292 17454
rect 54236 17350 54292 17388
rect 54348 17220 54404 17612
rect 54124 16942 54126 16994
rect 54178 16942 54180 16994
rect 53900 16146 53956 16156
rect 54124 16100 54180 16942
rect 54236 17164 54404 17220
rect 54572 17220 54628 20636
rect 54684 20468 54740 20862
rect 54684 20402 54740 20412
rect 54796 21698 54852 21710
rect 54796 21646 54798 21698
rect 54850 21646 54852 21698
rect 54796 20244 54852 21646
rect 55020 21700 55076 21710
rect 55020 21606 55076 21644
rect 54684 20188 54852 20244
rect 54908 21474 54964 21486
rect 54908 21422 54910 21474
rect 54962 21422 54964 21474
rect 54684 18340 54740 20188
rect 54796 20020 54852 20030
rect 54796 19926 54852 19964
rect 54908 19124 54964 21422
rect 55132 21476 55188 21868
rect 55244 21700 55300 21710
rect 55692 21700 55748 22764
rect 55916 24388 55972 24398
rect 55244 21588 55300 21644
rect 55580 21644 55748 21700
rect 55804 22372 55860 22382
rect 55468 21588 55524 21598
rect 55244 21586 55524 21588
rect 55244 21534 55470 21586
rect 55522 21534 55524 21586
rect 55244 21532 55524 21534
rect 55468 21522 55524 21532
rect 55132 21420 55300 21476
rect 55244 21364 55300 21420
rect 55244 21308 55412 21364
rect 54908 19058 54964 19068
rect 55020 21028 55076 21038
rect 55020 19122 55076 20972
rect 55132 20020 55188 20030
rect 55132 19348 55188 19964
rect 55244 20018 55300 20030
rect 55244 19966 55246 20018
rect 55298 19966 55300 20018
rect 55244 19460 55300 19966
rect 55356 19906 55412 21308
rect 55580 20804 55636 21644
rect 55692 21476 55748 21486
rect 55692 21382 55748 21420
rect 55692 20804 55748 20814
rect 55580 20802 55748 20804
rect 55580 20750 55694 20802
rect 55746 20750 55748 20802
rect 55580 20748 55748 20750
rect 55580 20580 55636 20590
rect 55580 20486 55636 20524
rect 55356 19854 55358 19906
rect 55410 19854 55412 19906
rect 55356 19842 55412 19854
rect 55580 19794 55636 19806
rect 55580 19742 55582 19794
rect 55634 19742 55636 19794
rect 55580 19460 55636 19742
rect 55244 19404 55412 19460
rect 55356 19348 55412 19404
rect 55580 19394 55636 19404
rect 55132 19292 55300 19348
rect 55020 19070 55022 19122
rect 55074 19070 55076 19122
rect 54684 18274 54740 18284
rect 54796 18900 54852 18910
rect 54572 17164 54740 17220
rect 54236 16994 54292 17164
rect 54348 17108 54404 17164
rect 54348 17052 54628 17108
rect 54236 16942 54238 16994
rect 54290 16942 54292 16994
rect 54236 16930 54292 16942
rect 54460 16660 54516 16670
rect 54124 16034 54180 16044
rect 54348 16658 54516 16660
rect 54348 16606 54462 16658
rect 54514 16606 54516 16658
rect 54348 16604 54516 16606
rect 53676 15474 53732 15484
rect 54012 15988 54068 15998
rect 53676 15314 53732 15326
rect 53676 15262 53678 15314
rect 53730 15262 53732 15314
rect 53676 15204 53732 15262
rect 53900 15316 53956 15326
rect 54012 15316 54068 15932
rect 53900 15314 54068 15316
rect 53900 15262 53902 15314
rect 53954 15262 54068 15314
rect 53900 15260 54068 15262
rect 53900 15250 53956 15260
rect 53676 15138 53732 15148
rect 53340 14700 53508 14756
rect 53788 14868 53844 14878
rect 53116 13806 53118 13858
rect 53170 13806 53172 13858
rect 53116 12292 53172 13806
rect 53228 14308 53284 14318
rect 53228 12740 53284 14252
rect 53228 12674 53284 12684
rect 53340 12404 53396 14700
rect 53452 14530 53508 14542
rect 53452 14478 53454 14530
rect 53506 14478 53508 14530
rect 53452 13860 53508 14478
rect 53452 13766 53508 13804
rect 53564 14308 53620 14318
rect 53564 14084 53620 14252
rect 53564 13636 53620 14028
rect 53452 13580 53620 13636
rect 53788 13636 53844 14812
rect 53452 12852 53508 13580
rect 53788 13570 53844 13580
rect 53900 14642 53956 14654
rect 53900 14590 53902 14642
rect 53954 14590 53956 14642
rect 53900 13300 53956 14590
rect 54012 13412 54068 15260
rect 54124 15426 54180 15438
rect 54124 15374 54126 15426
rect 54178 15374 54180 15426
rect 54124 15092 54180 15374
rect 54124 15026 54180 15036
rect 54236 15316 54292 15326
rect 54236 15090 54292 15260
rect 54236 15038 54238 15090
rect 54290 15038 54292 15090
rect 54236 14530 54292 15038
rect 54236 14478 54238 14530
rect 54290 14478 54292 14530
rect 54236 14466 54292 14478
rect 54124 14420 54180 14430
rect 54124 14084 54180 14364
rect 54348 14308 54404 16604
rect 54460 16594 54516 16604
rect 54460 16324 54516 16334
rect 54460 15874 54516 16268
rect 54460 15822 54462 15874
rect 54514 15822 54516 15874
rect 54460 15428 54516 15822
rect 54460 15362 54516 15372
rect 54348 14242 54404 14252
rect 54460 14084 54516 14094
rect 54124 14028 54404 14084
rect 54124 13860 54180 13870
rect 54124 13858 54292 13860
rect 54124 13806 54126 13858
rect 54178 13806 54292 13858
rect 54124 13804 54292 13806
rect 54124 13794 54180 13804
rect 54236 13636 54292 13804
rect 54236 13570 54292 13580
rect 54012 13346 54068 13356
rect 54124 13524 54180 13534
rect 53900 13234 53956 13244
rect 53788 13076 53844 13086
rect 53788 13074 54068 13076
rect 53788 13022 53790 13074
rect 53842 13022 54068 13074
rect 53788 13020 54068 13022
rect 53788 13010 53844 13020
rect 53452 12758 53508 12796
rect 53788 12850 53844 12862
rect 53788 12798 53790 12850
rect 53842 12798 53844 12850
rect 53676 12740 53732 12750
rect 53676 12646 53732 12684
rect 53452 12404 53508 12414
rect 53340 12402 53508 12404
rect 53340 12350 53454 12402
rect 53506 12350 53508 12402
rect 53340 12348 53508 12350
rect 53004 12236 53172 12292
rect 53452 12292 53508 12348
rect 52780 10882 52836 10892
rect 52892 11284 52948 11294
rect 52780 10724 52836 10734
rect 52780 10630 52836 10668
rect 52892 10722 52948 11228
rect 52892 10670 52894 10722
rect 52946 10670 52948 10722
rect 52892 10658 52948 10670
rect 52668 9090 52724 9100
rect 52780 10386 52836 10398
rect 52780 10334 52782 10386
rect 52834 10334 52836 10386
rect 52780 9044 52836 10334
rect 53004 9604 53060 12236
rect 53452 12226 53508 12236
rect 53676 12292 53732 12302
rect 53228 12178 53284 12190
rect 53228 12126 53230 12178
rect 53282 12126 53284 12178
rect 53004 9538 53060 9548
rect 53116 11956 53172 11966
rect 52892 9044 52948 9054
rect 52780 9042 52948 9044
rect 52780 8990 52894 9042
rect 52946 8990 52948 9042
rect 52780 8988 52948 8990
rect 52668 8932 52724 8942
rect 52444 8930 52724 8932
rect 52444 8878 52670 8930
rect 52722 8878 52724 8930
rect 52444 8876 52724 8878
rect 52444 8260 52500 8876
rect 52668 8866 52724 8876
rect 52780 8708 52836 8988
rect 52892 8978 52948 8988
rect 52444 8128 52500 8204
rect 52556 8652 52836 8708
rect 52556 8146 52612 8652
rect 52556 8094 52558 8146
rect 52610 8094 52612 8146
rect 52556 8082 52612 8094
rect 53004 8260 53060 8270
rect 52780 8036 52836 8046
rect 52780 7586 52836 7980
rect 52780 7534 52782 7586
rect 52834 7534 52836 7586
rect 52780 7522 52836 7534
rect 52780 7362 52836 7374
rect 52780 7310 52782 7362
rect 52834 7310 52836 7362
rect 52556 6692 52612 6702
rect 52556 6598 52612 6636
rect 52332 6412 52612 6468
rect 52444 6132 52500 6142
rect 52220 6130 52500 6132
rect 52220 6078 52446 6130
rect 52498 6078 52500 6130
rect 52220 6076 52500 6078
rect 52444 6066 52500 6076
rect 52108 5182 52110 5234
rect 52162 5182 52164 5234
rect 52108 5170 52164 5182
rect 52444 5236 52500 5246
rect 52556 5236 52612 6412
rect 52444 5234 52612 5236
rect 52444 5182 52446 5234
rect 52498 5182 52612 5234
rect 52444 5180 52612 5182
rect 52444 5170 52500 5180
rect 50204 5068 50484 5124
rect 50204 5012 50260 5068
rect 50204 4946 50260 4956
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 52780 4564 52836 7310
rect 53004 7252 53060 8204
rect 53004 7186 53060 7196
rect 53004 6020 53060 6030
rect 53004 5926 53060 5964
rect 52780 4498 52836 4508
rect 50652 4452 50708 4462
rect 49868 3332 50036 3388
rect 50428 3668 50484 3678
rect 49868 2996 49924 3332
rect 49868 2930 49924 2940
rect 49084 2818 49140 2828
rect 50428 800 50484 3612
rect 50652 3554 50708 4396
rect 51324 3668 51380 3678
rect 51324 3574 51380 3612
rect 50652 3502 50654 3554
rect 50706 3502 50708 3554
rect 50652 3490 50708 3502
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 53116 2548 53172 11900
rect 53228 11284 53284 12126
rect 53564 12180 53620 12190
rect 53228 11218 53284 11228
rect 53452 12068 53508 12078
rect 53340 10724 53396 10734
rect 53340 10630 53396 10668
rect 53340 9828 53396 9838
rect 53340 9734 53396 9772
rect 53452 9604 53508 12012
rect 53564 11394 53620 12124
rect 53564 11342 53566 11394
rect 53618 11342 53620 11394
rect 53564 11330 53620 11342
rect 53676 11394 53732 12236
rect 53788 11620 53844 12798
rect 53788 11554 53844 11564
rect 53676 11342 53678 11394
rect 53730 11342 53732 11394
rect 53676 11330 53732 11342
rect 53788 11396 53844 11406
rect 53788 11302 53844 11340
rect 54012 11394 54068 13020
rect 54124 12402 54180 13468
rect 54236 12962 54292 12974
rect 54236 12910 54238 12962
rect 54290 12910 54292 12962
rect 54236 12852 54292 12910
rect 54236 12786 54292 12796
rect 54124 12350 54126 12402
rect 54178 12350 54180 12402
rect 54124 12338 54180 12350
rect 54236 12516 54292 12526
rect 54236 12292 54292 12460
rect 54236 12198 54292 12236
rect 54012 11342 54014 11394
rect 54066 11342 54068 11394
rect 53564 11172 53620 11182
rect 53564 10834 53620 11116
rect 53900 11172 53956 11182
rect 53900 11078 53956 11116
rect 54012 10948 54068 11342
rect 53564 10782 53566 10834
rect 53618 10782 53620 10834
rect 53564 10770 53620 10782
rect 53676 10892 54068 10948
rect 54124 11732 54180 11742
rect 53676 10722 53732 10892
rect 54124 10834 54180 11676
rect 54124 10782 54126 10834
rect 54178 10782 54180 10834
rect 54124 10770 54180 10782
rect 53676 10670 53678 10722
rect 53730 10670 53732 10722
rect 53676 10658 53732 10670
rect 54348 10500 54404 14028
rect 54460 13858 54516 14028
rect 54460 13806 54462 13858
rect 54514 13806 54516 13858
rect 54460 13794 54516 13806
rect 54460 13636 54516 13646
rect 54460 11620 54516 13580
rect 54460 11554 54516 11564
rect 54572 11618 54628 17052
rect 54684 16882 54740 17164
rect 54684 16830 54686 16882
rect 54738 16830 54740 16882
rect 54684 16818 54740 16830
rect 54796 16772 54852 18844
rect 54908 17668 54964 17678
rect 54908 17574 54964 17612
rect 54796 16706 54852 16716
rect 54908 17332 54964 17342
rect 54796 15874 54852 15886
rect 54796 15822 54798 15874
rect 54850 15822 54852 15874
rect 54796 15314 54852 15822
rect 54796 15262 54798 15314
rect 54850 15262 54852 15314
rect 54796 15092 54852 15262
rect 54684 14532 54740 14542
rect 54684 12852 54740 14476
rect 54796 14308 54852 15036
rect 54796 14242 54852 14252
rect 54684 12786 54740 12796
rect 54796 13412 54852 13422
rect 54684 12404 54740 12414
rect 54684 12310 54740 12348
rect 54572 11566 54574 11618
rect 54626 11566 54628 11618
rect 54572 11554 54628 11566
rect 54572 11172 54628 11182
rect 53900 10444 54404 10500
rect 54460 11170 54628 11172
rect 54460 11118 54574 11170
rect 54626 11118 54628 11170
rect 54460 11116 54628 11118
rect 53788 9940 53844 9950
rect 53788 9846 53844 9884
rect 53340 9548 53508 9604
rect 53340 8260 53396 9548
rect 53340 8194 53396 8204
rect 53452 9156 53508 9166
rect 53228 8036 53284 8046
rect 53228 7474 53284 7980
rect 53228 7422 53230 7474
rect 53282 7422 53284 7474
rect 53228 7410 53284 7422
rect 53340 7364 53396 7374
rect 53340 6130 53396 7308
rect 53452 6692 53508 9100
rect 53564 8932 53620 8942
rect 53564 8838 53620 8876
rect 53788 8372 53844 8382
rect 53788 8278 53844 8316
rect 53676 8260 53732 8270
rect 53564 8258 53732 8260
rect 53564 8206 53678 8258
rect 53730 8206 53732 8258
rect 53564 8204 53732 8206
rect 53564 7474 53620 8204
rect 53676 8194 53732 8204
rect 53564 7422 53566 7474
rect 53618 7422 53620 7474
rect 53564 6916 53620 7422
rect 53788 7924 53844 7934
rect 53788 7140 53844 7868
rect 53788 7074 53844 7084
rect 53564 6850 53620 6860
rect 53452 6560 53508 6636
rect 53788 6692 53844 6702
rect 53900 6692 53956 10444
rect 53788 6690 53956 6692
rect 53788 6638 53790 6690
rect 53842 6638 53956 6690
rect 53788 6636 53956 6638
rect 53788 6626 53844 6636
rect 53340 6078 53342 6130
rect 53394 6078 53396 6130
rect 53340 6066 53396 6078
rect 53788 6132 53844 6142
rect 53788 6038 53844 6076
rect 53900 5682 53956 6636
rect 54012 10276 54068 10286
rect 54012 6132 54068 10220
rect 54348 9716 54404 9726
rect 54348 9622 54404 9660
rect 54460 9268 54516 11116
rect 54572 11106 54628 11116
rect 54684 11060 54740 11070
rect 54572 10836 54628 10846
rect 54572 10742 54628 10780
rect 54572 10500 54628 10510
rect 54572 9716 54628 10444
rect 54684 9938 54740 11004
rect 54684 9886 54686 9938
rect 54738 9886 54740 9938
rect 54684 9874 54740 9886
rect 54796 9828 54852 13356
rect 54908 13300 54964 17276
rect 55020 15876 55076 19070
rect 55132 19124 55188 19134
rect 55132 18450 55188 19068
rect 55244 19122 55300 19292
rect 55356 19282 55412 19292
rect 55468 19236 55524 19246
rect 55468 19142 55524 19180
rect 55244 19070 55246 19122
rect 55298 19070 55300 19122
rect 55244 19058 55300 19070
rect 55356 19010 55412 19022
rect 55692 19012 55748 20748
rect 55356 18958 55358 19010
rect 55410 18958 55412 19010
rect 55132 18398 55134 18450
rect 55186 18398 55188 18450
rect 55132 18386 55188 18398
rect 55244 18900 55300 18910
rect 55132 16884 55188 16894
rect 55132 16790 55188 16828
rect 55020 15810 55076 15820
rect 55020 15652 55076 15662
rect 55020 15538 55076 15596
rect 55020 15486 55022 15538
rect 55074 15486 55076 15538
rect 55020 15474 55076 15486
rect 55244 15148 55300 18844
rect 55356 16994 55412 18958
rect 55468 18956 55748 19012
rect 55468 17108 55524 18956
rect 55692 18676 55748 18686
rect 55692 18450 55748 18620
rect 55692 18398 55694 18450
rect 55746 18398 55748 18450
rect 55692 18386 55748 18398
rect 55468 17042 55524 17052
rect 55356 16942 55358 16994
rect 55410 16942 55412 16994
rect 55356 16930 55412 16942
rect 55132 15092 55300 15148
rect 55356 16772 55412 16782
rect 55020 14532 55076 14542
rect 55020 14438 55076 14476
rect 55132 14420 55188 15092
rect 55356 14532 55412 16716
rect 55580 16658 55636 16670
rect 55580 16606 55582 16658
rect 55634 16606 55636 16658
rect 55580 16436 55636 16606
rect 55580 16370 55636 16380
rect 55692 16660 55748 16670
rect 55692 16210 55748 16604
rect 55692 16158 55694 16210
rect 55746 16158 55748 16210
rect 55692 16146 55748 16158
rect 55692 15988 55748 15998
rect 55580 15932 55692 15988
rect 55580 15148 55636 15932
rect 55692 15894 55748 15932
rect 55804 15876 55860 22316
rect 55916 21698 55972 24332
rect 56700 24050 56756 25452
rect 56700 23998 56702 24050
rect 56754 23998 56756 24050
rect 56700 23986 56756 23998
rect 56028 23826 56084 23838
rect 56028 23774 56030 23826
rect 56082 23774 56084 23826
rect 56028 23604 56084 23774
rect 56028 23538 56084 23548
rect 55916 21646 55918 21698
rect 55970 21646 55972 21698
rect 55916 18900 55972 21646
rect 56140 23380 56196 23390
rect 56028 21586 56084 21598
rect 56028 21534 56030 21586
rect 56082 21534 56084 21586
rect 56028 21028 56084 21534
rect 56028 20962 56084 20972
rect 56140 19236 56196 23324
rect 56476 23380 56532 23390
rect 56476 23154 56532 23324
rect 56476 23102 56478 23154
rect 56530 23102 56532 23154
rect 56476 23090 56532 23102
rect 56700 23042 56756 23054
rect 56700 22990 56702 23042
rect 56754 22990 56756 23042
rect 56700 22372 56756 22990
rect 56700 22306 56756 22316
rect 56812 22370 56868 25564
rect 56924 24164 56980 29596
rect 57148 25060 57204 31500
rect 57708 31556 57764 31566
rect 57708 31462 57764 31500
rect 57484 30882 57540 30894
rect 57484 30830 57486 30882
rect 57538 30830 57540 30882
rect 57484 30212 57540 30830
rect 57820 30884 57876 30894
rect 57820 30790 57876 30828
rect 57484 30156 57988 30212
rect 57372 29986 57428 29998
rect 57820 29988 57876 29998
rect 57372 29934 57374 29986
rect 57426 29934 57428 29986
rect 57372 29540 57428 29934
rect 57708 29986 57876 29988
rect 57708 29934 57822 29986
rect 57874 29934 57876 29986
rect 57708 29932 57876 29934
rect 57484 29540 57540 29550
rect 57428 29538 57540 29540
rect 57428 29486 57486 29538
rect 57538 29486 57540 29538
rect 57428 29484 57540 29486
rect 57372 29474 57428 29484
rect 57484 29474 57540 29484
rect 57596 28644 57652 28654
rect 57596 28550 57652 28588
rect 57260 28532 57316 28542
rect 57316 28476 57540 28532
rect 57260 28438 57316 28476
rect 57372 27972 57428 27982
rect 57372 27878 57428 27916
rect 57372 26852 57428 26862
rect 57372 26758 57428 26796
rect 57372 26404 57428 26414
rect 57372 26310 57428 26348
rect 57036 25004 57204 25060
rect 57484 25732 57540 28476
rect 57708 27074 57764 29932
rect 57820 29922 57876 29932
rect 57820 29540 57876 29550
rect 57932 29540 57988 30156
rect 57820 29538 57988 29540
rect 57820 29486 57822 29538
rect 57874 29486 57988 29538
rect 57820 29484 57988 29486
rect 57820 28420 57876 29484
rect 58044 28644 58100 28654
rect 58044 28550 58100 28588
rect 57820 28354 57876 28364
rect 57820 27748 57876 27758
rect 57820 27654 57876 27692
rect 57708 27022 57710 27074
rect 57762 27022 57764 27074
rect 57708 26628 57764 27022
rect 57708 26562 57764 26572
rect 57820 26178 57876 26190
rect 57820 26126 57822 26178
rect 57874 26126 57876 26178
rect 57596 25732 57652 25742
rect 57484 25730 57652 25732
rect 57484 25678 57598 25730
rect 57650 25678 57652 25730
rect 57484 25676 57652 25678
rect 57036 24500 57092 25004
rect 57484 24948 57540 25676
rect 57596 25666 57652 25676
rect 57708 25284 57764 25294
rect 57036 24434 57092 24444
rect 57148 24946 57540 24948
rect 57148 24894 57486 24946
rect 57538 24894 57540 24946
rect 57148 24892 57540 24894
rect 56924 24098 56980 24108
rect 57148 24162 57204 24892
rect 57484 24882 57540 24892
rect 57596 25282 57764 25284
rect 57596 25230 57710 25282
rect 57762 25230 57764 25282
rect 57596 25228 57764 25230
rect 57596 24724 57652 25228
rect 57708 25218 57764 25228
rect 57820 25172 57876 26126
rect 57820 25106 57876 25116
rect 57932 26066 57988 26078
rect 57932 26014 57934 26066
rect 57986 26014 57988 26066
rect 57932 25506 57988 26014
rect 57932 25454 57934 25506
rect 57986 25454 57988 25506
rect 57148 24110 57150 24162
rect 57202 24110 57204 24162
rect 57148 24098 57204 24110
rect 57260 24668 57652 24724
rect 56924 23938 56980 23950
rect 56924 23886 56926 23938
rect 56978 23886 56980 23938
rect 56924 23380 56980 23886
rect 56924 22484 56980 23324
rect 57036 22484 57092 22494
rect 56924 22482 57092 22484
rect 56924 22430 57038 22482
rect 57090 22430 57092 22482
rect 56924 22428 57092 22430
rect 57036 22418 57092 22428
rect 56812 22318 56814 22370
rect 56866 22318 56868 22370
rect 56812 22260 56868 22318
rect 56476 22146 56532 22158
rect 56476 22094 56478 22146
rect 56530 22094 56532 22146
rect 56476 21700 56532 22094
rect 56476 21634 56532 21644
rect 56588 21474 56644 21486
rect 56588 21422 56590 21474
rect 56642 21422 56644 21474
rect 56364 21364 56420 21374
rect 56364 20242 56420 21308
rect 56588 20356 56644 21422
rect 56588 20290 56644 20300
rect 56364 20190 56366 20242
rect 56418 20190 56420 20242
rect 56364 20178 56420 20190
rect 56252 19236 56308 19246
rect 56196 19234 56308 19236
rect 56196 19182 56254 19234
rect 56306 19182 56308 19234
rect 56196 19180 56308 19182
rect 56140 19104 56196 19180
rect 56252 19170 56308 19180
rect 55916 18844 56420 18900
rect 56252 18564 56308 18574
rect 56252 18470 56308 18508
rect 56028 18338 56084 18350
rect 56028 18286 56030 18338
rect 56082 18286 56084 18338
rect 55916 18228 55972 18238
rect 55916 17778 55972 18172
rect 55916 17726 55918 17778
rect 55970 17726 55972 17778
rect 55916 17714 55972 17726
rect 56028 17780 56084 18286
rect 56028 17714 56084 17724
rect 56364 16884 56420 18844
rect 56812 18788 56868 22204
rect 57260 21476 57316 24668
rect 57372 24500 57428 24510
rect 57372 21700 57428 24444
rect 57596 24164 57652 24174
rect 57596 24070 57652 24108
rect 57820 24052 57876 24062
rect 57820 23716 57876 23996
rect 57932 23940 57988 25454
rect 58044 25172 58100 25182
rect 58044 24722 58100 25116
rect 58044 24670 58046 24722
rect 58098 24670 58100 24722
rect 58044 24658 58100 24670
rect 57932 23884 58100 23940
rect 57932 23716 57988 23726
rect 57820 23714 57988 23716
rect 57820 23662 57934 23714
rect 57986 23662 57988 23714
rect 57820 23660 57988 23662
rect 57932 23650 57988 23660
rect 57484 23380 57540 23390
rect 57484 22260 57540 23324
rect 57932 23044 57988 23054
rect 57708 23042 57988 23044
rect 57708 22990 57934 23042
rect 57986 22990 57988 23042
rect 57708 22988 57988 22990
rect 57596 22260 57652 22270
rect 57484 22258 57652 22260
rect 57484 22206 57598 22258
rect 57650 22206 57652 22258
rect 57484 22204 57652 22206
rect 57596 22194 57652 22204
rect 57708 21924 57764 22988
rect 57932 22978 57988 22988
rect 58044 22820 58100 23884
rect 58156 22932 58212 48860
rect 58380 32452 58436 32462
rect 58268 30884 58324 30894
rect 58268 26066 58324 30828
rect 58268 26014 58270 26066
rect 58322 26014 58324 26066
rect 58268 26002 58324 26014
rect 58156 22866 58212 22876
rect 57372 21644 57652 21700
rect 57260 21420 57428 21476
rect 57260 21140 57316 21150
rect 57260 20802 57316 21084
rect 57260 20750 57262 20802
rect 57314 20750 57316 20802
rect 57260 19348 57316 20750
rect 57260 19282 57316 19292
rect 57148 19234 57204 19246
rect 57148 19182 57150 19234
rect 57202 19182 57204 19234
rect 56812 18732 56980 18788
rect 56476 18452 56532 18462
rect 56476 18358 56532 18396
rect 56588 18340 56644 18350
rect 56476 17444 56532 17454
rect 56476 16884 56532 17388
rect 56588 16996 56644 18284
rect 56812 17666 56868 17678
rect 56812 17614 56814 17666
rect 56866 17614 56868 17666
rect 56700 17556 56756 17566
rect 56700 17462 56756 17500
rect 56700 16996 56756 17006
rect 56588 16994 56756 16996
rect 56588 16942 56702 16994
rect 56754 16942 56756 16994
rect 56588 16940 56756 16942
rect 56700 16884 56756 16940
rect 56476 16828 56644 16884
rect 56364 16818 56420 16828
rect 56028 16658 56084 16670
rect 56028 16606 56030 16658
rect 56082 16606 56084 16658
rect 56028 16548 56084 16606
rect 56028 16482 56084 16492
rect 56252 16658 56308 16670
rect 56476 16660 56532 16670
rect 56252 16606 56254 16658
rect 56306 16606 56308 16658
rect 55916 16212 55972 16222
rect 56252 16212 56308 16606
rect 55916 16210 56308 16212
rect 55916 16158 55918 16210
rect 55970 16158 56308 16210
rect 55916 16156 56308 16158
rect 55916 16146 55972 16156
rect 56028 15876 56084 15886
rect 55804 15820 55972 15876
rect 55804 15316 55860 15326
rect 55132 14288 55188 14364
rect 55244 14476 55412 14532
rect 55468 15092 55636 15148
rect 55692 15204 55748 15242
rect 55804 15222 55860 15260
rect 55692 15138 55748 15148
rect 55132 14084 55188 14094
rect 55132 13970 55188 14028
rect 55132 13918 55134 13970
rect 55186 13918 55188 13970
rect 55132 13906 55188 13918
rect 55020 13746 55076 13758
rect 55020 13694 55022 13746
rect 55074 13694 55076 13746
rect 55020 13524 55076 13694
rect 55020 13458 55076 13468
rect 54908 13244 55188 13300
rect 54908 13076 54964 13086
rect 54908 12982 54964 13020
rect 54572 9660 54740 9716
rect 54460 9202 54516 9212
rect 54460 9042 54516 9054
rect 54460 8990 54462 9042
rect 54514 8990 54516 9042
rect 54348 8484 54404 8494
rect 54348 7698 54404 8428
rect 54460 7924 54516 8990
rect 54572 8260 54628 8270
rect 54572 8166 54628 8204
rect 54460 7858 54516 7868
rect 54348 7646 54350 7698
rect 54402 7646 54404 7698
rect 54348 7634 54404 7646
rect 54348 7140 54404 7150
rect 54236 6692 54292 6702
rect 54236 6598 54292 6636
rect 54012 6066 54068 6076
rect 54124 6580 54180 6590
rect 53900 5630 53902 5682
rect 53954 5630 53956 5682
rect 53900 5618 53956 5630
rect 54012 5908 54068 5918
rect 53900 5236 53956 5246
rect 54012 5236 54068 5852
rect 53900 5234 54068 5236
rect 53900 5182 53902 5234
rect 53954 5182 54068 5234
rect 53900 5180 54068 5182
rect 53900 5170 53956 5180
rect 53116 2482 53172 2492
rect 54124 1652 54180 6524
rect 54348 5236 54404 7084
rect 54460 6132 54516 6142
rect 54684 6132 54740 9660
rect 54796 6690 54852 9772
rect 54908 12852 54964 12862
rect 54908 11956 54964 12796
rect 55132 12402 55188 13244
rect 55132 12350 55134 12402
rect 55186 12350 55188 12402
rect 55132 12338 55188 12350
rect 54908 8148 54964 11900
rect 55020 11620 55076 11630
rect 55020 10500 55076 11564
rect 55132 11508 55188 11518
rect 55132 11414 55188 11452
rect 55132 10836 55188 10846
rect 55244 10836 55300 14476
rect 55356 14308 55412 14318
rect 55356 14214 55412 14252
rect 55468 14084 55524 15092
rect 55580 14418 55636 14430
rect 55580 14366 55582 14418
rect 55634 14366 55636 14418
rect 55580 14196 55636 14366
rect 55580 14130 55636 14140
rect 55468 14018 55524 14028
rect 55804 13972 55860 13982
rect 55916 13972 55972 15820
rect 55804 13970 55972 13972
rect 55804 13918 55806 13970
rect 55858 13918 55972 13970
rect 55804 13916 55972 13918
rect 56028 13972 56084 15820
rect 56252 15876 56308 16156
rect 56364 16658 56532 16660
rect 56364 16606 56478 16658
rect 56530 16606 56532 16658
rect 56364 16604 56532 16606
rect 56364 15988 56420 16604
rect 56476 16594 56532 16604
rect 56588 16436 56644 16828
rect 56700 16818 56756 16828
rect 56364 15922 56420 15932
rect 56476 16380 56644 16436
rect 56700 16660 56756 16670
rect 56252 15810 56308 15820
rect 56476 15874 56532 16380
rect 56700 15876 56756 16604
rect 56812 16098 56868 17614
rect 56812 16046 56814 16098
rect 56866 16046 56868 16098
rect 56812 15988 56868 16046
rect 56812 15922 56868 15932
rect 56476 15822 56478 15874
rect 56530 15822 56532 15874
rect 56364 15316 56420 15326
rect 56364 15222 56420 15260
rect 56476 15148 56532 15822
rect 56252 15092 56532 15148
rect 56588 15820 56756 15876
rect 56140 14420 56196 14430
rect 56140 14326 56196 14364
rect 56140 13972 56196 13982
rect 56028 13970 56196 13972
rect 56028 13918 56142 13970
rect 56194 13918 56196 13970
rect 56028 13916 56196 13918
rect 55804 13906 55860 13916
rect 56140 13906 56196 13916
rect 55356 13860 55412 13870
rect 55356 13766 55412 13804
rect 55580 13524 55636 13534
rect 55132 10834 55300 10836
rect 55132 10782 55134 10834
rect 55186 10782 55300 10834
rect 55132 10780 55300 10782
rect 55356 12292 55412 12302
rect 55132 10770 55188 10780
rect 55020 10434 55076 10444
rect 55244 9940 55300 9950
rect 55244 9846 55300 9884
rect 55020 9042 55076 9054
rect 55020 8990 55022 9042
rect 55074 8990 55076 9042
rect 55020 8932 55076 8990
rect 55020 8260 55076 8876
rect 55132 8932 55188 8942
rect 55132 8930 55300 8932
rect 55132 8878 55134 8930
rect 55186 8878 55300 8930
rect 55132 8876 55300 8878
rect 55132 8866 55188 8876
rect 55132 8260 55188 8270
rect 55020 8258 55188 8260
rect 55020 8206 55134 8258
rect 55186 8206 55188 8258
rect 55020 8204 55188 8206
rect 55132 8194 55188 8204
rect 55244 8260 55300 8876
rect 55244 8194 55300 8204
rect 54908 8092 55076 8148
rect 54796 6638 54798 6690
rect 54850 6638 54852 6690
rect 54796 6626 54852 6638
rect 54908 7252 54964 7262
rect 54908 6468 54964 7196
rect 54460 6130 54740 6132
rect 54460 6078 54462 6130
rect 54514 6078 54740 6130
rect 54460 6076 54740 6078
rect 54796 6412 54964 6468
rect 54460 6066 54516 6076
rect 54348 5104 54404 5180
rect 54796 5234 54852 6412
rect 54908 6020 54964 6030
rect 54908 5926 54964 5964
rect 54796 5182 54798 5234
rect 54850 5182 54852 5234
rect 54796 5170 54852 5182
rect 55020 5236 55076 8092
rect 55244 8034 55300 8046
rect 55244 7982 55246 8034
rect 55298 7982 55300 8034
rect 55244 7924 55300 7982
rect 55244 7858 55300 7868
rect 55356 7700 55412 12236
rect 55468 11618 55524 11630
rect 55468 11566 55470 11618
rect 55522 11566 55524 11618
rect 55468 9268 55524 11566
rect 55580 11506 55636 13468
rect 55804 13076 55860 13086
rect 55692 12068 55748 12106
rect 55692 12002 55748 12012
rect 55804 11788 55860 13020
rect 56140 12850 56196 12862
rect 56140 12798 56142 12850
rect 56194 12798 56196 12850
rect 56028 12404 56084 12414
rect 56028 12310 56084 12348
rect 55580 11454 55582 11506
rect 55634 11454 55636 11506
rect 55580 11442 55636 11454
rect 55692 11732 55860 11788
rect 56140 12180 56196 12798
rect 55692 10834 55748 11732
rect 55916 11618 55972 11630
rect 55916 11566 55918 11618
rect 55970 11566 55972 11618
rect 55916 11506 55972 11566
rect 55916 11454 55918 11506
rect 55970 11454 55972 11506
rect 55916 11442 55972 11454
rect 55692 10782 55694 10834
rect 55746 10782 55748 10834
rect 55692 10770 55748 10782
rect 56028 10500 56084 10510
rect 56028 10406 56084 10444
rect 55580 10052 55636 10062
rect 55580 9938 55636 9996
rect 55580 9886 55582 9938
rect 55634 9886 55636 9938
rect 55580 9874 55636 9886
rect 56028 9604 56084 9642
rect 56028 9538 56084 9548
rect 56028 9380 56084 9390
rect 55580 9268 55636 9278
rect 55468 9266 55636 9268
rect 55468 9214 55582 9266
rect 55634 9214 55636 9266
rect 55468 9212 55636 9214
rect 55468 8484 55524 9212
rect 55580 9202 55636 9212
rect 56028 9266 56084 9324
rect 56028 9214 56030 9266
rect 56082 9214 56084 9266
rect 56028 9202 56084 9214
rect 55468 8418 55524 8428
rect 55916 8260 55972 8270
rect 55468 8036 55524 8046
rect 55468 7942 55524 7980
rect 55804 8036 55860 8046
rect 55356 7644 55524 7700
rect 55356 7362 55412 7374
rect 55356 7310 55358 7362
rect 55410 7310 55412 7362
rect 55356 6804 55412 7310
rect 55356 6738 55412 6748
rect 55356 6580 55412 6590
rect 55356 6486 55412 6524
rect 55468 5908 55524 7644
rect 55804 7476 55860 7980
rect 55804 7410 55860 7420
rect 55916 6690 55972 8204
rect 55916 6638 55918 6690
rect 55970 6638 55972 6690
rect 55916 6626 55972 6638
rect 56028 8148 56084 8158
rect 56140 8148 56196 12124
rect 56252 8372 56308 15092
rect 56476 14308 56532 14318
rect 56588 14308 56644 15820
rect 56924 15764 56980 18732
rect 57148 18340 57204 19182
rect 57148 18274 57204 18284
rect 57372 18004 57428 21420
rect 57484 21474 57540 21486
rect 57484 21422 57486 21474
rect 57538 21422 57540 21474
rect 57484 21252 57540 21422
rect 57484 21186 57540 21196
rect 57596 20356 57652 21644
rect 57708 20690 57764 21868
rect 57820 22764 58100 22820
rect 57820 22372 57876 22764
rect 57820 21698 57876 22316
rect 57932 22372 57988 22382
rect 58380 22372 58436 32396
rect 59388 24612 59444 24622
rect 57932 22370 58436 22372
rect 57932 22318 57934 22370
rect 57986 22318 58436 22370
rect 57932 22316 58436 22318
rect 58604 22932 58660 22942
rect 57932 22306 57988 22316
rect 57820 21646 57822 21698
rect 57874 21646 57876 21698
rect 57820 21588 57876 21646
rect 57932 21588 57988 21598
rect 57820 21586 57988 21588
rect 57820 21534 57934 21586
rect 57986 21534 57988 21586
rect 57820 21532 57988 21534
rect 57932 21522 57988 21532
rect 58268 21588 58324 21598
rect 58268 21586 58436 21588
rect 58268 21534 58270 21586
rect 58322 21534 58436 21586
rect 58268 21532 58436 21534
rect 58268 21522 58324 21532
rect 57708 20638 57710 20690
rect 57762 20638 57764 20690
rect 57708 20626 57764 20638
rect 57596 20300 57876 20356
rect 57484 20244 57540 20254
rect 57484 20150 57540 20188
rect 57708 20018 57764 20030
rect 57708 19966 57710 20018
rect 57762 19966 57764 20018
rect 57484 18564 57540 18574
rect 57484 18470 57540 18508
rect 57708 18340 57764 19966
rect 57708 18274 57764 18284
rect 57820 18562 57876 20300
rect 57820 18510 57822 18562
rect 57874 18510 57876 18562
rect 57148 17948 57428 18004
rect 56812 15708 56980 15764
rect 57036 17556 57092 17566
rect 56476 14306 56644 14308
rect 56476 14254 56478 14306
rect 56530 14254 56644 14306
rect 56476 14252 56644 14254
rect 56700 15428 56756 15438
rect 56364 13860 56420 13870
rect 56364 11618 56420 13804
rect 56476 13748 56532 14252
rect 56700 14196 56756 15372
rect 56700 14130 56756 14140
rect 56476 13682 56532 13692
rect 56588 13636 56644 13646
rect 56588 13524 56644 13580
rect 56364 11566 56366 11618
rect 56418 11566 56420 11618
rect 56364 11554 56420 11566
rect 56476 13468 56644 13524
rect 56476 11508 56532 13468
rect 56812 12964 56868 15708
rect 57036 15652 57092 17500
rect 57148 16548 57204 17948
rect 57260 17668 57316 17678
rect 57820 17668 57876 18510
rect 57932 19796 57988 19806
rect 57932 17778 57988 19740
rect 58044 19122 58100 19134
rect 58044 19070 58046 19122
rect 58098 19070 58100 19122
rect 58044 18340 58100 19070
rect 58044 18116 58100 18284
rect 58044 18050 58100 18060
rect 58268 18788 58324 18798
rect 57932 17726 57934 17778
rect 57986 17726 57988 17778
rect 57932 17714 57988 17726
rect 57260 17666 57876 17668
rect 57260 17614 57262 17666
rect 57314 17614 57876 17666
rect 57260 17612 57876 17614
rect 57260 17602 57316 17612
rect 57484 17108 57540 17612
rect 57484 17106 57652 17108
rect 57484 17054 57486 17106
rect 57538 17054 57652 17106
rect 57484 17052 57652 17054
rect 57484 17042 57540 17052
rect 57148 16482 57204 16492
rect 57372 15988 57428 15998
rect 57372 15894 57428 15932
rect 56812 12898 56868 12908
rect 56924 15596 57092 15652
rect 57260 15652 57316 15662
rect 56812 12738 56868 12750
rect 56812 12686 56814 12738
rect 56866 12686 56868 12738
rect 56812 12628 56868 12686
rect 56812 12562 56868 12572
rect 56588 12404 56644 12414
rect 56924 12404 56980 15596
rect 57036 14308 57092 14318
rect 57036 14214 57092 14252
rect 57260 13972 57316 15596
rect 57484 15316 57540 15326
rect 57372 14532 57428 14542
rect 57484 14532 57540 15260
rect 57372 14530 57540 14532
rect 57372 14478 57374 14530
rect 57426 14478 57540 14530
rect 57372 14476 57540 14478
rect 57372 14466 57428 14476
rect 57484 14196 57540 14206
rect 57372 13972 57428 13982
rect 57260 13970 57428 13972
rect 57260 13918 57374 13970
rect 57426 13918 57428 13970
rect 57260 13916 57428 13918
rect 57372 13906 57428 13916
rect 57372 13748 57428 13758
rect 57260 13076 57316 13086
rect 57260 12982 57316 13020
rect 56588 12402 56980 12404
rect 56588 12350 56590 12402
rect 56642 12350 56980 12402
rect 56588 12348 56980 12350
rect 57036 12964 57092 12974
rect 56588 12338 56644 12348
rect 57036 12068 57092 12908
rect 57036 12002 57092 12012
rect 57148 12516 57204 12526
rect 56476 11442 56532 11452
rect 56812 11618 56868 11630
rect 56812 11566 56814 11618
rect 56866 11566 56868 11618
rect 56812 11506 56868 11566
rect 56812 11454 56814 11506
rect 56866 11454 56868 11506
rect 56812 11442 56868 11454
rect 56364 11170 56420 11182
rect 56364 11118 56366 11170
rect 56418 11118 56420 11170
rect 56364 10612 56420 11118
rect 56476 10948 56532 10958
rect 56476 10834 56532 10892
rect 56476 10782 56478 10834
rect 56530 10782 56532 10834
rect 56476 10770 56532 10782
rect 57036 10836 57092 10846
rect 57148 10836 57204 12460
rect 57372 12402 57428 13692
rect 57372 12350 57374 12402
rect 57426 12350 57428 12402
rect 57372 12338 57428 12350
rect 57372 11508 57428 11518
rect 57372 11414 57428 11452
rect 57372 10836 57428 10846
rect 57148 10834 57428 10836
rect 57148 10782 57374 10834
rect 57426 10782 57428 10834
rect 57148 10780 57428 10782
rect 56364 10546 56420 10556
rect 57036 9938 57092 10780
rect 57372 10386 57428 10780
rect 57372 10334 57374 10386
rect 57426 10334 57428 10386
rect 57372 10322 57428 10334
rect 57036 9886 57038 9938
rect 57090 9886 57092 9938
rect 57036 9874 57092 9886
rect 57372 10052 57428 10062
rect 57372 9938 57428 9996
rect 57372 9886 57374 9938
rect 57426 9886 57428 9938
rect 57372 9716 57428 9886
rect 57372 9650 57428 9660
rect 56476 9604 56532 9614
rect 56532 9548 56644 9604
rect 56476 9472 56532 9548
rect 56476 9268 56532 9278
rect 56476 9174 56532 9212
rect 56364 8372 56420 8382
rect 56252 8370 56420 8372
rect 56252 8318 56366 8370
rect 56418 8318 56420 8370
rect 56252 8316 56420 8318
rect 56364 8306 56420 8316
rect 56140 8092 56420 8148
rect 55916 6132 55972 6142
rect 56028 6132 56084 8092
rect 56140 7474 56196 7486
rect 56140 7422 56142 7474
rect 56194 7422 56196 7474
rect 56140 6580 56196 7422
rect 56252 6580 56308 6590
rect 56140 6578 56308 6580
rect 56140 6526 56254 6578
rect 56306 6526 56308 6578
rect 56140 6524 56308 6526
rect 56252 6514 56308 6524
rect 55916 6130 56084 6132
rect 55916 6078 55918 6130
rect 55970 6078 56084 6130
rect 55916 6076 56084 6078
rect 55916 6066 55972 6076
rect 55468 5842 55524 5852
rect 55244 5794 55300 5806
rect 55244 5742 55246 5794
rect 55298 5742 55300 5794
rect 55244 5682 55300 5742
rect 55244 5630 55246 5682
rect 55298 5630 55300 5682
rect 55244 5618 55300 5630
rect 56028 5682 56084 6076
rect 56364 6130 56420 8092
rect 56588 8036 56644 9548
rect 57372 9268 57428 9278
rect 57484 9268 57540 14140
rect 57372 9266 57540 9268
rect 57372 9214 57374 9266
rect 57426 9214 57540 9266
rect 57372 9212 57540 9214
rect 57372 9202 57428 9212
rect 57484 8372 57540 8382
rect 57484 8278 57540 8316
rect 56924 8036 56980 8046
rect 56588 8034 56980 8036
rect 56588 7982 56926 8034
rect 56978 7982 56980 8034
rect 56588 7980 56980 7982
rect 56812 7700 56868 7710
rect 56812 7606 56868 7644
rect 56812 6692 56868 6702
rect 56812 6598 56868 6636
rect 56364 6078 56366 6130
rect 56418 6078 56420 6130
rect 56364 6066 56420 6078
rect 56028 5630 56030 5682
rect 56082 5630 56084 5682
rect 56028 5618 56084 5630
rect 56812 5794 56868 5806
rect 56812 5742 56814 5794
rect 56866 5742 56868 5794
rect 56812 5682 56868 5742
rect 56812 5630 56814 5682
rect 56866 5630 56868 5682
rect 56812 5618 56868 5630
rect 55244 5236 55300 5246
rect 55020 5234 55300 5236
rect 55020 5182 55246 5234
rect 55298 5182 55300 5234
rect 55020 5180 55300 5182
rect 55244 5170 55300 5180
rect 55580 5236 55636 5246
rect 55580 5142 55636 5180
rect 56924 5012 56980 7980
rect 57596 7700 57652 17052
rect 57708 16884 57764 16894
rect 57708 16660 57764 16828
rect 57820 16884 57876 16894
rect 57820 16882 58100 16884
rect 57820 16830 57822 16882
rect 57874 16830 58100 16882
rect 57820 16828 58100 16830
rect 57820 16818 57876 16828
rect 57708 16604 57876 16660
rect 57708 15986 57764 15998
rect 57708 15934 57710 15986
rect 57762 15934 57764 15986
rect 57708 13860 57764 15934
rect 57820 15538 57876 16604
rect 57820 15486 57822 15538
rect 57874 15486 57876 15538
rect 57820 15474 57876 15486
rect 58044 14644 58100 16828
rect 58044 14550 58100 14588
rect 57932 14306 57988 14318
rect 57932 14254 57934 14306
rect 57986 14254 57988 14306
rect 57932 14084 57988 14254
rect 57932 14018 57988 14028
rect 57708 13794 57764 13804
rect 58044 13860 58100 13870
rect 57820 13636 57876 13646
rect 57708 13634 57876 13636
rect 57708 13582 57822 13634
rect 57874 13582 57876 13634
rect 57708 13580 57876 13582
rect 57708 12740 57764 13580
rect 57820 13570 57876 13580
rect 57708 12646 57764 12684
rect 57932 12628 57988 12638
rect 57820 12068 57876 12078
rect 57820 11974 57876 12012
rect 57708 11844 57764 11854
rect 57708 11620 57764 11788
rect 57932 11620 57988 12572
rect 58044 12292 58100 13804
rect 58044 12226 58100 12236
rect 58156 12404 58212 12414
rect 57708 11564 57876 11620
rect 57708 11170 57764 11182
rect 57708 11118 57710 11170
rect 57762 11118 57764 11170
rect 57708 9940 57764 11118
rect 57820 10836 57876 11564
rect 57932 11554 57988 11564
rect 57820 10704 57876 10780
rect 57708 9874 57764 9884
rect 57932 10386 57988 10398
rect 57932 10334 57934 10386
rect 57986 10334 57988 10386
rect 57932 9268 57988 10334
rect 58044 9828 58100 9838
rect 58044 9734 58100 9772
rect 58044 9268 58100 9278
rect 57932 9266 58100 9268
rect 57932 9214 58046 9266
rect 58098 9214 58100 9266
rect 57932 9212 58100 9214
rect 57932 8148 57988 9212
rect 58044 9202 58100 9212
rect 57932 8082 57988 8092
rect 58044 8372 58100 8382
rect 58156 8372 58212 12348
rect 58268 9380 58324 18732
rect 58380 11508 58436 21532
rect 58380 11442 58436 11452
rect 58492 18340 58548 18350
rect 58492 10052 58548 18284
rect 58492 9986 58548 9996
rect 58268 9314 58324 9324
rect 58044 8370 58212 8372
rect 58044 8318 58046 8370
rect 58098 8318 58212 8370
rect 58044 8316 58212 8318
rect 58044 7700 58100 8316
rect 57596 7698 57876 7700
rect 57596 7646 57598 7698
rect 57650 7646 57876 7698
rect 57596 7644 57876 7646
rect 57596 7634 57652 7644
rect 57148 7028 57204 7038
rect 57148 6466 57204 6972
rect 57820 6802 57876 7644
rect 58044 7568 58100 7644
rect 57820 6750 57822 6802
rect 57874 6750 57876 6802
rect 57820 6738 57876 6750
rect 57148 6414 57150 6466
rect 57202 6414 57204 6466
rect 57148 6132 57204 6414
rect 57932 6132 57988 6142
rect 57148 6130 57988 6132
rect 57148 6078 57934 6130
rect 57986 6078 57988 6130
rect 57148 6076 57988 6078
rect 57932 6066 57988 6076
rect 57372 5908 57428 5918
rect 57372 5814 57428 5852
rect 56924 4946 56980 4956
rect 54236 4900 54292 4910
rect 54236 4564 54292 4844
rect 54348 4564 54404 4574
rect 54236 4562 54404 4564
rect 54236 4510 54350 4562
rect 54402 4510 54404 4562
rect 54236 4508 54404 4510
rect 54348 4340 54404 4508
rect 55916 4452 55972 4462
rect 54348 4274 54404 4284
rect 54908 4340 54964 4350
rect 54908 4246 54964 4284
rect 55804 4226 55860 4238
rect 55804 4174 55806 4226
rect 55858 4174 55860 4226
rect 54124 1586 54180 1596
rect 55244 3666 55300 3678
rect 55244 3614 55246 3666
rect 55298 3614 55300 3666
rect 55244 1428 55300 3614
rect 55244 1362 55300 1372
rect 55804 800 55860 4174
rect 55916 3554 55972 4396
rect 57484 4452 57540 4462
rect 57484 4358 57540 4396
rect 55916 3502 55918 3554
rect 55970 3502 55972 3554
rect 55916 3490 55972 3502
rect 56700 4340 56756 4350
rect 56700 2772 56756 4284
rect 57708 4340 57764 4350
rect 57708 4246 57764 4284
rect 58604 4228 58660 22876
rect 58828 18564 58884 18574
rect 58716 16996 58772 17006
rect 58716 8036 58772 16940
rect 58828 8372 58884 18508
rect 58940 16884 58996 16894
rect 58940 12404 58996 16828
rect 59388 13188 59444 24556
rect 59388 13122 59444 13132
rect 58940 12338 58996 12348
rect 58828 8306 58884 8316
rect 58716 7970 58772 7980
rect 58604 4162 58660 4172
rect 56700 2706 56756 2716
rect 0 200 112 800
rect 5376 200 5488 800
rect 10752 200 10864 800
rect 16800 200 16912 800
rect 22176 200 22288 800
rect 27552 200 27664 800
rect 33600 200 33712 800
rect 38976 200 39088 800
rect 44352 200 44464 800
rect 50400 200 50512 800
rect 55776 200 55888 800
<< via2 >>
rect 2604 58380 2660 58436
rect 1372 58044 1428 58100
rect 2268 58044 2324 58100
rect 1260 55916 1316 55972
rect 1148 52220 1204 52276
rect 1148 47180 1204 47236
rect 1932 55804 1988 55860
rect 1820 53618 1876 53620
rect 1820 53566 1822 53618
rect 1822 53566 1874 53618
rect 1874 53566 1876 53618
rect 1820 53564 1876 53566
rect 2492 54402 2548 54404
rect 2492 54350 2494 54402
rect 2494 54350 2546 54402
rect 2546 54350 2548 54402
rect 2492 54348 2548 54350
rect 2268 53506 2324 53508
rect 2268 53454 2270 53506
rect 2270 53454 2322 53506
rect 2322 53454 2324 53506
rect 2268 53452 2324 53454
rect 2044 53340 2100 53396
rect 1484 53228 1540 53284
rect 1372 52780 1428 52836
rect 2492 53116 2548 53172
rect 2156 52834 2212 52836
rect 2156 52782 2158 52834
rect 2158 52782 2210 52834
rect 2210 52782 2212 52834
rect 2156 52780 2212 52782
rect 1820 52556 1876 52612
rect 1932 51938 1988 51940
rect 1932 51886 1934 51938
rect 1934 51886 1986 51938
rect 1986 51886 1988 51938
rect 1932 51884 1988 51886
rect 1932 50482 1988 50484
rect 1932 50430 1934 50482
rect 1934 50430 1986 50482
rect 1986 50430 1988 50482
rect 1932 50428 1988 50430
rect 2156 51884 2212 51940
rect 1820 48914 1876 48916
rect 1820 48862 1822 48914
rect 1822 48862 1874 48914
rect 1874 48862 1876 48914
rect 1820 48860 1876 48862
rect 2044 48860 2100 48916
rect 1484 48412 1540 48468
rect 1596 48300 1652 48356
rect 1372 42924 1428 42980
rect 1484 47180 1540 47236
rect 1596 44492 1652 44548
rect 1708 47068 1764 47124
rect 2268 50764 2324 50820
rect 2380 50652 2436 50708
rect 2156 48076 2212 48132
rect 4620 57372 4676 57428
rect 6636 57260 6692 57316
rect 5852 57148 5908 57204
rect 3052 55970 3108 55972
rect 3052 55918 3054 55970
rect 3054 55918 3106 55970
rect 3106 55918 3108 55970
rect 3052 55916 3108 55918
rect 2828 55298 2884 55300
rect 2828 55246 2830 55298
rect 2830 55246 2882 55298
rect 2882 55246 2884 55298
rect 2828 55244 2884 55246
rect 5068 55970 5124 55972
rect 5068 55918 5070 55970
rect 5070 55918 5122 55970
rect 5122 55918 5124 55970
rect 5068 55916 5124 55918
rect 5404 55916 5460 55972
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 4172 55244 4228 55300
rect 5180 55580 5236 55636
rect 5068 55186 5124 55188
rect 5068 55134 5070 55186
rect 5070 55134 5122 55186
rect 5122 55134 5124 55186
rect 5068 55132 5124 55134
rect 3724 54460 3780 54516
rect 3948 54684 4004 54740
rect 2716 53228 2772 53284
rect 2940 52556 2996 52612
rect 2604 52220 2660 52276
rect 2716 51996 2772 52052
rect 2716 49026 2772 49028
rect 2716 48974 2718 49026
rect 2718 48974 2770 49026
rect 2770 48974 2772 49026
rect 2716 48972 2772 48974
rect 2828 49084 2884 49140
rect 2044 47458 2100 47460
rect 2044 47406 2046 47458
rect 2046 47406 2098 47458
rect 2098 47406 2100 47458
rect 2044 47404 2100 47406
rect 2156 47516 2212 47572
rect 1932 46002 1988 46004
rect 1932 45950 1934 46002
rect 1934 45950 1986 46002
rect 1986 45950 1988 46002
rect 1932 45948 1988 45950
rect 1932 44380 1988 44436
rect 2044 44940 2100 44996
rect 1820 43372 1876 43428
rect 1932 43260 1988 43316
rect 2268 46844 2324 46900
rect 2492 46956 2548 47012
rect 2604 46844 2660 46900
rect 2604 46172 2660 46228
rect 3388 53788 3444 53844
rect 3164 52780 3220 52836
rect 3276 52162 3332 52164
rect 3276 52110 3278 52162
rect 3278 52110 3330 52162
rect 3330 52110 3332 52162
rect 3276 52108 3332 52110
rect 3052 51212 3108 51268
rect 3052 50594 3108 50596
rect 3052 50542 3054 50594
rect 3054 50542 3106 50594
rect 3106 50542 3108 50594
rect 3052 50540 3108 50542
rect 3164 50428 3220 50484
rect 3164 49644 3220 49700
rect 3836 54402 3892 54404
rect 3836 54350 3838 54402
rect 3838 54350 3890 54402
rect 3890 54350 3892 54402
rect 3836 54348 3892 54350
rect 3500 53676 3556 53732
rect 3500 53228 3556 53284
rect 3612 53116 3668 53172
rect 3388 49532 3444 49588
rect 3276 49196 3332 49252
rect 3052 48802 3108 48804
rect 3052 48750 3054 48802
rect 3054 48750 3106 48802
rect 3106 48750 3108 48802
rect 3052 48748 3108 48750
rect 2828 47852 2884 47908
rect 3052 47628 3108 47684
rect 3164 47458 3220 47460
rect 3164 47406 3166 47458
rect 3166 47406 3218 47458
rect 3218 47406 3220 47458
rect 3164 47404 3220 47406
rect 2828 46898 2884 46900
rect 2828 46846 2830 46898
rect 2830 46846 2882 46898
rect 2882 46846 2884 46898
rect 2828 46844 2884 46846
rect 3052 47234 3108 47236
rect 3052 47182 3054 47234
rect 3054 47182 3106 47234
rect 3106 47182 3108 47234
rect 3052 47180 3108 47182
rect 3612 50876 3668 50932
rect 3500 47852 3556 47908
rect 3612 50316 3668 50372
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 5068 54012 5124 54068
rect 4284 53004 4340 53060
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4060 51436 4116 51492
rect 4172 51548 4228 51604
rect 3948 50988 4004 51044
rect 3724 49980 3780 50036
rect 4172 50316 4228 50372
rect 4844 51490 4900 51492
rect 4844 51438 4846 51490
rect 4846 51438 4898 51490
rect 4898 51438 4900 51490
rect 4844 51436 4900 51438
rect 5180 53452 5236 53508
rect 5516 55692 5572 55748
rect 5964 56140 6020 56196
rect 5516 54012 5572 54068
rect 5628 53788 5684 53844
rect 5740 53730 5796 53732
rect 5740 53678 5742 53730
rect 5742 53678 5794 53730
rect 5794 53678 5796 53730
rect 5740 53676 5796 53678
rect 6076 55970 6132 55972
rect 6076 55918 6078 55970
rect 6078 55918 6130 55970
rect 6130 55918 6132 55970
rect 6076 55916 6132 55918
rect 6524 55970 6580 55972
rect 6524 55918 6526 55970
rect 6526 55918 6578 55970
rect 6578 55918 6580 55970
rect 6524 55916 6580 55918
rect 6300 54796 6356 54852
rect 6076 53676 6132 53732
rect 5628 53170 5684 53172
rect 5628 53118 5630 53170
rect 5630 53118 5682 53170
rect 5682 53118 5684 53170
rect 5628 53116 5684 53118
rect 5180 52220 5236 52276
rect 4956 51212 5012 51268
rect 5068 51996 5124 52052
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 5068 50988 5124 51044
rect 4396 50428 4452 50484
rect 4508 50370 4564 50372
rect 4508 50318 4510 50370
rect 4510 50318 4562 50370
rect 4562 50318 4564 50370
rect 4508 50316 4564 50318
rect 4284 50204 4340 50260
rect 3948 49980 4004 50036
rect 3948 49756 4004 49812
rect 3724 48748 3780 48804
rect 2940 46620 2996 46676
rect 3052 46732 3108 46788
rect 2716 45388 2772 45444
rect 2828 45106 2884 45108
rect 2828 45054 2830 45106
rect 2830 45054 2882 45106
rect 2882 45054 2884 45106
rect 2828 45052 2884 45054
rect 2492 44492 2548 44548
rect 2940 44322 2996 44324
rect 2940 44270 2942 44322
rect 2942 44270 2994 44322
rect 2994 44270 2996 44322
rect 2940 44268 2996 44270
rect 3500 46396 3556 46452
rect 3612 46844 3668 46900
rect 4060 49644 4116 49700
rect 4060 49420 4116 49476
rect 5068 50428 5124 50484
rect 4956 49756 5012 49812
rect 4620 49532 4676 49588
rect 3948 48018 4004 48020
rect 3948 47966 3950 48018
rect 3950 47966 4002 48018
rect 4002 47966 4004 48018
rect 3948 47964 4004 47966
rect 3836 46674 3892 46676
rect 3836 46622 3838 46674
rect 3838 46622 3890 46674
rect 3890 46622 3892 46674
rect 3836 46620 3892 46622
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4844 48972 4900 49028
rect 4732 48914 4788 48916
rect 4732 48862 4734 48914
rect 4734 48862 4786 48914
rect 4786 48862 4788 48914
rect 4732 48860 4788 48862
rect 4620 48748 4676 48804
rect 5068 48636 5124 48692
rect 4284 48412 4340 48468
rect 4844 48466 4900 48468
rect 4844 48414 4846 48466
rect 4846 48414 4898 48466
rect 4898 48414 4900 48466
rect 4844 48412 4900 48414
rect 4284 48188 4340 48244
rect 5068 48242 5124 48244
rect 5068 48190 5070 48242
rect 5070 48190 5122 48242
rect 5122 48190 5124 48242
rect 5068 48188 5124 48190
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4508 47570 4564 47572
rect 4508 47518 4510 47570
rect 4510 47518 4562 47570
rect 4562 47518 4564 47570
rect 4508 47516 4564 47518
rect 4732 47404 4788 47460
rect 4284 46786 4340 46788
rect 4284 46734 4286 46786
rect 4286 46734 4338 46786
rect 4338 46734 4340 46786
rect 4284 46732 4340 46734
rect 3724 46284 3780 46340
rect 3948 46172 4004 46228
rect 4172 46450 4228 46452
rect 4172 46398 4174 46450
rect 4174 46398 4226 46450
rect 4226 46398 4228 46450
rect 4172 46396 4228 46398
rect 3388 45890 3444 45892
rect 3388 45838 3390 45890
rect 3390 45838 3442 45890
rect 3442 45838 3444 45890
rect 3388 45836 3444 45838
rect 3612 45836 3668 45892
rect 3836 46060 3892 46116
rect 4060 45724 4116 45780
rect 2716 43708 2772 43764
rect 2268 43484 2324 43540
rect 2268 42700 2324 42756
rect 2156 42642 2212 42644
rect 2156 42590 2158 42642
rect 2158 42590 2210 42642
rect 2210 42590 2212 42642
rect 2156 42588 2212 42590
rect 2156 42364 2212 42420
rect 1932 41692 1988 41748
rect 1820 40908 1876 40964
rect 1820 40626 1876 40628
rect 1820 40574 1822 40626
rect 1822 40574 1874 40626
rect 1874 40574 1876 40626
rect 1820 40572 1876 40574
rect 2380 41858 2436 41860
rect 2380 41806 2382 41858
rect 2382 41806 2434 41858
rect 2434 41806 2436 41858
rect 2380 41804 2436 41806
rect 2604 42866 2660 42868
rect 2604 42814 2606 42866
rect 2606 42814 2658 42866
rect 2658 42814 2660 42866
rect 2604 42812 2660 42814
rect 2828 43650 2884 43652
rect 2828 43598 2830 43650
rect 2830 43598 2882 43650
rect 2882 43598 2884 43650
rect 2828 43596 2884 43598
rect 2940 43484 2996 43540
rect 2828 42588 2884 42644
rect 2828 42194 2884 42196
rect 2828 42142 2830 42194
rect 2830 42142 2882 42194
rect 2882 42142 2884 42194
rect 2828 42140 2884 42142
rect 2380 40236 2436 40292
rect 2492 40460 2548 40516
rect 1484 35868 1540 35924
rect 1596 39564 1652 39620
rect 1932 39004 1988 39060
rect 1820 38892 1876 38948
rect 1932 38834 1988 38836
rect 1932 38782 1934 38834
rect 1934 38782 1986 38834
rect 1986 38782 1988 38834
rect 1932 38780 1988 38782
rect 1708 37324 1764 37380
rect 1932 36652 1988 36708
rect 1820 36594 1876 36596
rect 1820 36542 1822 36594
rect 1822 36542 1874 36594
rect 1874 36542 1876 36594
rect 1820 36540 1876 36542
rect 1820 34636 1876 34692
rect 1932 33628 1988 33684
rect 1932 33458 1988 33460
rect 1932 33406 1934 33458
rect 1934 33406 1986 33458
rect 1986 33406 1988 33458
rect 1932 33404 1988 33406
rect 2156 38444 2212 38500
rect 2380 37938 2436 37940
rect 2380 37886 2382 37938
rect 2382 37886 2434 37938
rect 2434 37886 2436 37938
rect 2380 37884 2436 37886
rect 2604 39004 2660 39060
rect 3164 43932 3220 43988
rect 3276 45052 3332 45108
rect 3276 44156 3332 44212
rect 3276 43036 3332 43092
rect 3164 42082 3220 42084
rect 3164 42030 3166 42082
rect 3166 42030 3218 42082
rect 3218 42030 3220 42082
rect 3164 42028 3220 42030
rect 3052 40962 3108 40964
rect 3052 40910 3054 40962
rect 3054 40910 3106 40962
rect 3106 40910 3108 40962
rect 3052 40908 3108 40910
rect 2940 39676 2996 39732
rect 2828 39618 2884 39620
rect 2828 39566 2830 39618
rect 2830 39566 2882 39618
rect 2882 39566 2884 39618
rect 2828 39564 2884 39566
rect 2716 38444 2772 38500
rect 2716 37324 2772 37380
rect 2380 36370 2436 36372
rect 2380 36318 2382 36370
rect 2382 36318 2434 36370
rect 2434 36318 2436 36370
rect 2380 36316 2436 36318
rect 2268 35922 2324 35924
rect 2268 35870 2270 35922
rect 2270 35870 2322 35922
rect 2322 35870 2324 35922
rect 2268 35868 2324 35870
rect 2156 34914 2212 34916
rect 2156 34862 2158 34914
rect 2158 34862 2210 34914
rect 2210 34862 2212 34914
rect 2156 34860 2212 34862
rect 2380 33852 2436 33908
rect 2492 36092 2548 36148
rect 2380 33628 2436 33684
rect 2940 36370 2996 36372
rect 2940 36318 2942 36370
rect 2942 36318 2994 36370
rect 2994 36318 2996 36370
rect 2940 36316 2996 36318
rect 3164 39116 3220 39172
rect 3052 36092 3108 36148
rect 3164 38834 3220 38836
rect 3164 38782 3166 38834
rect 3166 38782 3218 38834
rect 3218 38782 3220 38834
rect 3164 38780 3220 38782
rect 3388 41244 3444 41300
rect 3948 45106 4004 45108
rect 3948 45054 3950 45106
rect 3950 45054 4002 45106
rect 4002 45054 4004 45106
rect 3948 45052 4004 45054
rect 3948 44268 4004 44324
rect 3724 43260 3780 43316
rect 3612 43148 3668 43204
rect 3612 42754 3668 42756
rect 3612 42702 3614 42754
rect 3614 42702 3666 42754
rect 3666 42702 3668 42754
rect 3612 42700 3668 42702
rect 3836 42866 3892 42868
rect 3836 42814 3838 42866
rect 3838 42814 3890 42866
rect 3890 42814 3892 42866
rect 3836 42812 3892 42814
rect 3724 42588 3780 42644
rect 3836 42252 3892 42308
rect 3276 38162 3332 38164
rect 3276 38110 3278 38162
rect 3278 38110 3330 38162
rect 3330 38110 3332 38162
rect 3276 38108 3332 38110
rect 3724 41244 3780 41300
rect 3276 37266 3332 37268
rect 3276 37214 3278 37266
rect 3278 37214 3330 37266
rect 3330 37214 3332 37266
rect 3276 37212 3332 37214
rect 3276 36370 3332 36372
rect 3276 36318 3278 36370
rect 3278 36318 3330 36370
rect 3330 36318 3332 36370
rect 3276 36316 3332 36318
rect 2716 35084 2772 35140
rect 2940 35196 2996 35252
rect 2604 34690 2660 34692
rect 2604 34638 2606 34690
rect 2606 34638 2658 34690
rect 2658 34638 2660 34690
rect 2604 34636 2660 34638
rect 1932 31276 1988 31332
rect 2044 31218 2100 31220
rect 2044 31166 2046 31218
rect 2046 31166 2098 31218
rect 2098 31166 2100 31218
rect 2044 31164 2100 31166
rect 2268 31276 2324 31332
rect 2380 31052 2436 31108
rect 2492 32956 2548 33012
rect 2940 33740 2996 33796
rect 3164 35084 3220 35140
rect 3164 33628 3220 33684
rect 3276 33404 3332 33460
rect 3276 33180 3332 33236
rect 3052 32956 3108 33012
rect 2940 32508 2996 32564
rect 3052 31836 3108 31892
rect 2716 31612 2772 31668
rect 3724 40572 3780 40628
rect 3836 41132 3892 41188
rect 5964 52892 6020 52948
rect 5852 52274 5908 52276
rect 5852 52222 5854 52274
rect 5854 52222 5906 52274
rect 5906 52222 5908 52274
rect 5852 52220 5908 52222
rect 5628 51884 5684 51940
rect 5292 51772 5348 51828
rect 5628 51660 5684 51716
rect 5404 51548 5460 51604
rect 5292 51100 5348 51156
rect 5740 51602 5796 51604
rect 5740 51550 5742 51602
rect 5742 51550 5794 51602
rect 5794 51550 5796 51602
rect 5740 51548 5796 51550
rect 5852 51436 5908 51492
rect 5964 50482 6020 50484
rect 5964 50430 5966 50482
rect 5966 50430 6018 50482
rect 6018 50430 6020 50482
rect 5964 50428 6020 50430
rect 6188 53170 6244 53172
rect 6188 53118 6190 53170
rect 6190 53118 6242 53170
rect 6242 53118 6244 53170
rect 6188 53116 6244 53118
rect 6300 52780 6356 52836
rect 6524 54124 6580 54180
rect 6524 53564 6580 53620
rect 10892 58156 10948 58212
rect 7532 57932 7588 57988
rect 7420 57820 7476 57876
rect 6860 55244 6916 55300
rect 6748 55074 6804 55076
rect 6748 55022 6750 55074
rect 6750 55022 6802 55074
rect 6802 55022 6804 55074
rect 6748 55020 6804 55022
rect 6748 53618 6804 53620
rect 6748 53566 6750 53618
rect 6750 53566 6802 53618
rect 6802 53566 6804 53618
rect 6748 53564 6804 53566
rect 6524 52220 6580 52276
rect 6636 51996 6692 52052
rect 6524 51884 6580 51940
rect 6412 50764 6468 50820
rect 9324 57596 9380 57652
rect 7868 57484 7924 57540
rect 6972 53900 7028 53956
rect 7756 53676 7812 53732
rect 7644 53618 7700 53620
rect 7644 53566 7646 53618
rect 7646 53566 7698 53618
rect 7698 53566 7700 53618
rect 7644 53564 7700 53566
rect 6972 52892 7028 52948
rect 7196 52946 7252 52948
rect 7196 52894 7198 52946
rect 7198 52894 7250 52946
rect 7250 52894 7252 52946
rect 7196 52892 7252 52894
rect 7196 52444 7252 52500
rect 6972 52220 7028 52276
rect 5852 50370 5908 50372
rect 5852 50318 5854 50370
rect 5854 50318 5906 50370
rect 5906 50318 5908 50370
rect 5852 50316 5908 50318
rect 5628 49868 5684 49924
rect 5404 48300 5460 48356
rect 5404 47964 5460 48020
rect 4844 46956 4900 47012
rect 4956 46844 5012 46900
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4620 46060 4676 46116
rect 4284 45948 4340 46004
rect 4508 46002 4564 46004
rect 4508 45950 4510 46002
rect 4510 45950 4562 46002
rect 4562 45950 4564 46002
rect 4508 45948 4564 45950
rect 4172 45500 4228 45556
rect 4396 45890 4452 45892
rect 4396 45838 4398 45890
rect 4398 45838 4450 45890
rect 4450 45838 4452 45890
rect 4396 45836 4452 45838
rect 4508 45276 4564 45332
rect 5068 46562 5124 46564
rect 5068 46510 5070 46562
rect 5070 46510 5122 46562
rect 5122 46510 5124 46562
rect 5068 46508 5124 46510
rect 5404 46956 5460 47012
rect 5292 46060 5348 46116
rect 5404 45724 5460 45780
rect 4172 44828 4228 44884
rect 4844 44828 4900 44884
rect 4172 43538 4228 43540
rect 4172 43486 4174 43538
rect 4174 43486 4226 43538
rect 4226 43486 4228 43538
rect 4172 43484 4228 43486
rect 4172 41916 4228 41972
rect 4060 41074 4116 41076
rect 4060 41022 4062 41074
rect 4062 41022 4114 41074
rect 4114 41022 4116 41074
rect 4060 41020 4116 41022
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4508 44492 4564 44548
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4844 43148 4900 43204
rect 4844 42082 4900 42084
rect 4844 42030 4846 42082
rect 4846 42030 4898 42082
rect 4898 42030 4900 42082
rect 4844 42028 4900 42030
rect 4620 41916 4676 41972
rect 4732 41804 4788 41860
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4620 41186 4676 41188
rect 4620 41134 4622 41186
rect 4622 41134 4674 41186
rect 4674 41134 4676 41186
rect 4620 41132 4676 41134
rect 5292 43708 5348 43764
rect 4956 41244 5012 41300
rect 5068 41692 5124 41748
rect 4732 41020 4788 41076
rect 4284 40684 4340 40740
rect 4508 40908 4564 40964
rect 3500 39618 3556 39620
rect 3500 39566 3502 39618
rect 3502 39566 3554 39618
rect 3554 39566 3556 39618
rect 3500 39564 3556 39566
rect 3500 37324 3556 37380
rect 3724 39788 3780 39844
rect 3836 39676 3892 39732
rect 4284 40236 4340 40292
rect 3948 39564 4004 39620
rect 4172 39676 4228 39732
rect 3836 39116 3892 39172
rect 3836 38946 3892 38948
rect 3836 38894 3838 38946
rect 3838 38894 3890 38946
rect 3890 38894 3892 38946
rect 3836 38892 3892 38894
rect 4172 39004 4228 39060
rect 4956 41074 5012 41076
rect 4956 41022 4958 41074
rect 4958 41022 5010 41074
rect 5010 41022 5012 41074
rect 4956 41020 5012 41022
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4844 40012 4900 40068
rect 4956 40684 5012 40740
rect 4684 39956 4740 39958
rect 4284 38780 4340 38836
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 3948 37826 4004 37828
rect 3948 37774 3950 37826
rect 3950 37774 4002 37826
rect 4002 37774 4004 37826
rect 3948 37772 4004 37774
rect 4956 39228 5012 39284
rect 5180 39676 5236 39732
rect 5180 39452 5236 39508
rect 5180 38722 5236 38724
rect 5180 38670 5182 38722
rect 5182 38670 5234 38722
rect 5234 38670 5236 38722
rect 5180 38668 5236 38670
rect 5180 38444 5236 38500
rect 4956 37772 5012 37828
rect 5180 37772 5236 37828
rect 4060 36706 4116 36708
rect 4060 36654 4062 36706
rect 4062 36654 4114 36706
rect 4114 36654 4116 36706
rect 4060 36652 4116 36654
rect 4508 37266 4564 37268
rect 4508 37214 4510 37266
rect 4510 37214 4562 37266
rect 4562 37214 4564 37266
rect 4508 37212 4564 37214
rect 4172 36316 4228 36372
rect 3948 36204 4004 36260
rect 3500 34972 3556 35028
rect 3612 34300 3668 34356
rect 3948 33964 4004 34020
rect 4172 34076 4228 34132
rect 3612 33292 3668 33348
rect 4060 33404 4116 33460
rect 3276 32562 3332 32564
rect 3276 32510 3278 32562
rect 3278 32510 3330 32562
rect 3330 32510 3332 32562
rect 3276 32508 3332 32510
rect 3388 32450 3444 32452
rect 3388 32398 3390 32450
rect 3390 32398 3442 32450
rect 3442 32398 3444 32450
rect 3388 32396 3444 32398
rect 2492 30940 2548 30996
rect 1932 30210 1988 30212
rect 1932 30158 1934 30210
rect 1934 30158 1986 30210
rect 1986 30158 1988 30210
rect 1932 30156 1988 30158
rect 1708 29596 1764 29652
rect 1596 29372 1652 29428
rect 2044 29260 2100 29316
rect 1260 28140 1316 28196
rect 1932 27580 1988 27636
rect 1932 22258 1988 22260
rect 1932 22206 1934 22258
rect 1934 22206 1986 22258
rect 1986 22206 1988 22258
rect 1932 22204 1988 22206
rect 2940 31052 2996 31108
rect 2828 30828 2884 30884
rect 2716 29932 2772 29988
rect 2156 28418 2212 28420
rect 2156 28366 2158 28418
rect 2158 28366 2210 28418
rect 2210 28366 2212 28418
rect 2156 28364 2212 28366
rect 2604 28754 2660 28756
rect 2604 28702 2606 28754
rect 2606 28702 2658 28754
rect 2658 28702 2660 28754
rect 2604 28700 2660 28702
rect 2380 28028 2436 28084
rect 3164 31218 3220 31220
rect 3164 31166 3166 31218
rect 3166 31166 3218 31218
rect 3218 31166 3220 31218
rect 3164 31164 3220 31166
rect 3276 29986 3332 29988
rect 3276 29934 3278 29986
rect 3278 29934 3330 29986
rect 3330 29934 3332 29986
rect 3276 29932 3332 29934
rect 3276 29650 3332 29652
rect 3276 29598 3278 29650
rect 3278 29598 3330 29650
rect 3330 29598 3332 29650
rect 3276 29596 3332 29598
rect 3612 32620 3668 32676
rect 3612 32396 3668 32452
rect 3612 31666 3668 31668
rect 3612 31614 3614 31666
rect 3614 31614 3666 31666
rect 3666 31614 3668 31666
rect 3612 31612 3668 31614
rect 3724 30156 3780 30212
rect 3612 29596 3668 29652
rect 3948 32508 4004 32564
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4508 36316 4564 36372
rect 4732 35922 4788 35924
rect 4732 35870 4734 35922
rect 4734 35870 4786 35922
rect 4786 35870 4788 35922
rect 4732 35868 4788 35870
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4844 35308 4900 35364
rect 4956 37212 5012 37268
rect 4684 35252 4740 35254
rect 5068 35196 5124 35252
rect 4732 34914 4788 34916
rect 4732 34862 4734 34914
rect 4734 34862 4786 34914
rect 4786 34862 4788 34914
rect 4732 34860 4788 34862
rect 4396 34354 4452 34356
rect 4396 34302 4398 34354
rect 4398 34302 4450 34354
rect 4450 34302 4452 34354
rect 4396 34300 4452 34302
rect 4956 34524 5012 34580
rect 5628 49308 5684 49364
rect 5628 47292 5684 47348
rect 5628 47068 5684 47124
rect 5516 45612 5572 45668
rect 5628 46732 5684 46788
rect 5964 49138 6020 49140
rect 5964 49086 5966 49138
rect 5966 49086 6018 49138
rect 6018 49086 6020 49138
rect 5964 49084 6020 49086
rect 5740 46620 5796 46676
rect 5964 46284 6020 46340
rect 5740 45388 5796 45444
rect 5628 44044 5684 44100
rect 5516 43426 5572 43428
rect 5516 43374 5518 43426
rect 5518 43374 5570 43426
rect 5570 43374 5572 43426
rect 5516 43372 5572 43374
rect 5404 42924 5460 42980
rect 5516 42082 5572 42084
rect 5516 42030 5518 42082
rect 5518 42030 5570 42082
rect 5570 42030 5572 42082
rect 5516 42028 5572 42030
rect 5292 36092 5348 36148
rect 5516 41804 5572 41860
rect 5180 34412 5236 34468
rect 6188 49196 6244 49252
rect 6412 48354 6468 48356
rect 6412 48302 6414 48354
rect 6414 48302 6466 48354
rect 6466 48302 6468 48354
rect 6412 48300 6468 48302
rect 6412 47404 6468 47460
rect 6636 48412 6692 48468
rect 6636 48242 6692 48244
rect 6636 48190 6638 48242
rect 6638 48190 6690 48242
rect 6690 48190 6692 48242
rect 6636 48188 6692 48190
rect 6636 47068 6692 47124
rect 6076 45052 6132 45108
rect 6188 46060 6244 46116
rect 5964 44716 6020 44772
rect 5964 44098 6020 44100
rect 5964 44046 5966 44098
rect 5966 44046 6018 44098
rect 6018 44046 6020 44098
rect 5964 44044 6020 44046
rect 5852 43708 5908 43764
rect 6524 46786 6580 46788
rect 6524 46734 6526 46786
rect 6526 46734 6578 46786
rect 6578 46734 6580 46786
rect 6524 46732 6580 46734
rect 6412 46674 6468 46676
rect 6412 46622 6414 46674
rect 6414 46622 6466 46674
rect 6466 46622 6468 46674
rect 6412 46620 6468 46622
rect 6636 46396 6692 46452
rect 6860 51660 6916 51716
rect 7532 52108 7588 52164
rect 7644 51884 7700 51940
rect 7756 52780 7812 52836
rect 7308 51548 7364 51604
rect 7420 51436 7476 51492
rect 7084 50370 7140 50372
rect 7084 50318 7086 50370
rect 7086 50318 7138 50370
rect 7138 50318 7140 50370
rect 7084 50316 7140 50318
rect 6860 49868 6916 49924
rect 7084 49810 7140 49812
rect 7084 49758 7086 49810
rect 7086 49758 7138 49810
rect 7138 49758 7140 49810
rect 7084 49756 7140 49758
rect 6972 49420 7028 49476
rect 6860 49196 6916 49252
rect 6860 48524 6916 48580
rect 7084 48972 7140 49028
rect 6972 48300 7028 48356
rect 7420 50428 7476 50484
rect 7644 50988 7700 51044
rect 7532 50316 7588 50372
rect 7532 49810 7588 49812
rect 7532 49758 7534 49810
rect 7534 49758 7586 49810
rect 7586 49758 7588 49810
rect 7532 49756 7588 49758
rect 7644 49196 7700 49252
rect 7644 49026 7700 49028
rect 7644 48974 7646 49026
rect 7646 48974 7698 49026
rect 7698 48974 7700 49026
rect 7644 48972 7700 48974
rect 9212 56252 9268 56308
rect 8988 55804 9044 55860
rect 7980 54012 8036 54068
rect 7980 53506 8036 53508
rect 7980 53454 7982 53506
rect 7982 53454 8034 53506
rect 8034 53454 8036 53506
rect 7980 53452 8036 53454
rect 8540 54684 8596 54740
rect 8652 54908 8708 54964
rect 8876 54796 8932 54852
rect 8092 53116 8148 53172
rect 8204 54348 8260 54404
rect 8428 53788 8484 53844
rect 9100 54348 9156 54404
rect 9100 53842 9156 53844
rect 9100 53790 9102 53842
rect 9102 53790 9154 53842
rect 9154 53790 9156 53842
rect 9100 53788 9156 53790
rect 8204 52892 8260 52948
rect 8204 52332 8260 52388
rect 8092 52108 8148 52164
rect 7980 51490 8036 51492
rect 7980 51438 7982 51490
rect 7982 51438 8034 51490
rect 8034 51438 8036 51490
rect 7980 51436 8036 51438
rect 8204 51996 8260 52052
rect 8876 53452 8932 53508
rect 8540 52668 8596 52724
rect 9100 52108 9156 52164
rect 8316 51324 8372 51380
rect 10444 56028 10500 56084
rect 10220 55970 10276 55972
rect 10220 55918 10222 55970
rect 10222 55918 10274 55970
rect 10274 55918 10276 55970
rect 10220 55916 10276 55918
rect 9772 55468 9828 55524
rect 10668 56028 10724 56084
rect 10668 55692 10724 55748
rect 9436 55186 9492 55188
rect 9436 55134 9438 55186
rect 9438 55134 9490 55186
rect 9490 55134 9492 55186
rect 9436 55132 9492 55134
rect 9884 55132 9940 55188
rect 9772 54908 9828 54964
rect 9772 54348 9828 54404
rect 9436 53954 9492 53956
rect 9436 53902 9438 53954
rect 9438 53902 9490 53954
rect 9490 53902 9492 53954
rect 9436 53900 9492 53902
rect 9884 54012 9940 54068
rect 10108 55020 10164 55076
rect 10332 54626 10388 54628
rect 10332 54574 10334 54626
rect 10334 54574 10386 54626
rect 10386 54574 10388 54626
rect 10332 54572 10388 54574
rect 10220 52780 10276 52836
rect 9996 52556 10052 52612
rect 9996 51772 10052 51828
rect 9212 51660 9268 51716
rect 9884 51602 9940 51604
rect 9884 51550 9886 51602
rect 9886 51550 9938 51602
rect 9938 51550 9940 51602
rect 9884 51548 9940 51550
rect 7980 51100 8036 51156
rect 7420 48354 7476 48356
rect 7420 48302 7422 48354
rect 7422 48302 7474 48354
rect 7474 48302 7476 48354
rect 7420 48300 7476 48302
rect 6860 47404 6916 47460
rect 8204 50764 8260 50820
rect 8092 50428 8148 50484
rect 7980 49138 8036 49140
rect 7980 49086 7982 49138
rect 7982 49086 8034 49138
rect 8034 49086 8036 49138
rect 7980 49084 8036 49086
rect 8204 49196 8260 49252
rect 7980 47852 8036 47908
rect 7980 47404 8036 47460
rect 7308 47292 7364 47348
rect 6300 45276 6356 45332
rect 6412 46172 6468 46228
rect 6300 44604 6356 44660
rect 5740 41692 5796 41748
rect 5852 43484 5908 43540
rect 6076 43426 6132 43428
rect 6076 43374 6078 43426
rect 6078 43374 6130 43426
rect 6130 43374 6132 43426
rect 6076 43372 6132 43374
rect 5964 41804 6020 41860
rect 6860 46172 6916 46228
rect 6972 45666 7028 45668
rect 6972 45614 6974 45666
rect 6974 45614 7026 45666
rect 7026 45614 7028 45666
rect 6972 45612 7028 45614
rect 6748 45500 6804 45556
rect 6636 44268 6692 44324
rect 6748 45164 6804 45220
rect 6972 45218 7028 45220
rect 6972 45166 6974 45218
rect 6974 45166 7026 45218
rect 7026 45166 7028 45218
rect 6972 45164 7028 45166
rect 6860 45106 6916 45108
rect 6860 45054 6862 45106
rect 6862 45054 6914 45106
rect 6914 45054 6916 45106
rect 6860 45052 6916 45054
rect 7420 46508 7476 46564
rect 7196 45500 7252 45556
rect 7308 45612 7364 45668
rect 6860 44604 6916 44660
rect 6860 44434 6916 44436
rect 6860 44382 6862 44434
rect 6862 44382 6914 44434
rect 6914 44382 6916 44434
rect 6860 44380 6916 44382
rect 6972 43932 7028 43988
rect 6748 43820 6804 43876
rect 6524 42924 6580 42980
rect 6748 42924 6804 42980
rect 6412 42812 6468 42868
rect 6748 42754 6804 42756
rect 6748 42702 6750 42754
rect 6750 42702 6802 42754
rect 6802 42702 6804 42754
rect 6748 42700 6804 42702
rect 6300 41970 6356 41972
rect 6300 41918 6302 41970
rect 6302 41918 6354 41970
rect 6354 41918 6356 41970
rect 6300 41916 6356 41918
rect 6188 41804 6244 41860
rect 6076 41468 6132 41524
rect 5964 41298 6020 41300
rect 5964 41246 5966 41298
rect 5966 41246 6018 41298
rect 6018 41246 6020 41298
rect 5964 41244 6020 41246
rect 5740 38834 5796 38836
rect 5740 38782 5742 38834
rect 5742 38782 5794 38834
rect 5794 38782 5796 38834
rect 5740 38780 5796 38782
rect 6636 42642 6692 42644
rect 6636 42590 6638 42642
rect 6638 42590 6690 42642
rect 6690 42590 6692 42642
rect 6636 42588 6692 42590
rect 6524 41580 6580 41636
rect 6860 41244 6916 41300
rect 6412 40460 6468 40516
rect 6636 41132 6692 41188
rect 5964 38332 6020 38388
rect 6076 38556 6132 38612
rect 5740 37884 5796 37940
rect 5852 37826 5908 37828
rect 5852 37774 5854 37826
rect 5854 37774 5906 37826
rect 5906 37774 5908 37826
rect 5852 37772 5908 37774
rect 6076 36876 6132 36932
rect 6076 36594 6132 36596
rect 6076 36542 6078 36594
rect 6078 36542 6130 36594
rect 6130 36542 6132 36594
rect 6076 36540 6132 36542
rect 6412 36428 6468 36484
rect 6300 36316 6356 36372
rect 6524 35756 6580 35812
rect 4956 34354 5012 34356
rect 4956 34302 4958 34354
rect 4958 34302 5010 34354
rect 5010 34302 5012 34354
rect 4956 34300 5012 34302
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4620 33458 4676 33460
rect 4620 33406 4622 33458
rect 4622 33406 4674 33458
rect 4674 33406 4676 33458
rect 4620 33404 4676 33406
rect 4284 32562 4340 32564
rect 4284 32510 4286 32562
rect 4286 32510 4338 32562
rect 4338 32510 4340 32562
rect 4284 32508 4340 32510
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4956 33404 5012 33460
rect 5628 35420 5684 35476
rect 5516 35196 5572 35252
rect 5852 34860 5908 34916
rect 5516 34412 5572 34468
rect 5740 34636 5796 34692
rect 5404 34354 5460 34356
rect 5404 34302 5406 34354
rect 5406 34302 5458 34354
rect 5458 34302 5460 34354
rect 5404 34300 5460 34302
rect 5516 34188 5572 34244
rect 5404 32562 5460 32564
rect 5404 32510 5406 32562
rect 5406 32510 5458 32562
rect 5458 32510 5460 32562
rect 5404 32508 5460 32510
rect 5180 31948 5236 32004
rect 4956 31666 5012 31668
rect 4956 31614 4958 31666
rect 4958 31614 5010 31666
rect 5010 31614 5012 31666
rect 4956 31612 5012 31614
rect 4956 31388 5012 31444
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4172 30156 4228 30212
rect 4284 29708 4340 29764
rect 3724 29372 3780 29428
rect 4844 29596 4900 29652
rect 5068 30994 5124 30996
rect 5068 30942 5070 30994
rect 5070 30942 5122 30994
rect 5122 30942 5124 30994
rect 5068 30940 5124 30942
rect 5068 29932 5124 29988
rect 3276 28588 3332 28644
rect 3052 28028 3108 28084
rect 3500 28082 3556 28084
rect 3500 28030 3502 28082
rect 3502 28030 3554 28082
rect 3554 28030 3556 28082
rect 3500 28028 3556 28030
rect 3276 25116 3332 25172
rect 2940 24892 2996 24948
rect 2716 20524 2772 20580
rect 3276 20578 3332 20580
rect 3276 20526 3278 20578
rect 3278 20526 3330 20578
rect 3330 20526 3332 20578
rect 3276 20524 3332 20526
rect 1932 16828 1988 16884
rect 1932 10780 1988 10836
rect 2716 17052 2772 17108
rect 3276 17106 3332 17108
rect 3276 17054 3278 17106
rect 3278 17054 3330 17106
rect 3330 17054 3332 17106
rect 3276 17052 3332 17054
rect 2716 12402 2772 12404
rect 2716 12350 2718 12402
rect 2718 12350 2770 12402
rect 2770 12350 2772 12402
rect 2716 12348 2772 12350
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4508 28642 4564 28644
rect 4508 28590 4510 28642
rect 4510 28590 4562 28642
rect 4562 28590 4564 28642
rect 4508 28588 4564 28590
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 5180 29538 5236 29540
rect 5180 29486 5182 29538
rect 5182 29486 5234 29538
rect 5234 29486 5236 29538
rect 5180 29484 5236 29486
rect 6188 34914 6244 34916
rect 6188 34862 6190 34914
rect 6190 34862 6242 34914
rect 6242 34862 6244 34914
rect 6188 34860 6244 34862
rect 6188 34412 6244 34468
rect 5852 33234 5908 33236
rect 5852 33182 5854 33234
rect 5854 33182 5906 33234
rect 5906 33182 5908 33234
rect 5852 33180 5908 33182
rect 5628 32172 5684 32228
rect 5516 30940 5572 30996
rect 5180 28700 5236 28756
rect 6076 32844 6132 32900
rect 5964 32508 6020 32564
rect 5964 31612 6020 31668
rect 5628 29708 5684 29764
rect 6300 34354 6356 34356
rect 6300 34302 6302 34354
rect 6302 34302 6354 34354
rect 6354 34302 6356 34354
rect 6300 34300 6356 34302
rect 6860 40908 6916 40964
rect 6860 39788 6916 39844
rect 6748 39676 6804 39732
rect 7084 41804 7140 41860
rect 7420 45500 7476 45556
rect 7532 45276 7588 45332
rect 7532 45106 7588 45108
rect 7532 45054 7534 45106
rect 7534 45054 7586 45106
rect 7586 45054 7588 45106
rect 7532 45052 7588 45054
rect 7532 44716 7588 44772
rect 8092 47292 8148 47348
rect 8092 46898 8148 46900
rect 8092 46846 8094 46898
rect 8094 46846 8146 46898
rect 8146 46846 8148 46898
rect 8092 46844 8148 46846
rect 8092 46450 8148 46452
rect 8092 46398 8094 46450
rect 8094 46398 8146 46450
rect 8146 46398 8148 46450
rect 8092 46396 8148 46398
rect 7980 45948 8036 46004
rect 7868 45612 7924 45668
rect 8316 48972 8372 49028
rect 8428 47404 8484 47460
rect 8876 51212 8932 51268
rect 9660 50876 9716 50932
rect 8652 50204 8708 50260
rect 8652 49644 8708 49700
rect 9436 50316 9492 50372
rect 9100 49644 9156 49700
rect 9324 49868 9380 49924
rect 8652 49420 8708 49476
rect 8988 49138 9044 49140
rect 8988 49086 8990 49138
rect 8990 49086 9042 49138
rect 9042 49086 9044 49138
rect 8988 49084 9044 49086
rect 8652 48188 8708 48244
rect 8764 48076 8820 48132
rect 8540 46060 8596 46116
rect 8428 45890 8484 45892
rect 8428 45838 8430 45890
rect 8430 45838 8482 45890
rect 8482 45838 8484 45890
rect 8428 45836 8484 45838
rect 8204 45218 8260 45220
rect 8204 45166 8206 45218
rect 8206 45166 8258 45218
rect 8258 45166 8260 45218
rect 8204 45164 8260 45166
rect 7756 44716 7812 44772
rect 8204 44716 8260 44772
rect 7980 44380 8036 44436
rect 7532 44044 7588 44100
rect 7420 43538 7476 43540
rect 7420 43486 7422 43538
rect 7422 43486 7474 43538
rect 7474 43486 7476 43538
rect 7420 43484 7476 43486
rect 7308 42588 7364 42644
rect 7420 42082 7476 42084
rect 7420 42030 7422 42082
rect 7422 42030 7474 42082
rect 7474 42030 7476 42082
rect 7420 42028 7476 42030
rect 7308 41132 7364 41188
rect 7084 40514 7140 40516
rect 7084 40462 7086 40514
rect 7086 40462 7138 40514
rect 7138 40462 7140 40514
rect 7084 40460 7140 40462
rect 7196 40290 7252 40292
rect 7196 40238 7198 40290
rect 7198 40238 7250 40290
rect 7250 40238 7252 40290
rect 7196 40236 7252 40238
rect 7308 40178 7364 40180
rect 7308 40126 7310 40178
rect 7310 40126 7362 40178
rect 7362 40126 7364 40178
rect 7308 40124 7364 40126
rect 7644 43932 7700 43988
rect 7868 43932 7924 43988
rect 8092 43820 8148 43876
rect 8092 43596 8148 43652
rect 7868 43484 7924 43540
rect 7756 43372 7812 43428
rect 7756 42252 7812 42308
rect 7644 41132 7700 41188
rect 7756 42028 7812 42084
rect 7532 41020 7588 41076
rect 7980 41298 8036 41300
rect 7980 41246 7982 41298
rect 7982 41246 8034 41298
rect 8034 41246 8036 41298
rect 7980 41244 8036 41246
rect 7084 39564 7140 39620
rect 7084 39004 7140 39060
rect 7084 38050 7140 38052
rect 7084 37998 7086 38050
rect 7086 37998 7138 38050
rect 7138 37998 7140 38050
rect 7084 37996 7140 37998
rect 8876 47628 8932 47684
rect 9212 47628 9268 47684
rect 8988 47346 9044 47348
rect 8988 47294 8990 47346
rect 8990 47294 9042 47346
rect 9042 47294 9044 47346
rect 8988 47292 9044 47294
rect 9212 47292 9268 47348
rect 8876 46898 8932 46900
rect 8876 46846 8878 46898
rect 8878 46846 8930 46898
rect 8930 46846 8932 46898
rect 8876 46844 8932 46846
rect 8652 45836 8708 45892
rect 8988 45890 9044 45892
rect 8988 45838 8990 45890
rect 8990 45838 9042 45890
rect 9042 45838 9044 45890
rect 8988 45836 9044 45838
rect 8652 45612 8708 45668
rect 8652 45106 8708 45108
rect 8652 45054 8654 45106
rect 8654 45054 8706 45106
rect 8706 45054 8708 45106
rect 8652 45052 8708 45054
rect 8428 44604 8484 44660
rect 8428 44322 8484 44324
rect 8428 44270 8430 44322
rect 8430 44270 8482 44322
rect 8482 44270 8484 44322
rect 8428 44268 8484 44270
rect 8540 43650 8596 43652
rect 8540 43598 8542 43650
rect 8542 43598 8594 43650
rect 8594 43598 8596 43650
rect 8540 43596 8596 43598
rect 8316 43372 8372 43428
rect 8316 42476 8372 42532
rect 8428 43260 8484 43316
rect 8540 42530 8596 42532
rect 8540 42478 8542 42530
rect 8542 42478 8594 42530
rect 8594 42478 8596 42530
rect 8540 42476 8596 42478
rect 8204 42140 8260 42196
rect 8428 41468 8484 41524
rect 8428 40684 8484 40740
rect 9212 45388 9268 45444
rect 9212 45052 9268 45108
rect 8988 44156 9044 44212
rect 8988 43820 9044 43876
rect 8988 43426 9044 43428
rect 8988 43374 8990 43426
rect 8990 43374 9042 43426
rect 9042 43374 9044 43426
rect 8988 43372 9044 43374
rect 8988 41804 9044 41860
rect 9212 44044 9268 44100
rect 9212 43372 9268 43428
rect 9772 49980 9828 50036
rect 9436 49196 9492 49252
rect 9548 49644 9604 49700
rect 9436 47458 9492 47460
rect 9436 47406 9438 47458
rect 9438 47406 9490 47458
rect 9490 47406 9492 47458
rect 9436 47404 9492 47406
rect 9548 47068 9604 47124
rect 9772 48300 9828 48356
rect 9660 46898 9716 46900
rect 9660 46846 9662 46898
rect 9662 46846 9714 46898
rect 9714 46846 9716 46898
rect 9660 46844 9716 46846
rect 10108 51266 10164 51268
rect 10108 51214 10110 51266
rect 10110 51214 10162 51266
rect 10162 51214 10164 51266
rect 10108 51212 10164 51214
rect 10108 50428 10164 50484
rect 10444 51378 10500 51380
rect 10444 51326 10446 51378
rect 10446 51326 10498 51378
rect 10498 51326 10500 51378
rect 10444 51324 10500 51326
rect 10556 54012 10612 54068
rect 10780 53788 10836 53844
rect 11116 55970 11172 55972
rect 11116 55918 11118 55970
rect 11118 55918 11170 55970
rect 11170 55918 11172 55970
rect 11116 55916 11172 55918
rect 13356 58380 13412 58436
rect 13244 57708 13300 57764
rect 12796 56700 12852 56756
rect 12908 55410 12964 55412
rect 12908 55358 12910 55410
rect 12910 55358 12962 55410
rect 12962 55358 12964 55410
rect 12908 55356 12964 55358
rect 12124 55186 12180 55188
rect 12124 55134 12126 55186
rect 12126 55134 12178 55186
rect 12178 55134 12180 55186
rect 12124 55132 12180 55134
rect 11004 54572 11060 54628
rect 11116 54348 11172 54404
rect 10892 52220 10948 52276
rect 11228 52892 11284 52948
rect 10444 50764 10500 50820
rect 9996 49698 10052 49700
rect 9996 49646 9998 49698
rect 9998 49646 10050 49698
rect 10050 49646 10052 49698
rect 9996 49644 10052 49646
rect 9996 48354 10052 48356
rect 9996 48302 9998 48354
rect 9998 48302 10050 48354
rect 10050 48302 10052 48354
rect 9996 48300 10052 48302
rect 9884 47628 9940 47684
rect 10108 47740 10164 47796
rect 9996 47570 10052 47572
rect 9996 47518 9998 47570
rect 9998 47518 10050 47570
rect 10050 47518 10052 47570
rect 9996 47516 10052 47518
rect 9884 47404 9940 47460
rect 10332 49980 10388 50036
rect 11228 51772 11284 51828
rect 11452 51996 11508 52052
rect 11340 51660 11396 51716
rect 10332 49084 10388 49140
rect 10332 48354 10388 48356
rect 10332 48302 10334 48354
rect 10334 48302 10386 48354
rect 10386 48302 10388 48354
rect 10332 48300 10388 48302
rect 10332 47346 10388 47348
rect 10332 47294 10334 47346
rect 10334 47294 10386 47346
rect 10386 47294 10388 47346
rect 10332 47292 10388 47294
rect 9996 46284 10052 46340
rect 10108 45778 10164 45780
rect 10108 45726 10110 45778
rect 10110 45726 10162 45778
rect 10162 45726 10164 45778
rect 10108 45724 10164 45726
rect 10668 49698 10724 49700
rect 10668 49646 10670 49698
rect 10670 49646 10722 49698
rect 10722 49646 10724 49698
rect 10668 49644 10724 49646
rect 10780 49084 10836 49140
rect 10556 48914 10612 48916
rect 10556 48862 10558 48914
rect 10558 48862 10610 48914
rect 10610 48862 10612 48914
rect 10556 48860 10612 48862
rect 10780 48748 10836 48804
rect 10556 47516 10612 47572
rect 10332 46284 10388 46340
rect 9772 45218 9828 45220
rect 9772 45166 9774 45218
rect 9774 45166 9826 45218
rect 9826 45166 9828 45218
rect 9772 45164 9828 45166
rect 9660 44322 9716 44324
rect 9660 44270 9662 44322
rect 9662 44270 9714 44322
rect 9714 44270 9716 44322
rect 9660 44268 9716 44270
rect 9436 44210 9492 44212
rect 9436 44158 9438 44210
rect 9438 44158 9490 44210
rect 9490 44158 9492 44210
rect 9436 44156 9492 44158
rect 9772 44156 9828 44212
rect 9772 43820 9828 43876
rect 9548 43036 9604 43092
rect 9548 42140 9604 42196
rect 9324 42028 9380 42084
rect 9884 42700 9940 42756
rect 9772 41916 9828 41972
rect 9772 41132 9828 41188
rect 8876 40626 8932 40628
rect 8876 40574 8878 40626
rect 8878 40574 8930 40626
rect 8930 40574 8932 40626
rect 8876 40572 8932 40574
rect 9884 40572 9940 40628
rect 7980 39618 8036 39620
rect 7980 39566 7982 39618
rect 7982 39566 8034 39618
rect 8034 39566 8036 39618
rect 7980 39564 8036 39566
rect 8204 39340 8260 39396
rect 8428 39340 8484 39396
rect 7756 39228 7812 39284
rect 8092 39058 8148 39060
rect 8092 39006 8094 39058
rect 8094 39006 8146 39058
rect 8146 39006 8148 39058
rect 8092 39004 8148 39006
rect 7420 38556 7476 38612
rect 6972 37436 7028 37492
rect 7308 38220 7364 38276
rect 6748 37212 6804 37268
rect 7196 37378 7252 37380
rect 7196 37326 7198 37378
rect 7198 37326 7250 37378
rect 7250 37326 7252 37378
rect 7196 37324 7252 37326
rect 7420 38108 7476 38164
rect 7532 38050 7588 38052
rect 7532 37998 7534 38050
rect 7534 37998 7586 38050
rect 7586 37998 7588 38050
rect 7532 37996 7588 37998
rect 6860 36652 6916 36708
rect 6972 36764 7028 36820
rect 6748 36428 6804 36484
rect 7420 36876 7476 36932
rect 7532 36540 7588 36596
rect 7308 35084 7364 35140
rect 6860 34636 6916 34692
rect 6636 33906 6692 33908
rect 6636 33854 6638 33906
rect 6638 33854 6690 33906
rect 6690 33854 6692 33906
rect 6636 33852 6692 33854
rect 7308 33852 7364 33908
rect 6748 33234 6804 33236
rect 6748 33182 6750 33234
rect 6750 33182 6802 33234
rect 6802 33182 6804 33234
rect 6748 33180 6804 33182
rect 6412 32786 6468 32788
rect 6412 32734 6414 32786
rect 6414 32734 6466 32786
rect 6466 32734 6468 32786
rect 6412 32732 6468 32734
rect 7196 32786 7252 32788
rect 7196 32734 7198 32786
rect 7198 32734 7250 32786
rect 7250 32734 7252 32786
rect 7196 32732 7252 32734
rect 6412 32172 6468 32228
rect 6636 31388 6692 31444
rect 7420 33234 7476 33236
rect 7420 33182 7422 33234
rect 7422 33182 7474 33234
rect 7474 33182 7476 33234
rect 7420 33180 7476 33182
rect 7420 31612 7476 31668
rect 6748 30828 6804 30884
rect 7308 30210 7364 30212
rect 7308 30158 7310 30210
rect 7310 30158 7362 30210
rect 7362 30158 7364 30210
rect 7308 30156 7364 30158
rect 6412 30098 6468 30100
rect 6412 30046 6414 30098
rect 6414 30046 6466 30098
rect 6466 30046 6468 30098
rect 6412 30044 6468 30046
rect 6636 30044 6692 30100
rect 7644 35084 7700 35140
rect 7980 38444 8036 38500
rect 8204 38332 8260 38388
rect 8204 38108 8260 38164
rect 8092 36482 8148 36484
rect 8092 36430 8094 36482
rect 8094 36430 8146 36482
rect 8146 36430 8148 36482
rect 8092 36428 8148 36430
rect 8876 40348 8932 40404
rect 8652 38834 8708 38836
rect 8652 38782 8654 38834
rect 8654 38782 8706 38834
rect 8706 38782 8708 38834
rect 8652 38780 8708 38782
rect 9772 40402 9828 40404
rect 9772 40350 9774 40402
rect 9774 40350 9826 40402
rect 9826 40350 9828 40402
rect 9772 40348 9828 40350
rect 10220 45388 10276 45444
rect 10444 45724 10500 45780
rect 10220 42812 10276 42868
rect 10108 42364 10164 42420
rect 10668 46956 10724 47012
rect 11340 50876 11396 50932
rect 12796 54908 12852 54964
rect 12236 54684 12292 54740
rect 12460 54626 12516 54628
rect 12460 54574 12462 54626
rect 12462 54574 12514 54626
rect 12514 54574 12516 54626
rect 12460 54572 12516 54574
rect 11676 51548 11732 51604
rect 11564 51100 11620 51156
rect 11340 49308 11396 49364
rect 11340 49084 11396 49140
rect 11452 50204 11508 50260
rect 11676 50204 11732 50260
rect 11564 49644 11620 49700
rect 11676 48914 11732 48916
rect 11676 48862 11678 48914
rect 11678 48862 11730 48914
rect 11730 48862 11732 48914
rect 11676 48860 11732 48862
rect 11228 48300 11284 48356
rect 11116 48242 11172 48244
rect 11116 48190 11118 48242
rect 11118 48190 11170 48242
rect 11170 48190 11172 48242
rect 11116 48188 11172 48190
rect 10892 47516 10948 47572
rect 11004 48076 11060 48132
rect 10780 45724 10836 45780
rect 10892 46284 10948 46340
rect 10780 43372 10836 43428
rect 10444 42642 10500 42644
rect 10444 42590 10446 42642
rect 10446 42590 10498 42642
rect 10498 42590 10500 42642
rect 10444 42588 10500 42590
rect 10332 41970 10388 41972
rect 10332 41918 10334 41970
rect 10334 41918 10386 41970
rect 10386 41918 10388 41970
rect 10332 41916 10388 41918
rect 10668 41916 10724 41972
rect 11340 47180 11396 47236
rect 11228 46674 11284 46676
rect 11228 46622 11230 46674
rect 11230 46622 11282 46674
rect 11282 46622 11284 46674
rect 11228 46620 11284 46622
rect 11676 48636 11732 48692
rect 11676 48242 11732 48244
rect 11676 48190 11678 48242
rect 11678 48190 11730 48242
rect 11730 48190 11732 48242
rect 11676 48188 11732 48190
rect 11900 52332 11956 52388
rect 12572 53506 12628 53508
rect 12572 53454 12574 53506
rect 12574 53454 12626 53506
rect 12626 53454 12628 53506
rect 12572 53452 12628 53454
rect 12572 52946 12628 52948
rect 12572 52894 12574 52946
rect 12574 52894 12626 52946
rect 12626 52894 12628 52946
rect 12572 52892 12628 52894
rect 12124 52220 12180 52276
rect 13132 54908 13188 54964
rect 13132 54684 13188 54740
rect 13132 54348 13188 54404
rect 13020 54236 13076 54292
rect 13020 53004 13076 53060
rect 13132 52946 13188 52948
rect 13132 52894 13134 52946
rect 13134 52894 13186 52946
rect 13186 52894 13188 52946
rect 13132 52892 13188 52894
rect 12796 52332 12852 52388
rect 13020 52332 13076 52388
rect 12684 52220 12740 52276
rect 12908 52274 12964 52276
rect 12908 52222 12910 52274
rect 12910 52222 12962 52274
rect 12962 52222 12964 52274
rect 12908 52220 12964 52222
rect 12572 52050 12628 52052
rect 12572 51998 12574 52050
rect 12574 51998 12626 52050
rect 12626 51998 12628 52050
rect 12572 51996 12628 51998
rect 12124 51884 12180 51940
rect 12348 51938 12404 51940
rect 12348 51886 12350 51938
rect 12350 51886 12402 51938
rect 12402 51886 12404 51938
rect 12348 51884 12404 51886
rect 12236 51490 12292 51492
rect 12236 51438 12238 51490
rect 12238 51438 12290 51490
rect 12290 51438 12292 51490
rect 12236 51436 12292 51438
rect 12124 51378 12180 51380
rect 12124 51326 12126 51378
rect 12126 51326 12178 51378
rect 12178 51326 12180 51378
rect 12124 51324 12180 51326
rect 12460 51378 12516 51380
rect 12460 51326 12462 51378
rect 12462 51326 12514 51378
rect 12514 51326 12516 51378
rect 12460 51324 12516 51326
rect 12236 51212 12292 51268
rect 12124 50876 12180 50932
rect 12012 50652 12068 50708
rect 11900 49420 11956 49476
rect 13020 51100 13076 51156
rect 12348 50092 12404 50148
rect 12124 48130 12180 48132
rect 12124 48078 12126 48130
rect 12126 48078 12178 48130
rect 12178 48078 12180 48130
rect 12124 48076 12180 48078
rect 12012 47570 12068 47572
rect 12012 47518 12014 47570
rect 12014 47518 12066 47570
rect 12066 47518 12068 47570
rect 12012 47516 12068 47518
rect 13020 50652 13076 50708
rect 12908 49810 12964 49812
rect 12908 49758 12910 49810
rect 12910 49758 12962 49810
rect 12962 49758 12964 49810
rect 12908 49756 12964 49758
rect 12460 48748 12516 48804
rect 12796 48412 12852 48468
rect 12236 47292 12292 47348
rect 12460 48188 12516 48244
rect 12460 46732 12516 46788
rect 13692 57820 13748 57876
rect 13468 57260 13524 57316
rect 16380 57820 16436 57876
rect 13692 57260 13748 57316
rect 13916 57372 13972 57428
rect 13468 56476 13524 56532
rect 13804 54348 13860 54404
rect 14924 57372 14980 57428
rect 14812 57148 14868 57204
rect 15036 57148 15092 57204
rect 14140 56194 14196 56196
rect 14140 56142 14142 56194
rect 14142 56142 14194 56194
rect 14194 56142 14196 56194
rect 14140 56140 14196 56142
rect 13692 54124 13748 54180
rect 13804 53618 13860 53620
rect 13804 53566 13806 53618
rect 13806 53566 13858 53618
rect 13858 53566 13860 53618
rect 13804 53564 13860 53566
rect 13356 53116 13412 53172
rect 14028 56028 14084 56084
rect 13244 52556 13300 52612
rect 13244 52332 13300 52388
rect 14140 55804 14196 55860
rect 14140 55074 14196 55076
rect 14140 55022 14142 55074
rect 14142 55022 14194 55074
rect 14194 55022 14196 55074
rect 14140 55020 14196 55022
rect 14140 54460 14196 54516
rect 14140 53506 14196 53508
rect 14140 53454 14142 53506
rect 14142 53454 14194 53506
rect 14194 53454 14196 53506
rect 14140 53452 14196 53454
rect 13356 51100 13412 51156
rect 13692 51772 13748 51828
rect 13468 50988 13524 51044
rect 13244 50876 13300 50932
rect 13356 49756 13412 49812
rect 12908 48354 12964 48356
rect 12908 48302 12910 48354
rect 12910 48302 12962 48354
rect 12962 48302 12964 48354
rect 12908 48300 12964 48302
rect 13244 48354 13300 48356
rect 13244 48302 13246 48354
rect 13246 48302 13298 48354
rect 13298 48302 13300 48354
rect 13244 48300 13300 48302
rect 13020 47740 13076 47796
rect 13356 47740 13412 47796
rect 13132 47628 13188 47684
rect 12796 47234 12852 47236
rect 12796 47182 12798 47234
rect 12798 47182 12850 47234
rect 12850 47182 12852 47234
rect 12796 47180 12852 47182
rect 12572 47068 12628 47124
rect 11564 46562 11620 46564
rect 11564 46510 11566 46562
rect 11566 46510 11618 46562
rect 11618 46510 11620 46562
rect 11564 46508 11620 46510
rect 11340 46060 11396 46116
rect 11228 45778 11284 45780
rect 11228 45726 11230 45778
rect 11230 45726 11282 45778
rect 11282 45726 11284 45778
rect 11228 45724 11284 45726
rect 11340 44716 11396 44772
rect 12124 46674 12180 46676
rect 12124 46622 12126 46674
rect 12126 46622 12178 46674
rect 12178 46622 12180 46674
rect 12124 46620 12180 46622
rect 12460 45724 12516 45780
rect 11452 44268 11508 44324
rect 10892 43036 10948 43092
rect 11004 43484 11060 43540
rect 10780 42364 10836 42420
rect 9100 40124 9156 40180
rect 9548 39618 9604 39620
rect 9548 39566 9550 39618
rect 9550 39566 9602 39618
rect 9602 39566 9604 39618
rect 9548 39564 9604 39566
rect 9100 39506 9156 39508
rect 9100 39454 9102 39506
rect 9102 39454 9154 39506
rect 9154 39454 9156 39506
rect 9100 39452 9156 39454
rect 8876 39228 8932 39284
rect 8540 37996 8596 38052
rect 8316 36428 8372 36484
rect 7980 35532 8036 35588
rect 7644 34242 7700 34244
rect 7644 34190 7646 34242
rect 7646 34190 7698 34242
rect 7698 34190 7700 34242
rect 7644 34188 7700 34190
rect 7756 33852 7812 33908
rect 7644 32956 7700 33012
rect 8428 35756 8484 35812
rect 8092 35084 8148 35140
rect 8204 34802 8260 34804
rect 8204 34750 8206 34802
rect 8206 34750 8258 34802
rect 8258 34750 8260 34802
rect 8204 34748 8260 34750
rect 8652 35698 8708 35700
rect 8652 35646 8654 35698
rect 8654 35646 8706 35698
rect 8706 35646 8708 35698
rect 8652 35644 8708 35646
rect 9100 38444 9156 38500
rect 9212 37884 9268 37940
rect 8988 37378 9044 37380
rect 8988 37326 8990 37378
rect 8990 37326 9042 37378
rect 9042 37326 9044 37378
rect 8988 37324 9044 37326
rect 9212 36594 9268 36596
rect 9212 36542 9214 36594
rect 9214 36542 9266 36594
rect 9266 36542 9268 36594
rect 9212 36540 9268 36542
rect 8876 35810 8932 35812
rect 8876 35758 8878 35810
rect 8878 35758 8930 35810
rect 8930 35758 8932 35810
rect 8876 35756 8932 35758
rect 9548 35756 9604 35812
rect 8764 35532 8820 35588
rect 9100 35644 9156 35700
rect 8876 35420 8932 35476
rect 8988 35084 9044 35140
rect 8876 33852 8932 33908
rect 7868 31388 7924 31444
rect 7980 32620 8036 32676
rect 7644 30828 7700 30884
rect 9324 35084 9380 35140
rect 9100 34748 9156 34804
rect 9436 33516 9492 33572
rect 8540 32450 8596 32452
rect 8540 32398 8542 32450
rect 8542 32398 8594 32450
rect 8594 32398 8596 32450
rect 8540 32396 8596 32398
rect 8652 32172 8708 32228
rect 8988 32562 9044 32564
rect 8988 32510 8990 32562
rect 8990 32510 9042 32562
rect 9042 32510 9044 32562
rect 8988 32508 9044 32510
rect 8764 31836 8820 31892
rect 8764 31500 8820 31556
rect 8540 31388 8596 31444
rect 8092 31276 8148 31332
rect 8316 30156 8372 30212
rect 7980 30044 8036 30100
rect 7532 29820 7588 29876
rect 8204 29820 8260 29876
rect 6076 29484 6132 29540
rect 5516 28028 5572 28084
rect 5068 24332 5124 24388
rect 4956 23436 5012 23492
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 7196 29650 7252 29652
rect 7196 29598 7198 29650
rect 7198 29598 7250 29650
rect 7250 29598 7252 29650
rect 7196 29596 7252 29598
rect 7644 29650 7700 29652
rect 7644 29598 7646 29650
rect 7646 29598 7698 29650
rect 7698 29598 7700 29650
rect 7644 29596 7700 29598
rect 8652 30044 8708 30100
rect 9100 30994 9156 30996
rect 9100 30942 9102 30994
rect 9102 30942 9154 30994
rect 9154 30942 9156 30994
rect 9100 30940 9156 30942
rect 9212 30604 9268 30660
rect 9100 30098 9156 30100
rect 9100 30046 9102 30098
rect 9102 30046 9154 30098
rect 9154 30046 9156 30098
rect 9100 30044 9156 30046
rect 9100 29484 9156 29540
rect 6636 20860 6692 20916
rect 7532 26460 7588 26516
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 7532 17052 7588 17108
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 6972 14252 7028 14308
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 3724 12348 3780 12404
rect 2492 12012 2548 12068
rect 3164 12066 3220 12068
rect 3164 12014 3166 12066
rect 3166 12014 3218 12066
rect 3218 12014 3220 12066
rect 3164 12012 3220 12014
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 2716 10780 2772 10836
rect 3276 10834 3332 10836
rect 3276 10782 3278 10834
rect 3278 10782 3330 10834
rect 3330 10782 3332 10834
rect 3276 10780 3332 10782
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 2716 9714 2772 9716
rect 2716 9662 2718 9714
rect 2718 9662 2770 9714
rect 2770 9662 2772 9714
rect 2716 9660 2772 9662
rect 3276 9714 3332 9716
rect 3276 9662 3278 9714
rect 3278 9662 3330 9714
rect 3330 9662 3332 9714
rect 3276 9660 3332 9662
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 1932 5404 1988 5460
rect 2716 4508 2772 4564
rect 28 1820 84 1876
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 3276 4562 3332 4564
rect 3276 4510 3278 4562
rect 3278 4510 3330 4562
rect 3330 4510 3332 4562
rect 3276 4508 3332 4510
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 9996 39788 10052 39844
rect 10220 39452 10276 39508
rect 10668 41692 10724 41748
rect 11228 42700 11284 42756
rect 11340 42588 11396 42644
rect 11900 44994 11956 44996
rect 11900 44942 11902 44994
rect 11902 44942 11954 44994
rect 11954 44942 11956 44994
rect 11900 44940 11956 44942
rect 11676 44156 11732 44212
rect 11788 44828 11844 44884
rect 13692 51378 13748 51380
rect 13692 51326 13694 51378
rect 13694 51326 13746 51378
rect 13746 51326 13748 51378
rect 13692 51324 13748 51326
rect 13916 51660 13972 51716
rect 14028 51772 14084 51828
rect 13580 50876 13636 50932
rect 13804 50764 13860 50820
rect 14364 53116 14420 53172
rect 14476 53452 14532 53508
rect 14364 52834 14420 52836
rect 14364 52782 14366 52834
rect 14366 52782 14418 52834
rect 14418 52782 14420 52834
rect 14364 52780 14420 52782
rect 14700 54684 14756 54740
rect 14812 55020 14868 55076
rect 14924 56588 14980 56644
rect 14924 55132 14980 55188
rect 14812 54348 14868 54404
rect 14700 53730 14756 53732
rect 14700 53678 14702 53730
rect 14702 53678 14754 53730
rect 14754 53678 14756 53730
rect 14700 53676 14756 53678
rect 14588 53340 14644 53396
rect 14588 53004 14644 53060
rect 14364 51266 14420 51268
rect 14364 51214 14366 51266
rect 14366 51214 14418 51266
rect 14418 51214 14420 51266
rect 14364 51212 14420 51214
rect 14364 50764 14420 50820
rect 14252 50482 14308 50484
rect 14252 50430 14254 50482
rect 14254 50430 14306 50482
rect 14306 50430 14308 50482
rect 14252 50428 14308 50430
rect 14140 49868 14196 49924
rect 14028 49698 14084 49700
rect 14028 49646 14030 49698
rect 14030 49646 14082 49698
rect 14082 49646 14084 49698
rect 14028 49644 14084 49646
rect 14140 49308 14196 49364
rect 14252 49250 14308 49252
rect 14252 49198 14254 49250
rect 14254 49198 14306 49250
rect 14306 49198 14308 49250
rect 14252 49196 14308 49198
rect 14700 52946 14756 52948
rect 14700 52894 14702 52946
rect 14702 52894 14754 52946
rect 14754 52894 14756 52946
rect 14700 52892 14756 52894
rect 14812 52556 14868 52612
rect 14588 50428 14644 50484
rect 14700 52108 14756 52164
rect 14364 49084 14420 49140
rect 14140 49026 14196 49028
rect 14140 48974 14142 49026
rect 14142 48974 14194 49026
rect 14194 48974 14196 49026
rect 14140 48972 14196 48974
rect 13804 48412 13860 48468
rect 14364 48860 14420 48916
rect 14140 47964 14196 48020
rect 14028 47682 14084 47684
rect 14028 47630 14030 47682
rect 14030 47630 14082 47682
rect 14082 47630 14084 47682
rect 14028 47628 14084 47630
rect 14476 47628 14532 47684
rect 14476 47458 14532 47460
rect 14476 47406 14478 47458
rect 14478 47406 14530 47458
rect 14530 47406 14532 47458
rect 14476 47404 14532 47406
rect 13468 46844 13524 46900
rect 13468 46674 13524 46676
rect 13468 46622 13470 46674
rect 13470 46622 13522 46674
rect 13522 46622 13524 46674
rect 13468 46620 13524 46622
rect 13468 46060 13524 46116
rect 12684 45948 12740 46004
rect 12796 45500 12852 45556
rect 13020 45276 13076 45332
rect 14028 46844 14084 46900
rect 14028 46620 14084 46676
rect 14140 46732 14196 46788
rect 12236 44828 12292 44884
rect 14028 45948 14084 46004
rect 13804 45724 13860 45780
rect 13468 45164 13524 45220
rect 12012 44492 12068 44548
rect 11788 43932 11844 43988
rect 12572 44492 12628 44548
rect 12460 43932 12516 43988
rect 12348 43820 12404 43876
rect 12796 44828 12852 44884
rect 13468 44492 13524 44548
rect 12236 43596 12292 43652
rect 11564 42364 11620 42420
rect 11900 42924 11956 42980
rect 10108 39228 10164 39284
rect 9996 39116 10052 39172
rect 9884 38892 9940 38948
rect 10108 38946 10164 38948
rect 10108 38894 10110 38946
rect 10110 38894 10162 38946
rect 10162 38894 10164 38946
rect 10108 38892 10164 38894
rect 9884 38722 9940 38724
rect 9884 38670 9886 38722
rect 9886 38670 9938 38722
rect 9938 38670 9940 38722
rect 9884 38668 9940 38670
rect 9996 38556 10052 38612
rect 10108 37772 10164 37828
rect 9884 37660 9940 37716
rect 9884 37490 9940 37492
rect 9884 37438 9886 37490
rect 9886 37438 9938 37490
rect 9938 37438 9940 37490
rect 9884 37436 9940 37438
rect 9772 35756 9828 35812
rect 9660 35420 9716 35476
rect 9996 35868 10052 35924
rect 9884 35084 9940 35140
rect 10220 36428 10276 36484
rect 9884 34354 9940 34356
rect 9884 34302 9886 34354
rect 9886 34302 9938 34354
rect 9938 34302 9940 34354
rect 9884 34300 9940 34302
rect 10668 41020 10724 41076
rect 11116 40572 11172 40628
rect 10780 40236 10836 40292
rect 11452 41858 11508 41860
rect 11452 41806 11454 41858
rect 11454 41806 11506 41858
rect 11506 41806 11508 41858
rect 11452 41804 11508 41806
rect 11452 41468 11508 41524
rect 11564 40908 11620 40964
rect 11564 40460 11620 40516
rect 11564 40012 11620 40068
rect 10444 39452 10500 39508
rect 10444 39116 10500 39172
rect 10556 39228 10612 39284
rect 10780 39452 10836 39508
rect 11228 39228 11284 39284
rect 10444 37324 10500 37380
rect 10556 37100 10612 37156
rect 10668 36876 10724 36932
rect 10556 36482 10612 36484
rect 10556 36430 10558 36482
rect 10558 36430 10610 36482
rect 10610 36430 10612 36482
rect 10556 36428 10612 36430
rect 10668 36370 10724 36372
rect 10668 36318 10670 36370
rect 10670 36318 10722 36370
rect 10722 36318 10724 36370
rect 10668 36316 10724 36318
rect 10220 35196 10276 35252
rect 10332 35308 10388 35364
rect 9548 32732 9604 32788
rect 9996 32562 10052 32564
rect 9996 32510 9998 32562
rect 9998 32510 10050 32562
rect 10050 32510 10052 32562
rect 9996 32508 10052 32510
rect 9884 32172 9940 32228
rect 9996 31836 10052 31892
rect 9884 31612 9940 31668
rect 9772 31554 9828 31556
rect 9772 31502 9774 31554
rect 9774 31502 9826 31554
rect 9826 31502 9828 31554
rect 9772 31500 9828 31502
rect 9548 31388 9604 31444
rect 10332 32338 10388 32340
rect 10332 32286 10334 32338
rect 10334 32286 10386 32338
rect 10386 32286 10388 32338
rect 10332 32284 10388 32286
rect 10220 31836 10276 31892
rect 10108 31778 10164 31780
rect 10108 31726 10110 31778
rect 10110 31726 10162 31778
rect 10162 31726 10164 31778
rect 10108 31724 10164 31726
rect 9436 30044 9492 30100
rect 9996 30716 10052 30772
rect 9660 29986 9716 29988
rect 9660 29934 9662 29986
rect 9662 29934 9714 29986
rect 9714 29934 9716 29986
rect 9660 29932 9716 29934
rect 9660 29538 9716 29540
rect 9660 29486 9662 29538
rect 9662 29486 9714 29538
rect 9714 29486 9716 29538
rect 9660 29484 9716 29486
rect 9660 28252 9716 28308
rect 10332 30994 10388 30996
rect 10332 30942 10334 30994
rect 10334 30942 10386 30994
rect 10386 30942 10388 30994
rect 10332 30940 10388 30942
rect 10556 34802 10612 34804
rect 10556 34750 10558 34802
rect 10558 34750 10610 34802
rect 10610 34750 10612 34802
rect 10556 34748 10612 34750
rect 11116 38946 11172 38948
rect 11116 38894 11118 38946
rect 11118 38894 11170 38946
rect 11170 38894 11172 38946
rect 11116 38892 11172 38894
rect 11788 41916 11844 41972
rect 11676 39788 11732 39844
rect 11004 35810 11060 35812
rect 11004 35758 11006 35810
rect 11006 35758 11058 35810
rect 11058 35758 11060 35810
rect 11004 35756 11060 35758
rect 10780 34860 10836 34916
rect 11788 38050 11844 38052
rect 11788 37998 11790 38050
rect 11790 37998 11842 38050
rect 11842 37998 11844 38050
rect 11788 37996 11844 37998
rect 11676 37884 11732 37940
rect 11228 37660 11284 37716
rect 11564 37660 11620 37716
rect 11452 35698 11508 35700
rect 11452 35646 11454 35698
rect 11454 35646 11506 35698
rect 11506 35646 11508 35698
rect 11452 35644 11508 35646
rect 11340 35586 11396 35588
rect 11340 35534 11342 35586
rect 11342 35534 11394 35586
rect 11394 35534 11396 35586
rect 11340 35532 11396 35534
rect 12124 42754 12180 42756
rect 12124 42702 12126 42754
rect 12126 42702 12178 42754
rect 12178 42702 12180 42754
rect 12124 42700 12180 42702
rect 12124 42364 12180 42420
rect 12684 42028 12740 42084
rect 13692 44210 13748 44212
rect 13692 44158 13694 44210
rect 13694 44158 13746 44210
rect 13746 44158 13748 44210
rect 13692 44156 13748 44158
rect 13468 44044 13524 44100
rect 13356 43538 13412 43540
rect 13356 43486 13358 43538
rect 13358 43486 13410 43538
rect 13410 43486 13412 43538
rect 13356 43484 13412 43486
rect 13692 43708 13748 43764
rect 13580 43650 13636 43652
rect 13580 43598 13582 43650
rect 13582 43598 13634 43650
rect 13634 43598 13636 43650
rect 13580 43596 13636 43598
rect 13132 42476 13188 42532
rect 13132 42252 13188 42308
rect 13020 41916 13076 41972
rect 12012 41132 12068 41188
rect 12012 40908 12068 40964
rect 12124 41356 12180 41412
rect 12012 38722 12068 38724
rect 12012 38670 12014 38722
rect 12014 38670 12066 38722
rect 12066 38670 12068 38722
rect 12012 38668 12068 38670
rect 11900 36540 11956 36596
rect 11676 35980 11732 36036
rect 12012 35980 12068 36036
rect 11900 35810 11956 35812
rect 11900 35758 11902 35810
rect 11902 35758 11954 35810
rect 11954 35758 11956 35810
rect 11900 35756 11956 35758
rect 11116 34914 11172 34916
rect 11116 34862 11118 34914
rect 11118 34862 11170 34914
rect 11170 34862 11172 34914
rect 11116 34860 11172 34862
rect 11116 33404 11172 33460
rect 10668 31836 10724 31892
rect 11340 34860 11396 34916
rect 11452 34748 11508 34804
rect 11676 34860 11732 34916
rect 11676 34412 11732 34468
rect 12236 40796 12292 40852
rect 12908 40514 12964 40516
rect 12908 40462 12910 40514
rect 12910 40462 12962 40514
rect 12962 40462 12964 40514
rect 12908 40460 12964 40462
rect 12460 40012 12516 40068
rect 12348 39340 12404 39396
rect 12236 37996 12292 38052
rect 12348 37826 12404 37828
rect 12348 37774 12350 37826
rect 12350 37774 12402 37826
rect 12402 37774 12404 37826
rect 12348 37772 12404 37774
rect 12124 35644 12180 35700
rect 12236 36540 12292 36596
rect 11564 34076 11620 34132
rect 11676 33628 11732 33684
rect 10556 31666 10612 31668
rect 10556 31614 10558 31666
rect 10558 31614 10610 31666
rect 10610 31614 10612 31666
rect 10556 31612 10612 31614
rect 10780 31500 10836 31556
rect 10556 30940 10612 30996
rect 10892 30156 10948 30212
rect 11116 32002 11172 32004
rect 11116 31950 11118 32002
rect 11118 31950 11170 32002
rect 11170 31950 11172 32002
rect 11116 31948 11172 31950
rect 11676 32786 11732 32788
rect 11676 32734 11678 32786
rect 11678 32734 11730 32786
rect 11730 32734 11732 32786
rect 11676 32732 11732 32734
rect 11676 31836 11732 31892
rect 12572 39116 12628 39172
rect 12684 38834 12740 38836
rect 12684 38782 12686 38834
rect 12686 38782 12738 38834
rect 12738 38782 12740 38834
rect 12684 38780 12740 38782
rect 12684 38332 12740 38388
rect 12908 39730 12964 39732
rect 12908 39678 12910 39730
rect 12910 39678 12962 39730
rect 12962 39678 12964 39730
rect 12908 39676 12964 39678
rect 12796 38108 12852 38164
rect 12572 37436 12628 37492
rect 12460 36092 12516 36148
rect 13244 41746 13300 41748
rect 13244 41694 13246 41746
rect 13246 41694 13298 41746
rect 13298 41694 13300 41746
rect 13244 41692 13300 41694
rect 13132 41244 13188 41300
rect 13692 42642 13748 42644
rect 13692 42590 13694 42642
rect 13694 42590 13746 42642
rect 13746 42590 13748 42642
rect 13692 42588 13748 42590
rect 14476 46396 14532 46452
rect 14252 45330 14308 45332
rect 14252 45278 14254 45330
rect 14254 45278 14306 45330
rect 14306 45278 14308 45330
rect 14252 45276 14308 45278
rect 14364 45106 14420 45108
rect 14364 45054 14366 45106
rect 14366 45054 14418 45106
rect 14418 45054 14420 45106
rect 14364 45052 14420 45054
rect 14588 45500 14644 45556
rect 15148 55298 15204 55300
rect 15148 55246 15150 55298
rect 15150 55246 15202 55298
rect 15202 55246 15204 55298
rect 15148 55244 15204 55246
rect 15148 54684 15204 54740
rect 15260 53452 15316 53508
rect 15372 54236 15428 54292
rect 15148 53228 15204 53284
rect 15036 53116 15092 53172
rect 15148 52780 15204 52836
rect 15036 52332 15092 52388
rect 14924 51772 14980 51828
rect 14924 51100 14980 51156
rect 15372 51884 15428 51940
rect 15148 50316 15204 50372
rect 15036 49980 15092 50036
rect 15708 55916 15764 55972
rect 15596 55132 15652 55188
rect 15596 53730 15652 53732
rect 15596 53678 15598 53730
rect 15598 53678 15650 53730
rect 15650 53678 15652 53730
rect 15596 53676 15652 53678
rect 15596 52332 15652 52388
rect 15932 54514 15988 54516
rect 15932 54462 15934 54514
rect 15934 54462 15986 54514
rect 15986 54462 15988 54514
rect 15932 54460 15988 54462
rect 15820 53676 15876 53732
rect 17388 56476 17444 56532
rect 16828 55468 16884 55524
rect 16940 55804 16996 55860
rect 16156 55244 16212 55300
rect 16156 53900 16212 53956
rect 16604 55186 16660 55188
rect 16604 55134 16606 55186
rect 16606 55134 16658 55186
rect 16658 55134 16660 55186
rect 16604 55132 16660 55134
rect 16380 55020 16436 55076
rect 16492 54514 16548 54516
rect 16492 54462 16494 54514
rect 16494 54462 16546 54514
rect 16546 54462 16548 54514
rect 16492 54460 16548 54462
rect 16380 53900 16436 53956
rect 17276 55186 17332 55188
rect 17276 55134 17278 55186
rect 17278 55134 17330 55186
rect 17330 55134 17332 55186
rect 17276 55132 17332 55134
rect 17164 54908 17220 54964
rect 17164 54348 17220 54404
rect 17500 56082 17556 56084
rect 17500 56030 17502 56082
rect 17502 56030 17554 56082
rect 17554 56030 17556 56082
rect 17500 56028 17556 56030
rect 21868 58044 21924 58100
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 21868 56364 21924 56420
rect 18508 56082 18564 56084
rect 18508 56030 18510 56082
rect 18510 56030 18562 56082
rect 18562 56030 18564 56082
rect 18508 56028 18564 56030
rect 21644 56028 21700 56084
rect 18172 55916 18228 55972
rect 19068 55970 19124 55972
rect 19068 55918 19070 55970
rect 19070 55918 19122 55970
rect 19122 55918 19124 55970
rect 19068 55916 19124 55918
rect 17948 55804 18004 55860
rect 17836 55580 17892 55636
rect 19852 55580 19908 55636
rect 19516 55468 19572 55524
rect 19180 55132 19236 55188
rect 18172 54796 18228 54852
rect 17388 54236 17444 54292
rect 17948 54290 18004 54292
rect 17948 54238 17950 54290
rect 17950 54238 18002 54290
rect 18002 54238 18004 54290
rect 17948 54236 18004 54238
rect 18172 54236 18228 54292
rect 16268 53452 16324 53508
rect 16380 53340 16436 53396
rect 16156 52834 16212 52836
rect 16156 52782 16158 52834
rect 16158 52782 16210 52834
rect 16210 52782 16212 52834
rect 16156 52780 16212 52782
rect 16492 52834 16548 52836
rect 16492 52782 16494 52834
rect 16494 52782 16546 52834
rect 16546 52782 16548 52834
rect 16492 52780 16548 52782
rect 16828 53116 16884 53172
rect 17836 53788 17892 53844
rect 17052 53452 17108 53508
rect 16716 53004 16772 53060
rect 16380 52108 16436 52164
rect 16604 52556 16660 52612
rect 15708 51772 15764 51828
rect 16268 52050 16324 52052
rect 16268 51998 16270 52050
rect 16270 51998 16322 52050
rect 16322 51998 16324 52050
rect 16268 51996 16324 51998
rect 16492 52050 16548 52052
rect 16492 51998 16494 52050
rect 16494 51998 16546 52050
rect 16546 51998 16548 52050
rect 16492 51996 16548 51998
rect 16380 51660 16436 51716
rect 16492 51772 16548 51828
rect 16380 51324 16436 51380
rect 16492 50988 16548 51044
rect 16268 50876 16324 50932
rect 15372 49980 15428 50036
rect 15484 50204 15540 50260
rect 15484 49810 15540 49812
rect 15484 49758 15486 49810
rect 15486 49758 15538 49810
rect 15538 49758 15540 49810
rect 15484 49756 15540 49758
rect 15708 49532 15764 49588
rect 14924 48860 14980 48916
rect 15148 48524 15204 48580
rect 14476 44604 14532 44660
rect 14140 44380 14196 44436
rect 14140 44098 14196 44100
rect 14140 44046 14142 44098
rect 14142 44046 14194 44098
rect 14194 44046 14196 44098
rect 14140 44044 14196 44046
rect 14252 44268 14308 44324
rect 14028 43538 14084 43540
rect 14028 43486 14030 43538
rect 14030 43486 14082 43538
rect 14082 43486 14084 43538
rect 14028 43484 14084 43486
rect 14140 43426 14196 43428
rect 14140 43374 14142 43426
rect 14142 43374 14194 43426
rect 14194 43374 14196 43426
rect 14140 43372 14196 43374
rect 14364 43260 14420 43316
rect 14028 42812 14084 42868
rect 13916 42642 13972 42644
rect 13916 42590 13918 42642
rect 13918 42590 13970 42642
rect 13970 42590 13972 42642
rect 13916 42588 13972 42590
rect 13692 42364 13748 42420
rect 13580 41916 13636 41972
rect 13580 41132 13636 41188
rect 14140 42140 14196 42196
rect 14364 42700 14420 42756
rect 14588 43260 14644 43316
rect 14588 42252 14644 42308
rect 13916 41746 13972 41748
rect 13916 41694 13918 41746
rect 13918 41694 13970 41746
rect 13970 41694 13972 41746
rect 13916 41692 13972 41694
rect 14028 41410 14084 41412
rect 14028 41358 14030 41410
rect 14030 41358 14082 41410
rect 14082 41358 14084 41410
rect 14028 41356 14084 41358
rect 13580 40460 13636 40516
rect 14028 40908 14084 40964
rect 14252 41746 14308 41748
rect 14252 41694 14254 41746
rect 14254 41694 14306 41746
rect 14306 41694 14308 41746
rect 14252 41692 14308 41694
rect 14364 41356 14420 41412
rect 14252 41186 14308 41188
rect 14252 41134 14254 41186
rect 14254 41134 14306 41186
rect 14306 41134 14308 41186
rect 14252 41132 14308 41134
rect 13916 40348 13972 40404
rect 13356 40236 13412 40292
rect 13020 37436 13076 37492
rect 13356 40012 13412 40068
rect 13692 40012 13748 40068
rect 13916 40012 13972 40068
rect 13468 39564 13524 39620
rect 13580 39676 13636 39732
rect 12908 36482 12964 36484
rect 12908 36430 12910 36482
rect 12910 36430 12962 36482
rect 12962 36430 12964 36482
rect 12908 36428 12964 36430
rect 13020 36092 13076 36148
rect 12908 35980 12964 36036
rect 12460 35420 12516 35476
rect 12572 35026 12628 35028
rect 12572 34974 12574 35026
rect 12574 34974 12626 35026
rect 12626 34974 12628 35026
rect 12572 34972 12628 34974
rect 12908 35196 12964 35252
rect 12796 34748 12852 34804
rect 12572 34636 12628 34692
rect 12572 34354 12628 34356
rect 12572 34302 12574 34354
rect 12574 34302 12626 34354
rect 12626 34302 12628 34354
rect 12572 34300 12628 34302
rect 13244 35980 13300 36036
rect 13020 34018 13076 34020
rect 13020 33966 13022 34018
rect 13022 33966 13074 34018
rect 13074 33966 13076 34018
rect 13020 33964 13076 33966
rect 13132 35756 13188 35812
rect 12908 33346 12964 33348
rect 12908 33294 12910 33346
rect 12910 33294 12962 33346
rect 12962 33294 12964 33346
rect 12908 33292 12964 33294
rect 11900 32396 11956 32452
rect 11900 31948 11956 32004
rect 12236 33122 12292 33124
rect 12236 33070 12238 33122
rect 12238 33070 12290 33122
rect 12290 33070 12292 33122
rect 12236 33068 12292 33070
rect 12796 33068 12852 33124
rect 13468 38892 13524 38948
rect 13692 39340 13748 39396
rect 13580 38108 13636 38164
rect 14252 39618 14308 39620
rect 14252 39566 14254 39618
rect 14254 39566 14306 39618
rect 14306 39566 14308 39618
rect 14252 39564 14308 39566
rect 14252 38946 14308 38948
rect 14252 38894 14254 38946
rect 14254 38894 14306 38946
rect 14306 38894 14308 38946
rect 14252 38892 14308 38894
rect 14140 38668 14196 38724
rect 14476 39900 14532 39956
rect 14588 38946 14644 38948
rect 14588 38894 14590 38946
rect 14590 38894 14642 38946
rect 14642 38894 14644 38946
rect 14588 38892 14644 38894
rect 15036 47628 15092 47684
rect 14812 47180 14868 47236
rect 14924 46562 14980 46564
rect 14924 46510 14926 46562
rect 14926 46510 14978 46562
rect 14978 46510 14980 46562
rect 14924 46508 14980 46510
rect 15260 48466 15316 48468
rect 15260 48414 15262 48466
rect 15262 48414 15314 48466
rect 15314 48414 15316 48466
rect 15260 48412 15316 48414
rect 15260 47740 15316 47796
rect 15148 47234 15204 47236
rect 15148 47182 15150 47234
rect 15150 47182 15202 47234
rect 15202 47182 15204 47234
rect 15148 47180 15204 47182
rect 15260 47068 15316 47124
rect 15036 45724 15092 45780
rect 15148 45218 15204 45220
rect 15148 45166 15150 45218
rect 15150 45166 15202 45218
rect 15202 45166 15204 45218
rect 15148 45164 15204 45166
rect 15372 46562 15428 46564
rect 15372 46510 15374 46562
rect 15374 46510 15426 46562
rect 15426 46510 15428 46562
rect 15372 46508 15428 46510
rect 15484 46284 15540 46340
rect 15820 49980 15876 50036
rect 16156 50594 16212 50596
rect 16156 50542 16158 50594
rect 16158 50542 16210 50594
rect 16210 50542 16212 50594
rect 16156 50540 16212 50542
rect 16156 50316 16212 50372
rect 15932 49922 15988 49924
rect 15932 49870 15934 49922
rect 15934 49870 15986 49922
rect 15986 49870 15988 49922
rect 15932 49868 15988 49870
rect 16156 49026 16212 49028
rect 16156 48974 16158 49026
rect 16158 48974 16210 49026
rect 16210 48974 16212 49026
rect 16156 48972 16212 48974
rect 16492 49980 16548 50036
rect 16380 49810 16436 49812
rect 16380 49758 16382 49810
rect 16382 49758 16434 49810
rect 16434 49758 16436 49810
rect 16380 49756 16436 49758
rect 16268 49308 16324 49364
rect 15820 48860 15876 48916
rect 16044 48748 16100 48804
rect 15708 47068 15764 47124
rect 15596 46620 15652 46676
rect 15596 46060 15652 46116
rect 15708 46732 15764 46788
rect 15372 45836 15428 45892
rect 15932 46732 15988 46788
rect 15820 46562 15876 46564
rect 15820 46510 15822 46562
rect 15822 46510 15874 46562
rect 15874 46510 15876 46562
rect 15820 46508 15876 46510
rect 16940 52332 16996 52388
rect 16828 51996 16884 52052
rect 16716 51938 16772 51940
rect 16716 51886 16718 51938
rect 16718 51886 16770 51938
rect 16770 51886 16772 51938
rect 16716 51884 16772 51886
rect 16940 51378 16996 51380
rect 16940 51326 16942 51378
rect 16942 51326 16994 51378
rect 16994 51326 16996 51378
rect 16940 51324 16996 51326
rect 17164 52556 17220 52612
rect 17164 51996 17220 52052
rect 17500 53228 17556 53284
rect 17500 52668 17556 52724
rect 17724 52444 17780 52500
rect 16828 50316 16884 50372
rect 17388 50482 17444 50484
rect 17388 50430 17390 50482
rect 17390 50430 17442 50482
rect 17442 50430 17444 50482
rect 17388 50428 17444 50430
rect 16716 50034 16772 50036
rect 16716 49982 16718 50034
rect 16718 49982 16770 50034
rect 16770 49982 16772 50034
rect 16716 49980 16772 49982
rect 16940 49756 16996 49812
rect 17388 49868 17444 49924
rect 16604 48354 16660 48356
rect 16604 48302 16606 48354
rect 16606 48302 16658 48354
rect 16658 48302 16660 48354
rect 16604 48300 16660 48302
rect 16044 46172 16100 46228
rect 16156 45890 16212 45892
rect 16156 45838 16158 45890
rect 16158 45838 16210 45890
rect 16210 45838 16212 45890
rect 16156 45836 16212 45838
rect 15820 45724 15876 45780
rect 15372 45500 15428 45556
rect 15260 44546 15316 44548
rect 15260 44494 15262 44546
rect 15262 44494 15314 44546
rect 15314 44494 15316 44546
rect 15260 44492 15316 44494
rect 15148 44044 15204 44100
rect 15708 45388 15764 45444
rect 15596 45276 15652 45332
rect 15596 44994 15652 44996
rect 15596 44942 15598 44994
rect 15598 44942 15650 44994
rect 15650 44942 15652 44994
rect 15596 44940 15652 44942
rect 15148 43650 15204 43652
rect 15148 43598 15150 43650
rect 15150 43598 15202 43650
rect 15202 43598 15204 43650
rect 15148 43596 15204 43598
rect 14812 43484 14868 43540
rect 15260 43538 15316 43540
rect 15260 43486 15262 43538
rect 15262 43486 15314 43538
rect 15314 43486 15316 43538
rect 15260 43484 15316 43486
rect 15708 44210 15764 44212
rect 15708 44158 15710 44210
rect 15710 44158 15762 44210
rect 15762 44158 15764 44210
rect 15708 44156 15764 44158
rect 15596 43708 15652 43764
rect 15932 45500 15988 45556
rect 16044 45276 16100 45332
rect 15820 43596 15876 43652
rect 15596 43260 15652 43316
rect 15708 43148 15764 43204
rect 14812 42588 14868 42644
rect 15484 42924 15540 42980
rect 14812 40908 14868 40964
rect 14812 40236 14868 40292
rect 14924 41020 14980 41076
rect 14924 38892 14980 38948
rect 14028 38050 14084 38052
rect 14028 37998 14030 38050
rect 14030 37998 14082 38050
rect 14082 37998 14084 38050
rect 14028 37996 14084 37998
rect 13692 37884 13748 37940
rect 14700 38444 14756 38500
rect 14252 37266 14308 37268
rect 14252 37214 14254 37266
rect 14254 37214 14306 37266
rect 14306 37214 14308 37266
rect 14252 37212 14308 37214
rect 13468 36092 13524 36148
rect 14028 36370 14084 36372
rect 14028 36318 14030 36370
rect 14030 36318 14082 36370
rect 14082 36318 14084 36370
rect 14028 36316 14084 36318
rect 14028 35698 14084 35700
rect 14028 35646 14030 35698
rect 14030 35646 14082 35698
rect 14082 35646 14084 35698
rect 14028 35644 14084 35646
rect 14028 34860 14084 34916
rect 13804 34412 13860 34468
rect 14028 34354 14084 34356
rect 14028 34302 14030 34354
rect 14030 34302 14082 34354
rect 14082 34302 14084 34354
rect 14028 34300 14084 34302
rect 13468 34130 13524 34132
rect 13468 34078 13470 34130
rect 13470 34078 13522 34130
rect 13522 34078 13524 34130
rect 13468 34076 13524 34078
rect 13804 34130 13860 34132
rect 13804 34078 13806 34130
rect 13806 34078 13858 34130
rect 13858 34078 13860 34130
rect 13804 34076 13860 34078
rect 14364 36092 14420 36148
rect 15148 42364 15204 42420
rect 15148 40460 15204 40516
rect 15372 42252 15428 42308
rect 15820 42642 15876 42644
rect 15820 42590 15822 42642
rect 15822 42590 15874 42642
rect 15874 42590 15876 42642
rect 15820 42588 15876 42590
rect 16044 43932 16100 43988
rect 15932 42476 15988 42532
rect 16380 46898 16436 46900
rect 16380 46846 16382 46898
rect 16382 46846 16434 46898
rect 16434 46846 16436 46898
rect 16380 46844 16436 46846
rect 16604 47180 16660 47236
rect 16940 49138 16996 49140
rect 16940 49086 16942 49138
rect 16942 49086 16994 49138
rect 16994 49086 16996 49138
rect 16940 49084 16996 49086
rect 16828 48354 16884 48356
rect 16828 48302 16830 48354
rect 16830 48302 16882 48354
rect 16882 48302 16884 48354
rect 16828 48300 16884 48302
rect 17388 48636 17444 48692
rect 17164 47628 17220 47684
rect 17276 48188 17332 48244
rect 17164 47458 17220 47460
rect 17164 47406 17166 47458
rect 17166 47406 17218 47458
rect 17218 47406 17220 47458
rect 17164 47404 17220 47406
rect 17052 46844 17108 46900
rect 16828 46732 16884 46788
rect 16604 46284 16660 46340
rect 16828 46396 16884 46452
rect 16716 45164 16772 45220
rect 16716 44940 16772 44996
rect 16716 43932 16772 43988
rect 16716 43650 16772 43652
rect 16716 43598 16718 43650
rect 16718 43598 16770 43650
rect 16770 43598 16772 43650
rect 16716 43596 16772 43598
rect 16268 42812 16324 42868
rect 16156 42476 16212 42532
rect 16268 42252 16324 42308
rect 16492 42476 16548 42532
rect 16604 42194 16660 42196
rect 16604 42142 16606 42194
rect 16606 42142 16658 42194
rect 16658 42142 16660 42194
rect 16604 42140 16660 42142
rect 16044 41970 16100 41972
rect 16044 41918 16046 41970
rect 16046 41918 16098 41970
rect 16098 41918 16100 41970
rect 16044 41916 16100 41918
rect 15708 41804 15764 41860
rect 15596 41020 15652 41076
rect 15148 40290 15204 40292
rect 15148 40238 15150 40290
rect 15150 40238 15202 40290
rect 15202 40238 15204 40290
rect 15148 40236 15204 40238
rect 15820 40402 15876 40404
rect 15820 40350 15822 40402
rect 15822 40350 15874 40402
rect 15874 40350 15876 40402
rect 15820 40348 15876 40350
rect 15932 39506 15988 39508
rect 15932 39454 15934 39506
rect 15934 39454 15986 39506
rect 15986 39454 15988 39506
rect 15932 39452 15988 39454
rect 15484 39228 15540 39284
rect 15036 36428 15092 36484
rect 15148 37772 15204 37828
rect 15036 36092 15092 36148
rect 14812 35644 14868 35700
rect 14924 34972 14980 35028
rect 14700 34524 14756 34580
rect 15372 38108 15428 38164
rect 15708 39058 15764 39060
rect 15708 39006 15710 39058
rect 15710 39006 15762 39058
rect 15762 39006 15764 39058
rect 15708 39004 15764 39006
rect 15596 37996 15652 38052
rect 15820 37660 15876 37716
rect 15596 37436 15652 37492
rect 15484 36370 15540 36372
rect 15484 36318 15486 36370
rect 15486 36318 15538 36370
rect 15538 36318 15540 36370
rect 15484 36316 15540 36318
rect 15708 36316 15764 36372
rect 15596 35586 15652 35588
rect 15596 35534 15598 35586
rect 15598 35534 15650 35586
rect 15650 35534 15652 35586
rect 15596 35532 15652 35534
rect 15260 35308 15316 35364
rect 15596 35308 15652 35364
rect 15708 35026 15764 35028
rect 15708 34974 15710 35026
rect 15710 34974 15762 35026
rect 15762 34974 15764 35026
rect 15708 34972 15764 34974
rect 15820 34802 15876 34804
rect 15820 34750 15822 34802
rect 15822 34750 15874 34802
rect 15874 34750 15876 34802
rect 15820 34748 15876 34750
rect 15708 34354 15764 34356
rect 15708 34302 15710 34354
rect 15710 34302 15762 34354
rect 15762 34302 15764 34354
rect 15708 34300 15764 34302
rect 14252 33964 14308 34020
rect 14364 34076 14420 34132
rect 14140 33740 14196 33796
rect 14028 33628 14084 33684
rect 13356 33516 13412 33572
rect 13804 33292 13860 33348
rect 12572 32450 12628 32452
rect 12572 32398 12574 32450
rect 12574 32398 12626 32450
rect 12626 32398 12628 32450
rect 12572 32396 12628 32398
rect 12124 31948 12180 32004
rect 11452 31500 11508 31556
rect 11116 30882 11172 30884
rect 11116 30830 11118 30882
rect 11118 30830 11170 30882
rect 11170 30830 11172 30882
rect 11116 30828 11172 30830
rect 12012 30882 12068 30884
rect 12012 30830 12014 30882
rect 12014 30830 12066 30882
rect 12066 30830 12068 30882
rect 12012 30828 12068 30830
rect 14028 33122 14084 33124
rect 14028 33070 14030 33122
rect 14030 33070 14082 33122
rect 14082 33070 14084 33122
rect 14028 33068 14084 33070
rect 14140 32786 14196 32788
rect 14140 32734 14142 32786
rect 14142 32734 14194 32786
rect 14194 32734 14196 32786
rect 14140 32732 14196 32734
rect 13580 31724 13636 31780
rect 13020 31554 13076 31556
rect 13020 31502 13022 31554
rect 13022 31502 13074 31554
rect 13074 31502 13076 31554
rect 13020 31500 13076 31502
rect 13020 31276 13076 31332
rect 12796 30492 12852 30548
rect 11452 30156 11508 30212
rect 11900 30210 11956 30212
rect 11900 30158 11902 30210
rect 11902 30158 11954 30210
rect 11954 30158 11956 30210
rect 11900 30156 11956 30158
rect 11564 30044 11620 30100
rect 10556 29932 10612 29988
rect 11116 29986 11172 29988
rect 11116 29934 11118 29986
rect 11118 29934 11170 29986
rect 11170 29934 11172 29986
rect 11116 29932 11172 29934
rect 9996 24108 10052 24164
rect 10444 29426 10500 29428
rect 10444 29374 10446 29426
rect 10446 29374 10498 29426
rect 10498 29374 10500 29426
rect 10444 29372 10500 29374
rect 10332 28082 10388 28084
rect 10332 28030 10334 28082
rect 10334 28030 10386 28082
rect 10386 28030 10388 28082
rect 10332 28028 10388 28030
rect 10108 22652 10164 22708
rect 11452 29426 11508 29428
rect 11452 29374 11454 29426
rect 11454 29374 11506 29426
rect 11506 29374 11508 29426
rect 11452 29372 11508 29374
rect 11340 27858 11396 27860
rect 11340 27806 11342 27858
rect 11342 27806 11394 27858
rect 11394 27806 11396 27858
rect 11340 27804 11396 27806
rect 11340 27356 11396 27412
rect 12908 30098 12964 30100
rect 12908 30046 12910 30098
rect 12910 30046 12962 30098
rect 12962 30046 12964 30098
rect 12908 30044 12964 30046
rect 12348 29986 12404 29988
rect 12348 29934 12350 29986
rect 12350 29934 12402 29986
rect 12402 29934 12404 29986
rect 12348 29932 12404 29934
rect 13580 30940 13636 30996
rect 14588 33964 14644 34020
rect 14252 31836 14308 31892
rect 14812 33628 14868 33684
rect 16492 41916 16548 41972
rect 16604 41692 16660 41748
rect 16940 46674 16996 46676
rect 16940 46622 16942 46674
rect 16942 46622 16994 46674
rect 16994 46622 16996 46674
rect 16940 46620 16996 46622
rect 16940 46284 16996 46340
rect 17052 45890 17108 45892
rect 17052 45838 17054 45890
rect 17054 45838 17106 45890
rect 17106 45838 17108 45890
rect 17052 45836 17108 45838
rect 16940 45106 16996 45108
rect 16940 45054 16942 45106
rect 16942 45054 16994 45106
rect 16994 45054 16996 45106
rect 16940 45052 16996 45054
rect 16940 43708 16996 43764
rect 16940 43538 16996 43540
rect 16940 43486 16942 43538
rect 16942 43486 16994 43538
rect 16994 43486 16996 43538
rect 16940 43484 16996 43486
rect 16940 42866 16996 42868
rect 16940 42814 16942 42866
rect 16942 42814 16994 42866
rect 16994 42814 16996 42866
rect 16940 42812 16996 42814
rect 17612 51378 17668 51380
rect 17612 51326 17614 51378
rect 17614 51326 17666 51378
rect 17666 51326 17668 51378
rect 17612 51324 17668 51326
rect 17612 49868 17668 49924
rect 17948 53116 18004 53172
rect 18396 55074 18452 55076
rect 18396 55022 18398 55074
rect 18398 55022 18450 55074
rect 18450 55022 18452 55074
rect 18396 55020 18452 55022
rect 19068 54572 19124 54628
rect 19404 55074 19460 55076
rect 19404 55022 19406 55074
rect 19406 55022 19458 55074
rect 19458 55022 19460 55074
rect 19404 55020 19460 55022
rect 18620 54290 18676 54292
rect 18620 54238 18622 54290
rect 18622 54238 18674 54290
rect 18674 54238 18676 54290
rect 18620 54236 18676 54238
rect 18844 54012 18900 54068
rect 18284 53564 18340 53620
rect 18844 53618 18900 53620
rect 18844 53566 18846 53618
rect 18846 53566 18898 53618
rect 18898 53566 18900 53618
rect 18844 53564 18900 53566
rect 18396 53170 18452 53172
rect 18396 53118 18398 53170
rect 18398 53118 18450 53170
rect 18450 53118 18452 53170
rect 18396 53116 18452 53118
rect 18172 52556 18228 52612
rect 17948 52444 18004 52500
rect 18508 52668 18564 52724
rect 18396 52332 18452 52388
rect 18172 51938 18228 51940
rect 18172 51886 18174 51938
rect 18174 51886 18226 51938
rect 18226 51886 18228 51938
rect 18172 51884 18228 51886
rect 18284 51772 18340 51828
rect 17948 51602 18004 51604
rect 17948 51550 17950 51602
rect 17950 51550 18002 51602
rect 18002 51550 18004 51602
rect 17948 51548 18004 51550
rect 18172 51378 18228 51380
rect 18172 51326 18174 51378
rect 18174 51326 18226 51378
rect 18226 51326 18228 51378
rect 18172 51324 18228 51326
rect 17724 50316 17780 50372
rect 17724 48972 17780 49028
rect 18284 50482 18340 50484
rect 18284 50430 18286 50482
rect 18286 50430 18338 50482
rect 18338 50430 18340 50482
rect 18284 50428 18340 50430
rect 18508 49756 18564 49812
rect 17724 48242 17780 48244
rect 17724 48190 17726 48242
rect 17726 48190 17778 48242
rect 17778 48190 17780 48242
rect 17724 48188 17780 48190
rect 17836 48300 17892 48356
rect 17612 47516 17668 47572
rect 17500 47458 17556 47460
rect 17500 47406 17502 47458
rect 17502 47406 17554 47458
rect 17554 47406 17556 47458
rect 17500 47404 17556 47406
rect 17388 46844 17444 46900
rect 17500 47180 17556 47236
rect 17612 46844 17668 46900
rect 17500 46284 17556 46340
rect 17500 45164 17556 45220
rect 17500 44380 17556 44436
rect 17388 44098 17444 44100
rect 17388 44046 17390 44098
rect 17390 44046 17442 44098
rect 17442 44046 17444 44098
rect 17388 44044 17444 44046
rect 17500 43820 17556 43876
rect 18620 49644 18676 49700
rect 18508 49308 18564 49364
rect 18620 49138 18676 49140
rect 18620 49086 18622 49138
rect 18622 49086 18674 49138
rect 18674 49086 18676 49138
rect 18620 49084 18676 49086
rect 18508 48972 18564 49028
rect 18620 48802 18676 48804
rect 18620 48750 18622 48802
rect 18622 48750 18674 48802
rect 18674 48750 18676 48802
rect 18620 48748 18676 48750
rect 18508 48524 18564 48580
rect 18844 52444 18900 52500
rect 19180 53506 19236 53508
rect 19180 53454 19182 53506
rect 19182 53454 19234 53506
rect 19234 53454 19236 53506
rect 19180 53452 19236 53454
rect 18956 51548 19012 51604
rect 19180 51996 19236 52052
rect 18956 51100 19012 51156
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20860 54908 20916 54964
rect 20044 54852 20100 54854
rect 20412 54738 20468 54740
rect 20412 54686 20414 54738
rect 20414 54686 20466 54738
rect 20466 54686 20468 54738
rect 20412 54684 20468 54686
rect 20748 54514 20804 54516
rect 20748 54462 20750 54514
rect 20750 54462 20802 54514
rect 20802 54462 20804 54514
rect 20748 54460 20804 54462
rect 19964 53730 20020 53732
rect 19964 53678 19966 53730
rect 19966 53678 20018 53730
rect 20018 53678 20020 53730
rect 19964 53676 20020 53678
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19404 52386 19460 52388
rect 19404 52334 19406 52386
rect 19406 52334 19458 52386
rect 19458 52334 19460 52386
rect 19404 52332 19460 52334
rect 19292 51772 19348 51828
rect 20188 52834 20244 52836
rect 20188 52782 20190 52834
rect 20190 52782 20242 52834
rect 20242 52782 20244 52834
rect 20188 52780 20244 52782
rect 20076 52444 20132 52500
rect 19852 51996 19908 52052
rect 20188 52108 20244 52164
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19180 50876 19236 50932
rect 19404 50652 19460 50708
rect 20524 53170 20580 53172
rect 20524 53118 20526 53170
rect 20526 53118 20578 53170
rect 20578 53118 20580 53170
rect 20524 53116 20580 53118
rect 20524 52556 20580 52612
rect 20636 52892 20692 52948
rect 20524 52220 20580 52276
rect 20636 52108 20692 52164
rect 21084 55244 21140 55300
rect 20972 53116 21028 53172
rect 20860 52162 20916 52164
rect 20860 52110 20862 52162
rect 20862 52110 20914 52162
rect 20914 52110 20916 52162
rect 20860 52108 20916 52110
rect 22540 56082 22596 56084
rect 22540 56030 22542 56082
rect 22542 56030 22594 56082
rect 22594 56030 22596 56082
rect 22540 56028 22596 56030
rect 22652 55858 22708 55860
rect 22652 55806 22654 55858
rect 22654 55806 22706 55858
rect 22706 55806 22708 55858
rect 22652 55804 22708 55806
rect 22204 55132 22260 55188
rect 22092 55020 22148 55076
rect 22316 55074 22372 55076
rect 22316 55022 22318 55074
rect 22318 55022 22370 55074
rect 22370 55022 22372 55074
rect 22316 55020 22372 55022
rect 25900 57148 25956 57204
rect 24444 56082 24500 56084
rect 24444 56030 24446 56082
rect 24446 56030 24498 56082
rect 24498 56030 24500 56082
rect 24444 56028 24500 56030
rect 23548 55356 23604 55412
rect 22764 54908 22820 54964
rect 22204 54684 22260 54740
rect 21196 52946 21252 52948
rect 21196 52894 21198 52946
rect 21198 52894 21250 52946
rect 21250 52894 21252 52946
rect 21196 52892 21252 52894
rect 21308 54348 21364 54404
rect 21644 54124 21700 54180
rect 21868 54348 21924 54404
rect 22092 54460 22148 54516
rect 20748 51660 20804 51716
rect 21420 52780 21476 52836
rect 20524 51602 20580 51604
rect 20524 51550 20526 51602
rect 20526 51550 20578 51602
rect 20578 51550 20580 51602
rect 20524 51548 20580 51550
rect 20860 51324 20916 51380
rect 20972 51548 21028 51604
rect 20188 50876 20244 50932
rect 20076 50652 20132 50708
rect 18844 49980 18900 50036
rect 18956 49868 19012 49924
rect 18844 49698 18900 49700
rect 18844 49646 18846 49698
rect 18846 49646 18898 49698
rect 18898 49646 18900 49698
rect 18844 49644 18900 49646
rect 19628 50540 19684 50596
rect 19404 49868 19460 49924
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19852 50034 19908 50036
rect 19852 49982 19854 50034
rect 19854 49982 19906 50034
rect 19906 49982 19908 50034
rect 19852 49980 19908 49982
rect 20076 49810 20132 49812
rect 20076 49758 20078 49810
rect 20078 49758 20130 49810
rect 20130 49758 20132 49810
rect 20076 49756 20132 49758
rect 19628 49532 19684 49588
rect 18844 49026 18900 49028
rect 18844 48974 18846 49026
rect 18846 48974 18898 49026
rect 18898 48974 18900 49026
rect 18844 48972 18900 48974
rect 19068 49420 19124 49476
rect 18172 48354 18228 48356
rect 18172 48302 18174 48354
rect 18174 48302 18226 48354
rect 18226 48302 18228 48354
rect 18172 48300 18228 48302
rect 18060 46844 18116 46900
rect 18172 47628 18228 47684
rect 17948 46060 18004 46116
rect 17948 45612 18004 45668
rect 17724 44380 17780 44436
rect 17724 44044 17780 44100
rect 17724 43538 17780 43540
rect 17724 43486 17726 43538
rect 17726 43486 17778 43538
rect 17778 43486 17780 43538
rect 17724 43484 17780 43486
rect 18060 44940 18116 44996
rect 18396 48242 18452 48244
rect 18396 48190 18398 48242
rect 18398 48190 18450 48242
rect 18450 48190 18452 48242
rect 18396 48188 18452 48190
rect 19068 48300 19124 48356
rect 19180 49308 19236 49364
rect 18732 48076 18788 48132
rect 18396 46674 18452 46676
rect 18396 46622 18398 46674
rect 18398 46622 18450 46674
rect 18450 46622 18452 46674
rect 18396 46620 18452 46622
rect 18284 46508 18340 46564
rect 18620 46396 18676 46452
rect 18284 45500 18340 45556
rect 18284 44044 18340 44100
rect 18956 47740 19012 47796
rect 19068 46898 19124 46900
rect 19068 46846 19070 46898
rect 19070 46846 19122 46898
rect 19122 46846 19124 46898
rect 19068 46844 19124 46846
rect 19628 49308 19684 49364
rect 19404 49084 19460 49140
rect 19292 48636 19348 48692
rect 19292 48076 19348 48132
rect 19180 46060 19236 46116
rect 19292 47628 19348 47684
rect 18508 44828 18564 44884
rect 18508 43596 18564 43652
rect 18844 45500 18900 45556
rect 18844 45052 18900 45108
rect 18844 44828 18900 44884
rect 19068 44716 19124 44772
rect 20412 49868 20468 49924
rect 19964 49084 20020 49140
rect 20188 49084 20244 49140
rect 19516 48636 19572 48692
rect 19836 48634 19892 48636
rect 19628 48524 19684 48580
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19964 48300 20020 48356
rect 19852 47964 19908 48020
rect 19852 47628 19908 47684
rect 19628 47458 19684 47460
rect 19628 47406 19630 47458
rect 19630 47406 19682 47458
rect 19682 47406 19684 47458
rect 19628 47404 19684 47406
rect 20076 48076 20132 48132
rect 20188 47628 20244 47684
rect 20300 48748 20356 48804
rect 20524 48524 20580 48580
rect 20748 49644 20804 49700
rect 20748 48860 20804 48916
rect 20524 47964 20580 48020
rect 20524 47682 20580 47684
rect 20524 47630 20526 47682
rect 20526 47630 20578 47682
rect 20578 47630 20580 47682
rect 20524 47628 20580 47630
rect 19964 47292 20020 47348
rect 19740 47234 19796 47236
rect 19740 47182 19742 47234
rect 19742 47182 19794 47234
rect 19794 47182 19796 47234
rect 19740 47180 19796 47182
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19964 46844 20020 46900
rect 19628 46674 19684 46676
rect 19628 46622 19630 46674
rect 19630 46622 19682 46674
rect 19682 46622 19684 46674
rect 19628 46620 19684 46622
rect 19740 46562 19796 46564
rect 19740 46510 19742 46562
rect 19742 46510 19794 46562
rect 19794 46510 19796 46562
rect 19740 46508 19796 46510
rect 20076 46396 20132 46452
rect 20300 46060 20356 46116
rect 19516 45612 19572 45668
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19404 45164 19460 45220
rect 19740 45052 19796 45108
rect 19628 44828 19684 44884
rect 18956 44492 19012 44548
rect 19068 44380 19124 44436
rect 18844 43932 18900 43988
rect 18620 43820 18676 43876
rect 18284 43484 18340 43540
rect 17500 42924 17556 42980
rect 18060 42978 18116 42980
rect 18060 42926 18062 42978
rect 18062 42926 18114 42978
rect 18114 42926 18116 42978
rect 18060 42924 18116 42926
rect 17388 42530 17444 42532
rect 17388 42478 17390 42530
rect 17390 42478 17442 42530
rect 17442 42478 17444 42530
rect 17388 42476 17444 42478
rect 16940 41970 16996 41972
rect 16940 41918 16942 41970
rect 16942 41918 16994 41970
rect 16994 41918 16996 41970
rect 16940 41916 16996 41918
rect 16604 40796 16660 40852
rect 16156 39676 16212 39732
rect 16380 40460 16436 40516
rect 16604 40460 16660 40516
rect 16380 38946 16436 38948
rect 16380 38894 16382 38946
rect 16382 38894 16434 38946
rect 16434 38894 16436 38946
rect 16380 38892 16436 38894
rect 16492 39004 16548 39060
rect 16044 38556 16100 38612
rect 16044 37938 16100 37940
rect 16044 37886 16046 37938
rect 16046 37886 16098 37938
rect 16098 37886 16100 37938
rect 16044 37884 16100 37886
rect 16268 36482 16324 36484
rect 16268 36430 16270 36482
rect 16270 36430 16322 36482
rect 16322 36430 16324 36482
rect 16268 36428 16324 36430
rect 16156 36370 16212 36372
rect 16156 36318 16158 36370
rect 16158 36318 16210 36370
rect 16210 36318 16212 36370
rect 16156 36316 16212 36318
rect 16268 36092 16324 36148
rect 16268 35756 16324 35812
rect 16044 35420 16100 35476
rect 16044 34748 16100 34804
rect 16268 34748 16324 34804
rect 16156 34524 16212 34580
rect 16044 34076 16100 34132
rect 14924 33346 14980 33348
rect 14924 33294 14926 33346
rect 14926 33294 14978 33346
rect 14978 33294 14980 33346
rect 14924 33292 14980 33294
rect 15260 32956 15316 33012
rect 15148 32786 15204 32788
rect 15148 32734 15150 32786
rect 15150 32734 15202 32786
rect 15202 32734 15204 32786
rect 15148 32732 15204 32734
rect 15260 32396 15316 32452
rect 15708 32396 15764 32452
rect 14924 31890 14980 31892
rect 14924 31838 14926 31890
rect 14926 31838 14978 31890
rect 14978 31838 14980 31890
rect 14924 31836 14980 31838
rect 14140 31666 14196 31668
rect 14140 31614 14142 31666
rect 14142 31614 14194 31666
rect 14194 31614 14196 31666
rect 14140 31612 14196 31614
rect 14476 31724 14532 31780
rect 14140 31218 14196 31220
rect 14140 31166 14142 31218
rect 14142 31166 14194 31218
rect 14194 31166 14196 31218
rect 14140 31164 14196 31166
rect 14028 30940 14084 30996
rect 11676 29314 11732 29316
rect 11676 29262 11678 29314
rect 11678 29262 11730 29314
rect 11730 29262 11732 29314
rect 11676 29260 11732 29262
rect 12348 29148 12404 29204
rect 13356 28924 13412 28980
rect 13692 28476 13748 28532
rect 14028 29484 14084 29540
rect 15484 31218 15540 31220
rect 15484 31166 15486 31218
rect 15486 31166 15538 31218
rect 15538 31166 15540 31218
rect 15484 31164 15540 31166
rect 14588 31052 14644 31108
rect 15260 31106 15316 31108
rect 15260 31054 15262 31106
rect 15262 31054 15314 31106
rect 15314 31054 15316 31106
rect 15260 31052 15316 31054
rect 15036 30828 15092 30884
rect 14700 30434 14756 30436
rect 14700 30382 14702 30434
rect 14702 30382 14754 30434
rect 14754 30382 14756 30434
rect 14700 30380 14756 30382
rect 15148 30380 15204 30436
rect 15260 30828 15316 30884
rect 14924 30210 14980 30212
rect 14924 30158 14926 30210
rect 14926 30158 14978 30210
rect 14978 30158 14980 30210
rect 14924 30156 14980 30158
rect 14252 28028 14308 28084
rect 13468 27356 13524 27412
rect 13020 26962 13076 26964
rect 13020 26910 13022 26962
rect 13022 26910 13074 26962
rect 13074 26910 13076 26962
rect 13020 26908 13076 26910
rect 11676 24220 11732 24276
rect 13804 26962 13860 26964
rect 13804 26910 13806 26962
rect 13806 26910 13858 26962
rect 13858 26910 13860 26962
rect 13804 26908 13860 26910
rect 14812 29426 14868 29428
rect 14812 29374 14814 29426
rect 14814 29374 14866 29426
rect 14866 29374 14868 29426
rect 14812 29372 14868 29374
rect 14924 29260 14980 29316
rect 14700 28924 14756 28980
rect 14476 28642 14532 28644
rect 14476 28590 14478 28642
rect 14478 28590 14530 28642
rect 14530 28590 14532 28642
rect 14476 28588 14532 28590
rect 14588 27804 14644 27860
rect 15148 27356 15204 27412
rect 15708 30268 15764 30324
rect 15596 30210 15652 30212
rect 15596 30158 15598 30210
rect 15598 30158 15650 30210
rect 15650 30158 15652 30210
rect 15596 30156 15652 30158
rect 15932 32956 15988 33012
rect 15932 32732 15988 32788
rect 16156 33234 16212 33236
rect 16156 33182 16158 33234
rect 16158 33182 16210 33234
rect 16210 33182 16212 33234
rect 16156 33180 16212 33182
rect 16268 32956 16324 33012
rect 16604 37996 16660 38052
rect 16492 37938 16548 37940
rect 16492 37886 16494 37938
rect 16494 37886 16546 37938
rect 16546 37886 16548 37938
rect 16492 37884 16548 37886
rect 16604 37772 16660 37828
rect 17164 41132 17220 41188
rect 16940 40684 16996 40740
rect 17164 40684 17220 40740
rect 17500 41916 17556 41972
rect 16940 40402 16996 40404
rect 16940 40350 16942 40402
rect 16942 40350 16994 40402
rect 16994 40350 16996 40402
rect 16940 40348 16996 40350
rect 16940 39842 16996 39844
rect 16940 39790 16942 39842
rect 16942 39790 16994 39842
rect 16994 39790 16996 39842
rect 16940 39788 16996 39790
rect 17052 39676 17108 39732
rect 16940 38834 16996 38836
rect 16940 38782 16942 38834
rect 16942 38782 16994 38834
rect 16994 38782 16996 38834
rect 16940 38780 16996 38782
rect 16716 37436 16772 37492
rect 16604 36876 16660 36932
rect 16492 35308 16548 35364
rect 16716 35308 16772 35364
rect 16604 34802 16660 34804
rect 16604 34750 16606 34802
rect 16606 34750 16658 34802
rect 16658 34750 16660 34802
rect 16604 34748 16660 34750
rect 16604 33292 16660 33348
rect 16492 32956 16548 33012
rect 16940 37938 16996 37940
rect 16940 37886 16942 37938
rect 16942 37886 16994 37938
rect 16994 37886 16996 37938
rect 16940 37884 16996 37886
rect 16940 37490 16996 37492
rect 16940 37438 16942 37490
rect 16942 37438 16994 37490
rect 16994 37438 16996 37490
rect 16940 37436 16996 37438
rect 17164 36540 17220 36596
rect 17164 36204 17220 36260
rect 17052 35756 17108 35812
rect 16940 35698 16996 35700
rect 16940 35646 16942 35698
rect 16942 35646 16994 35698
rect 16994 35646 16996 35698
rect 16940 35644 16996 35646
rect 16940 35308 16996 35364
rect 16940 34524 16996 34580
rect 16940 33346 16996 33348
rect 16940 33294 16942 33346
rect 16942 33294 16994 33346
rect 16994 33294 16996 33346
rect 16940 33292 16996 33294
rect 16604 32450 16660 32452
rect 16604 32398 16606 32450
rect 16606 32398 16658 32450
rect 16658 32398 16660 32450
rect 16604 32396 16660 32398
rect 17388 40684 17444 40740
rect 17724 42082 17780 42084
rect 17724 42030 17726 42082
rect 17726 42030 17778 42082
rect 17778 42030 17780 42082
rect 17724 42028 17780 42030
rect 17948 42588 18004 42644
rect 18060 42028 18116 42084
rect 17612 41692 17668 41748
rect 17612 41410 17668 41412
rect 17612 41358 17614 41410
rect 17614 41358 17666 41410
rect 17666 41358 17668 41410
rect 17612 41356 17668 41358
rect 17836 41020 17892 41076
rect 17948 40908 18004 40964
rect 17500 37996 17556 38052
rect 17836 39394 17892 39396
rect 17836 39342 17838 39394
rect 17838 39342 17890 39394
rect 17890 39342 17892 39394
rect 17836 39340 17892 39342
rect 17724 39004 17780 39060
rect 18396 42978 18452 42980
rect 18396 42926 18398 42978
rect 18398 42926 18450 42978
rect 18450 42926 18452 42978
rect 18396 42924 18452 42926
rect 18844 43650 18900 43652
rect 18844 43598 18846 43650
rect 18846 43598 18898 43650
rect 18898 43598 18900 43650
rect 18844 43596 18900 43598
rect 18620 42588 18676 42644
rect 18172 39676 18228 39732
rect 18396 42476 18452 42532
rect 18508 40962 18564 40964
rect 18508 40910 18510 40962
rect 18510 40910 18562 40962
rect 18562 40910 18564 40962
rect 18508 40908 18564 40910
rect 17724 38668 17780 38724
rect 18732 43036 18788 43092
rect 18956 42978 19012 42980
rect 18956 42926 18958 42978
rect 18958 42926 19010 42978
rect 19010 42926 19012 42978
rect 18956 42924 19012 42926
rect 19180 42754 19236 42756
rect 19180 42702 19182 42754
rect 19182 42702 19234 42754
rect 19234 42702 19236 42754
rect 19180 42700 19236 42702
rect 19404 43036 19460 43092
rect 20188 44546 20244 44548
rect 20188 44494 20190 44546
rect 20190 44494 20242 44546
rect 20242 44494 20244 44546
rect 20188 44492 20244 44494
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19740 43708 19796 43764
rect 20636 46620 20692 46676
rect 20524 45778 20580 45780
rect 20524 45726 20526 45778
rect 20526 45726 20578 45778
rect 20578 45726 20580 45778
rect 20524 45724 20580 45726
rect 21084 49196 21140 49252
rect 20860 48300 20916 48356
rect 20972 48524 21028 48580
rect 20748 45500 20804 45556
rect 20860 47740 20916 47796
rect 20636 45052 20692 45108
rect 21420 51772 21476 51828
rect 21308 51602 21364 51604
rect 21308 51550 21310 51602
rect 21310 51550 21362 51602
rect 21362 51550 21364 51602
rect 21308 51548 21364 51550
rect 21308 50428 21364 50484
rect 21532 50764 21588 50820
rect 23436 55132 23492 55188
rect 23212 55074 23268 55076
rect 23212 55022 23214 55074
rect 23214 55022 23266 55074
rect 23266 55022 23268 55074
rect 23212 55020 23268 55022
rect 23324 54908 23380 54964
rect 23884 55244 23940 55300
rect 23660 54796 23716 54852
rect 23436 53900 23492 53956
rect 23100 53788 23156 53844
rect 22428 53564 22484 53620
rect 21756 51772 21812 51828
rect 22092 51884 22148 51940
rect 21868 51266 21924 51268
rect 21868 51214 21870 51266
rect 21870 51214 21922 51266
rect 21922 51214 21924 51266
rect 21868 51212 21924 51214
rect 21644 50540 21700 50596
rect 21756 50876 21812 50932
rect 21420 49420 21476 49476
rect 21532 49084 21588 49140
rect 21644 48412 21700 48468
rect 21980 49756 22036 49812
rect 23436 53564 23492 53620
rect 22764 53506 22820 53508
rect 22764 53454 22766 53506
rect 22766 53454 22818 53506
rect 22818 53454 22820 53506
rect 22764 53452 22820 53454
rect 22988 53340 23044 53396
rect 22428 52780 22484 52836
rect 22316 52556 22372 52612
rect 23100 52834 23156 52836
rect 23100 52782 23102 52834
rect 23102 52782 23154 52834
rect 23154 52782 23156 52834
rect 23100 52780 23156 52782
rect 23324 52780 23380 52836
rect 22876 52050 22932 52052
rect 22876 51998 22878 52050
rect 22878 51998 22930 52050
rect 22930 51998 22932 52050
rect 22876 51996 22932 51998
rect 22764 51772 22820 51828
rect 22428 51378 22484 51380
rect 22428 51326 22430 51378
rect 22430 51326 22482 51378
rect 22482 51326 22484 51378
rect 22428 51324 22484 51326
rect 22316 50764 22372 50820
rect 22652 51266 22708 51268
rect 22652 51214 22654 51266
rect 22654 51214 22706 51266
rect 22706 51214 22708 51266
rect 22652 51212 22708 51214
rect 22764 50876 22820 50932
rect 23212 51324 23268 51380
rect 22876 50482 22932 50484
rect 22876 50430 22878 50482
rect 22878 50430 22930 50482
rect 22930 50430 22932 50482
rect 22876 50428 22932 50430
rect 23548 53170 23604 53172
rect 23548 53118 23550 53170
rect 23550 53118 23602 53170
rect 23602 53118 23604 53170
rect 23548 53116 23604 53118
rect 23548 52274 23604 52276
rect 23548 52222 23550 52274
rect 23550 52222 23602 52274
rect 23602 52222 23604 52274
rect 23548 52220 23604 52222
rect 23660 52108 23716 52164
rect 23436 51772 23492 51828
rect 23772 51884 23828 51940
rect 24220 55298 24276 55300
rect 24220 55246 24222 55298
rect 24222 55246 24274 55298
rect 24274 55246 24276 55298
rect 24220 55244 24276 55246
rect 25676 56082 25732 56084
rect 25676 56030 25678 56082
rect 25678 56030 25730 56082
rect 25730 56030 25732 56082
rect 25676 56028 25732 56030
rect 24892 55804 24948 55860
rect 25228 55298 25284 55300
rect 25228 55246 25230 55298
rect 25230 55246 25282 55298
rect 25282 55246 25284 55298
rect 25228 55244 25284 55246
rect 25788 55916 25844 55972
rect 26460 56252 26516 56308
rect 26124 56194 26180 56196
rect 26124 56142 26126 56194
rect 26126 56142 26178 56194
rect 26178 56142 26180 56194
rect 26124 56140 26180 56142
rect 25340 55132 25396 55188
rect 26012 55580 26068 55636
rect 23996 54460 24052 54516
rect 24108 53730 24164 53732
rect 24108 53678 24110 53730
rect 24110 53678 24162 53730
rect 24162 53678 24164 53730
rect 24108 53676 24164 53678
rect 23996 53618 24052 53620
rect 23996 53566 23998 53618
rect 23998 53566 24050 53618
rect 24050 53566 24052 53618
rect 23996 53564 24052 53566
rect 23884 51548 23940 51604
rect 23996 53116 24052 53172
rect 24108 52444 24164 52500
rect 24108 52162 24164 52164
rect 24108 52110 24110 52162
rect 24110 52110 24162 52162
rect 24162 52110 24164 52162
rect 24108 52108 24164 52110
rect 23660 51490 23716 51492
rect 23660 51438 23662 51490
rect 23662 51438 23714 51490
rect 23714 51438 23716 51490
rect 23660 51436 23716 51438
rect 23548 51324 23604 51380
rect 23884 51378 23940 51380
rect 23884 51326 23886 51378
rect 23886 51326 23938 51378
rect 23938 51326 23940 51378
rect 23884 51324 23940 51326
rect 23324 51100 23380 51156
rect 23212 50204 23268 50260
rect 23436 50876 23492 50932
rect 22316 50034 22372 50036
rect 22316 49982 22318 50034
rect 22318 49982 22370 50034
rect 22370 49982 22372 50034
rect 22316 49980 22372 49982
rect 23324 50034 23380 50036
rect 23324 49982 23326 50034
rect 23326 49982 23378 50034
rect 23378 49982 23380 50034
rect 23324 49980 23380 49982
rect 23212 49922 23268 49924
rect 23212 49870 23214 49922
rect 23214 49870 23266 49922
rect 23266 49870 23268 49922
rect 23212 49868 23268 49870
rect 22652 49810 22708 49812
rect 22652 49758 22654 49810
rect 22654 49758 22706 49810
rect 22706 49758 22708 49810
rect 22652 49756 22708 49758
rect 22204 49420 22260 49476
rect 22876 49420 22932 49476
rect 22204 49250 22260 49252
rect 22204 49198 22206 49250
rect 22206 49198 22258 49250
rect 22258 49198 22260 49250
rect 22204 49196 22260 49198
rect 22652 48860 22708 48916
rect 22540 48802 22596 48804
rect 22540 48750 22542 48802
rect 22542 48750 22594 48802
rect 22594 48750 22596 48802
rect 22540 48748 22596 48750
rect 22092 48412 22148 48468
rect 21756 48300 21812 48356
rect 21196 47740 21252 47796
rect 21308 47852 21364 47908
rect 21084 47628 21140 47684
rect 21644 48076 21700 48132
rect 22540 47682 22596 47684
rect 22540 47630 22542 47682
rect 22542 47630 22594 47682
rect 22594 47630 22596 47682
rect 22540 47628 22596 47630
rect 21868 46956 21924 47012
rect 21308 46844 21364 46900
rect 20972 46508 21028 46564
rect 20524 44828 20580 44884
rect 20412 43820 20468 43876
rect 19964 43484 20020 43540
rect 20300 43484 20356 43540
rect 19628 42924 19684 42980
rect 19852 43148 19908 43204
rect 19516 42812 19572 42868
rect 19740 42866 19796 42868
rect 19740 42814 19742 42866
rect 19742 42814 19794 42866
rect 19794 42814 19796 42866
rect 19740 42812 19796 42814
rect 20076 42588 20132 42644
rect 19292 42252 19348 42308
rect 18844 41970 18900 41972
rect 18844 41918 18846 41970
rect 18846 41918 18898 41970
rect 18898 41918 18900 41970
rect 18844 41916 18900 41918
rect 19068 41916 19124 41972
rect 18956 41356 19012 41412
rect 19516 41020 19572 41076
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19852 41468 19908 41524
rect 20300 41858 20356 41860
rect 20300 41806 20302 41858
rect 20302 41806 20354 41858
rect 20354 41806 20356 41858
rect 20300 41804 20356 41806
rect 20412 43260 20468 43316
rect 19964 41356 20020 41412
rect 20636 43650 20692 43652
rect 20636 43598 20638 43650
rect 20638 43598 20690 43650
rect 20690 43598 20692 43650
rect 20636 43596 20692 43598
rect 20524 43036 20580 43092
rect 21308 44492 21364 44548
rect 21308 43932 21364 43988
rect 21084 43426 21140 43428
rect 21084 43374 21086 43426
rect 21086 43374 21138 43426
rect 21138 43374 21140 43426
rect 21084 43372 21140 43374
rect 20748 41692 20804 41748
rect 20524 41580 20580 41636
rect 20748 41356 20804 41412
rect 20636 41298 20692 41300
rect 20636 41246 20638 41298
rect 20638 41246 20690 41298
rect 20690 41246 20692 41298
rect 20636 41244 20692 41246
rect 19740 40908 19796 40964
rect 19516 40796 19572 40852
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 20412 41186 20468 41188
rect 20412 41134 20414 41186
rect 20414 41134 20466 41186
rect 20466 41134 20468 41186
rect 20412 41132 20468 41134
rect 20076 40514 20132 40516
rect 20076 40462 20078 40514
rect 20078 40462 20130 40514
rect 20130 40462 20132 40514
rect 20076 40460 20132 40462
rect 20412 40402 20468 40404
rect 20412 40350 20414 40402
rect 20414 40350 20466 40402
rect 20466 40350 20468 40402
rect 20412 40348 20468 40350
rect 18620 39116 18676 39172
rect 17500 37436 17556 37492
rect 17836 37212 17892 37268
rect 17724 36764 17780 36820
rect 17724 36540 17780 36596
rect 18732 38162 18788 38164
rect 18732 38110 18734 38162
rect 18734 38110 18786 38162
rect 18786 38110 18788 38162
rect 18732 38108 18788 38110
rect 19068 40236 19124 40292
rect 19068 38220 19124 38276
rect 18956 37772 19012 37828
rect 18620 37266 18676 37268
rect 18620 37214 18622 37266
rect 18622 37214 18674 37266
rect 18674 37214 18676 37266
rect 18620 37212 18676 37214
rect 17388 36092 17444 36148
rect 17276 35868 17332 35924
rect 17724 35810 17780 35812
rect 17724 35758 17726 35810
rect 17726 35758 17778 35810
rect 17778 35758 17780 35810
rect 17724 35756 17780 35758
rect 18284 36204 18340 36260
rect 17500 35308 17556 35364
rect 18172 35644 18228 35700
rect 17388 33180 17444 33236
rect 17276 32620 17332 32676
rect 16940 31724 16996 31780
rect 16380 30940 16436 30996
rect 16044 30882 16100 30884
rect 16044 30830 16046 30882
rect 16046 30830 16098 30882
rect 16098 30830 16100 30882
rect 16044 30828 16100 30830
rect 15820 29708 15876 29764
rect 16268 29484 16324 29540
rect 16940 30380 16996 30436
rect 16380 30156 16436 30212
rect 15596 29426 15652 29428
rect 15596 29374 15598 29426
rect 15598 29374 15650 29426
rect 15650 29374 15652 29426
rect 15596 29372 15652 29374
rect 17388 32060 17444 32116
rect 17948 34242 18004 34244
rect 17948 34190 17950 34242
rect 17950 34190 18002 34242
rect 18002 34190 18004 34242
rect 17948 34188 18004 34190
rect 17612 33292 17668 33348
rect 18508 36370 18564 36372
rect 18508 36318 18510 36370
rect 18510 36318 18562 36370
rect 18562 36318 18564 36370
rect 18508 36316 18564 36318
rect 18396 35308 18452 35364
rect 18396 34802 18452 34804
rect 18396 34750 18398 34802
rect 18398 34750 18450 34802
rect 18450 34750 18452 34802
rect 18396 34748 18452 34750
rect 18844 35980 18900 36036
rect 18732 35196 18788 35252
rect 18844 35644 18900 35700
rect 18284 34300 18340 34356
rect 18732 34524 18788 34580
rect 18620 34242 18676 34244
rect 18620 34190 18622 34242
rect 18622 34190 18674 34242
rect 18674 34190 18676 34242
rect 18620 34188 18676 34190
rect 19292 37938 19348 37940
rect 19292 37886 19294 37938
rect 19294 37886 19346 37938
rect 19346 37886 19348 37938
rect 19292 37884 19348 37886
rect 20524 40124 20580 40180
rect 19404 37212 19460 37268
rect 19516 40012 19572 40068
rect 19068 36258 19124 36260
rect 19068 36206 19070 36258
rect 19070 36206 19122 36258
rect 19122 36206 19124 36258
rect 19068 36204 19124 36206
rect 19068 35756 19124 35812
rect 19180 35532 19236 35588
rect 19404 35698 19460 35700
rect 19404 35646 19406 35698
rect 19406 35646 19458 35698
rect 19458 35646 19460 35698
rect 19404 35644 19460 35646
rect 19292 34524 19348 34580
rect 20860 40348 20916 40404
rect 21532 45330 21588 45332
rect 21532 45278 21534 45330
rect 21534 45278 21586 45330
rect 21586 45278 21588 45330
rect 21532 45276 21588 45278
rect 21868 45218 21924 45220
rect 21868 45166 21870 45218
rect 21870 45166 21922 45218
rect 21922 45166 21924 45218
rect 21868 45164 21924 45166
rect 21420 43708 21476 43764
rect 21532 43538 21588 43540
rect 21532 43486 21534 43538
rect 21534 43486 21586 43538
rect 21586 43486 21588 43538
rect 21532 43484 21588 43486
rect 22540 46898 22596 46900
rect 22540 46846 22542 46898
rect 22542 46846 22594 46898
rect 22594 46846 22596 46898
rect 22540 46844 22596 46846
rect 22428 45164 22484 45220
rect 21868 44322 21924 44324
rect 21868 44270 21870 44322
rect 21870 44270 21922 44322
rect 21922 44270 21924 44322
rect 21868 44268 21924 44270
rect 22092 44044 22148 44100
rect 21980 43708 22036 43764
rect 22092 43650 22148 43652
rect 22092 43598 22094 43650
rect 22094 43598 22146 43650
rect 22146 43598 22148 43650
rect 22092 43596 22148 43598
rect 21644 43260 21700 43316
rect 21532 43148 21588 43204
rect 21420 42028 21476 42084
rect 21196 41858 21252 41860
rect 21196 41806 21198 41858
rect 21198 41806 21250 41858
rect 21250 41806 21252 41858
rect 21196 41804 21252 41806
rect 21084 41468 21140 41524
rect 21308 41468 21364 41524
rect 20972 40236 21028 40292
rect 20972 39900 21028 39956
rect 19852 39842 19908 39844
rect 19852 39790 19854 39842
rect 19854 39790 19906 39842
rect 19906 39790 19908 39842
rect 19852 39788 19908 39790
rect 19628 39506 19684 39508
rect 19628 39454 19630 39506
rect 19630 39454 19682 39506
rect 19682 39454 19684 39506
rect 19628 39452 19684 39454
rect 19628 39228 19684 39284
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 20972 38892 21028 38948
rect 20748 38834 20804 38836
rect 20748 38782 20750 38834
rect 20750 38782 20802 38834
rect 20802 38782 20804 38834
rect 20748 38780 20804 38782
rect 20636 38668 20692 38724
rect 20300 38108 20356 38164
rect 19628 37938 19684 37940
rect 19628 37886 19630 37938
rect 19630 37886 19682 37938
rect 19682 37886 19684 37938
rect 19628 37884 19684 37886
rect 20636 37884 20692 37940
rect 19628 37660 19684 37716
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20860 37938 20916 37940
rect 20860 37886 20862 37938
rect 20862 37886 20914 37938
rect 20914 37886 20916 37938
rect 20860 37884 20916 37886
rect 20636 37324 20692 37380
rect 20076 37266 20132 37268
rect 20076 37214 20078 37266
rect 20078 37214 20130 37266
rect 20130 37214 20132 37266
rect 20076 37212 20132 37214
rect 19852 36764 19908 36820
rect 19628 36370 19684 36372
rect 19628 36318 19630 36370
rect 19630 36318 19682 36370
rect 19682 36318 19684 36370
rect 19628 36316 19684 36318
rect 19852 36204 19908 36260
rect 20524 36204 20580 36260
rect 21420 40348 21476 40404
rect 20972 36540 21028 36596
rect 21420 39900 21476 39956
rect 21420 39676 21476 39732
rect 21420 38722 21476 38724
rect 21420 38670 21422 38722
rect 21422 38670 21474 38722
rect 21474 38670 21476 38722
rect 21420 38668 21476 38670
rect 19628 36092 19684 36148
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 20860 36258 20916 36260
rect 20860 36206 20862 36258
rect 20862 36206 20914 36258
rect 20914 36206 20916 36258
rect 20860 36204 20916 36206
rect 19964 35474 20020 35476
rect 19964 35422 19966 35474
rect 19966 35422 20018 35474
rect 20018 35422 20020 35474
rect 19964 35420 20020 35422
rect 20076 34748 20132 34804
rect 20524 35196 20580 35252
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19740 34130 19796 34132
rect 19740 34078 19742 34130
rect 19742 34078 19794 34130
rect 19794 34078 19796 34130
rect 19740 34076 19796 34078
rect 20188 34076 20244 34132
rect 21084 35196 21140 35252
rect 19292 32844 19348 32900
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 18172 32786 18228 32788
rect 18172 32734 18174 32786
rect 18174 32734 18226 32786
rect 18226 32734 18228 32786
rect 18172 32732 18228 32734
rect 18956 32732 19012 32788
rect 19516 32562 19572 32564
rect 19516 32510 19518 32562
rect 19518 32510 19570 32562
rect 19570 32510 19572 32562
rect 19516 32508 19572 32510
rect 17612 32396 17668 32452
rect 20412 33964 20468 34020
rect 20748 33964 20804 34020
rect 20188 32284 20244 32340
rect 20860 32284 20916 32340
rect 20300 31890 20356 31892
rect 20300 31838 20302 31890
rect 20302 31838 20354 31890
rect 20354 31838 20356 31890
rect 20300 31836 20356 31838
rect 19852 31778 19908 31780
rect 19852 31726 19854 31778
rect 19854 31726 19906 31778
rect 19906 31726 19908 31778
rect 19852 31724 19908 31726
rect 16828 30268 16884 30324
rect 17724 30380 17780 30436
rect 16940 30210 16996 30212
rect 16940 30158 16942 30210
rect 16942 30158 16994 30210
rect 16994 30158 16996 30210
rect 16940 30156 16996 30158
rect 15372 28588 15428 28644
rect 16044 28924 16100 28980
rect 15484 28082 15540 28084
rect 15484 28030 15486 28082
rect 15486 28030 15538 28082
rect 15538 28030 15540 28082
rect 15484 28028 15540 28030
rect 15820 27356 15876 27412
rect 16268 27916 16324 27972
rect 16268 26908 16324 26964
rect 17948 29820 18004 29876
rect 18284 30380 18340 30436
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19180 30434 19236 30436
rect 19180 30382 19182 30434
rect 19182 30382 19234 30434
rect 19234 30382 19236 30434
rect 19180 30380 19236 30382
rect 18396 29932 18452 29988
rect 18956 29596 19012 29652
rect 17164 29036 17220 29092
rect 17612 29036 17668 29092
rect 17052 28476 17108 28532
rect 16940 28140 16996 28196
rect 14700 24834 14756 24836
rect 14700 24782 14702 24834
rect 14702 24782 14754 24834
rect 14754 24782 14756 24834
rect 14700 24780 14756 24782
rect 15260 24834 15316 24836
rect 15260 24782 15262 24834
rect 15262 24782 15314 24834
rect 15314 24782 15316 24834
rect 15260 24780 15316 24782
rect 14364 24332 14420 24388
rect 15372 23436 15428 23492
rect 16604 20524 16660 20580
rect 17612 28476 17668 28532
rect 17612 28252 17668 28308
rect 17948 28140 18004 28196
rect 17724 27132 17780 27188
rect 17948 27580 18004 27636
rect 17164 26962 17220 26964
rect 17164 26910 17166 26962
rect 17166 26910 17218 26962
rect 17218 26910 17220 26962
rect 17164 26908 17220 26910
rect 18284 27858 18340 27860
rect 18284 27806 18286 27858
rect 18286 27806 18338 27858
rect 18338 27806 18340 27858
rect 18284 27804 18340 27806
rect 18060 26908 18116 26964
rect 20524 30828 20580 30884
rect 20524 30268 20580 30324
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 21084 29708 21140 29764
rect 19628 29484 19684 29540
rect 19964 29596 20020 29652
rect 20412 29484 20468 29540
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 18844 27858 18900 27860
rect 18844 27806 18846 27858
rect 18846 27806 18898 27858
rect 18898 27806 18900 27858
rect 18844 27804 18900 27806
rect 19180 27580 19236 27636
rect 18508 27186 18564 27188
rect 18508 27134 18510 27186
rect 18510 27134 18562 27186
rect 18562 27134 18564 27186
rect 18508 27132 18564 27134
rect 20300 26908 20356 26964
rect 18172 26012 18228 26068
rect 18172 25676 18228 25732
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19180 26348 19236 26404
rect 18396 26290 18452 26292
rect 18396 26238 18398 26290
rect 18398 26238 18450 26290
rect 18450 26238 18452 26290
rect 18396 26236 18452 26238
rect 18956 26290 19012 26292
rect 18956 26238 18958 26290
rect 18958 26238 19010 26290
rect 19010 26238 19012 26290
rect 18956 26236 19012 26238
rect 18844 24834 18900 24836
rect 18844 24782 18846 24834
rect 18846 24782 18898 24834
rect 18898 24782 18900 24834
rect 18844 24780 18900 24782
rect 18284 24556 18340 24612
rect 17500 23938 17556 23940
rect 17500 23886 17502 23938
rect 17502 23886 17554 23938
rect 17554 23886 17556 23938
rect 17500 23884 17556 23886
rect 16604 18396 16660 18452
rect 15148 17778 15204 17780
rect 15148 17726 15150 17778
rect 15150 17726 15202 17778
rect 15202 17726 15204 17778
rect 15148 17724 15204 17726
rect 16268 17778 16324 17780
rect 16268 17726 16270 17778
rect 16270 17726 16322 17778
rect 16322 17726 16324 17778
rect 16268 17724 16324 17726
rect 14812 16322 14868 16324
rect 14812 16270 14814 16322
rect 14814 16270 14866 16322
rect 14866 16270 14868 16322
rect 14812 16268 14868 16270
rect 14700 15986 14756 15988
rect 14700 15934 14702 15986
rect 14702 15934 14754 15986
rect 14754 15934 14756 15986
rect 14700 15932 14756 15934
rect 14812 15874 14868 15876
rect 14812 15822 14814 15874
rect 14814 15822 14866 15874
rect 14866 15822 14868 15874
rect 14812 15820 14868 15822
rect 14252 14700 14308 14756
rect 14476 14476 14532 14532
rect 13804 14418 13860 14420
rect 13804 14366 13806 14418
rect 13806 14366 13858 14418
rect 13858 14366 13860 14418
rect 13804 14364 13860 14366
rect 13020 14252 13076 14308
rect 13916 13970 13972 13972
rect 13916 13918 13918 13970
rect 13918 13918 13970 13970
rect 13970 13918 13972 13970
rect 13916 13916 13972 13918
rect 14924 14754 14980 14756
rect 14924 14702 14926 14754
rect 14926 14702 14978 14754
rect 14978 14702 14980 14754
rect 14924 14700 14980 14702
rect 14700 14364 14756 14420
rect 14476 13916 14532 13972
rect 14924 14252 14980 14308
rect 14700 13746 14756 13748
rect 14700 13694 14702 13746
rect 14702 13694 14754 13746
rect 14754 13694 14756 13746
rect 14700 13692 14756 13694
rect 15036 13692 15092 13748
rect 14364 13132 14420 13188
rect 15932 17612 15988 17668
rect 15820 16268 15876 16324
rect 15372 13916 15428 13972
rect 15484 13804 15540 13860
rect 15260 13692 15316 13748
rect 15260 13186 15316 13188
rect 15260 13134 15262 13186
rect 15262 13134 15314 13186
rect 15314 13134 15316 13186
rect 15260 13132 15316 13134
rect 15484 12348 15540 12404
rect 16268 17388 16324 17444
rect 16716 17836 16772 17892
rect 16828 17666 16884 17668
rect 16828 17614 16830 17666
rect 16830 17614 16882 17666
rect 16882 17614 16884 17666
rect 16828 17612 16884 17614
rect 16940 17388 16996 17444
rect 16044 16268 16100 16324
rect 16044 16098 16100 16100
rect 16044 16046 16046 16098
rect 16046 16046 16098 16098
rect 16098 16046 16100 16098
rect 16044 16044 16100 16046
rect 16380 15932 16436 15988
rect 16380 15708 16436 15764
rect 16156 15484 16212 15540
rect 16156 14754 16212 14756
rect 16156 14702 16158 14754
rect 16158 14702 16210 14754
rect 16210 14702 16212 14754
rect 16156 14700 16212 14702
rect 15932 14418 15988 14420
rect 15932 14366 15934 14418
rect 15934 14366 15986 14418
rect 15986 14366 15988 14418
rect 15932 14364 15988 14366
rect 16044 14306 16100 14308
rect 16044 14254 16046 14306
rect 16046 14254 16098 14306
rect 16098 14254 16100 14306
rect 16044 14252 16100 14254
rect 16604 14306 16660 14308
rect 16604 14254 16606 14306
rect 16606 14254 16658 14306
rect 16658 14254 16660 14306
rect 16604 14252 16660 14254
rect 17164 16098 17220 16100
rect 17164 16046 17166 16098
rect 17166 16046 17218 16098
rect 17218 16046 17220 16098
rect 17164 16044 17220 16046
rect 17052 15874 17108 15876
rect 17052 15822 17054 15874
rect 17054 15822 17106 15874
rect 17106 15822 17108 15874
rect 17052 15820 17108 15822
rect 16828 15538 16884 15540
rect 16828 15486 16830 15538
rect 16830 15486 16882 15538
rect 16882 15486 16884 15538
rect 16828 15484 16884 15486
rect 17052 14418 17108 14420
rect 17052 14366 17054 14418
rect 17054 14366 17106 14418
rect 17106 14366 17108 14418
rect 17052 14364 17108 14366
rect 16492 13970 16548 13972
rect 16492 13918 16494 13970
rect 16494 13918 16546 13970
rect 16546 13918 16548 13970
rect 16492 13916 16548 13918
rect 15932 13468 15988 13524
rect 16492 13244 16548 13300
rect 15708 12178 15764 12180
rect 15708 12126 15710 12178
rect 15710 12126 15762 12178
rect 15762 12126 15764 12178
rect 15708 12124 15764 12126
rect 14252 12012 14308 12068
rect 10668 10780 10724 10836
rect 14812 10834 14868 10836
rect 14812 10782 14814 10834
rect 14814 10782 14866 10834
rect 14866 10782 14868 10834
rect 14812 10780 14868 10782
rect 15148 11394 15204 11396
rect 15148 11342 15150 11394
rect 15150 11342 15202 11394
rect 15202 11342 15204 11394
rect 15148 11340 15204 11342
rect 15708 11394 15764 11396
rect 15708 11342 15710 11394
rect 15710 11342 15762 11394
rect 15762 11342 15764 11394
rect 15708 11340 15764 11342
rect 15820 10780 15876 10836
rect 15036 10498 15092 10500
rect 15036 10446 15038 10498
rect 15038 10446 15090 10498
rect 15090 10446 15092 10498
rect 15036 10444 15092 10446
rect 14924 9996 14980 10052
rect 14700 9826 14756 9828
rect 14700 9774 14702 9826
rect 14702 9774 14754 9826
rect 14754 9774 14756 9826
rect 14700 9772 14756 9774
rect 16716 13858 16772 13860
rect 16716 13806 16718 13858
rect 16718 13806 16770 13858
rect 16770 13806 16772 13858
rect 16716 13804 16772 13806
rect 16828 13468 16884 13524
rect 18284 23884 18340 23940
rect 17948 23436 18004 23492
rect 19852 26290 19908 26292
rect 19852 26238 19854 26290
rect 19854 26238 19906 26290
rect 19906 26238 19908 26290
rect 19852 26236 19908 26238
rect 19628 26124 19684 26180
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19836 23546 19892 23548
rect 19404 23436 19460 23492
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20412 26290 20468 26292
rect 20412 26238 20414 26290
rect 20414 26238 20466 26290
rect 20466 26238 20468 26290
rect 20412 26236 20468 26238
rect 20524 26908 20580 26964
rect 20412 25282 20468 25284
rect 20412 25230 20414 25282
rect 20414 25230 20466 25282
rect 20466 25230 20468 25282
rect 20412 25228 20468 25230
rect 20860 26178 20916 26180
rect 20860 26126 20862 26178
rect 20862 26126 20914 26178
rect 20914 26126 20916 26178
rect 20860 26124 20916 26126
rect 20972 25730 21028 25732
rect 20972 25678 20974 25730
rect 20974 25678 21026 25730
rect 21026 25678 21028 25730
rect 20972 25676 21028 25678
rect 22316 43484 22372 43540
rect 21644 42140 21700 42196
rect 22764 46956 22820 47012
rect 22764 45388 22820 45444
rect 22764 45218 22820 45220
rect 22764 45166 22766 45218
rect 22766 45166 22818 45218
rect 22818 45166 22820 45218
rect 22764 45164 22820 45166
rect 22540 43372 22596 43428
rect 22428 43148 22484 43204
rect 22652 42924 22708 42980
rect 22652 42700 22708 42756
rect 22204 42530 22260 42532
rect 22204 42478 22206 42530
rect 22206 42478 22258 42530
rect 22258 42478 22260 42530
rect 22204 42476 22260 42478
rect 22540 42476 22596 42532
rect 22428 42140 22484 42196
rect 22652 42028 22708 42084
rect 21868 41468 21924 41524
rect 21644 41074 21700 41076
rect 21644 41022 21646 41074
rect 21646 41022 21698 41074
rect 21698 41022 21700 41074
rect 21644 41020 21700 41022
rect 21980 40908 22036 40964
rect 22204 41410 22260 41412
rect 22204 41358 22206 41410
rect 22206 41358 22258 41410
rect 22258 41358 22260 41410
rect 22204 41356 22260 41358
rect 22540 41020 22596 41076
rect 22204 40908 22260 40964
rect 21868 40348 21924 40404
rect 21644 39452 21700 39508
rect 21756 39788 21812 39844
rect 21644 38780 21700 38836
rect 21644 37938 21700 37940
rect 21644 37886 21646 37938
rect 21646 37886 21698 37938
rect 21698 37886 21700 37938
rect 21644 37884 21700 37886
rect 21420 37378 21476 37380
rect 21420 37326 21422 37378
rect 21422 37326 21474 37378
rect 21474 37326 21476 37378
rect 21420 37324 21476 37326
rect 21644 37378 21700 37380
rect 21644 37326 21646 37378
rect 21646 37326 21698 37378
rect 21698 37326 21700 37378
rect 21644 37324 21700 37326
rect 21868 39618 21924 39620
rect 21868 39566 21870 39618
rect 21870 39566 21922 39618
rect 21922 39566 21924 39618
rect 21868 39564 21924 39566
rect 22092 40402 22148 40404
rect 22092 40350 22094 40402
rect 22094 40350 22146 40402
rect 22146 40350 22148 40402
rect 22092 40348 22148 40350
rect 22092 40124 22148 40180
rect 22652 40348 22708 40404
rect 22428 39788 22484 39844
rect 22204 39676 22260 39732
rect 22540 39618 22596 39620
rect 22540 39566 22542 39618
rect 22542 39566 22594 39618
rect 22594 39566 22596 39618
rect 22540 39564 22596 39566
rect 22316 39452 22372 39508
rect 22652 38722 22708 38724
rect 22652 38670 22654 38722
rect 22654 38670 22706 38722
rect 22706 38670 22708 38722
rect 22652 38668 22708 38670
rect 22204 38108 22260 38164
rect 21980 37212 22036 37268
rect 21868 36652 21924 36708
rect 21644 36204 21700 36260
rect 21868 36092 21924 36148
rect 21644 35922 21700 35924
rect 21644 35870 21646 35922
rect 21646 35870 21698 35922
rect 21698 35870 21700 35922
rect 21644 35868 21700 35870
rect 21532 35810 21588 35812
rect 21532 35758 21534 35810
rect 21534 35758 21586 35810
rect 21586 35758 21588 35810
rect 21532 35756 21588 35758
rect 21868 35196 21924 35252
rect 22092 35308 22148 35364
rect 21644 34412 21700 34468
rect 21868 34130 21924 34132
rect 21868 34078 21870 34130
rect 21870 34078 21922 34130
rect 21922 34078 21924 34130
rect 21868 34076 21924 34078
rect 21532 33964 21588 34020
rect 21644 33234 21700 33236
rect 21644 33182 21646 33234
rect 21646 33182 21698 33234
rect 21698 33182 21700 33234
rect 21644 33180 21700 33182
rect 22092 32786 22148 32788
rect 22092 32734 22094 32786
rect 22094 32734 22146 32786
rect 22146 32734 22148 32786
rect 22092 32732 22148 32734
rect 21980 31890 22036 31892
rect 21980 31838 21982 31890
rect 21982 31838 22034 31890
rect 22034 31838 22036 31890
rect 21980 31836 22036 31838
rect 22540 38332 22596 38388
rect 22540 37660 22596 37716
rect 22652 36988 22708 37044
rect 22652 36258 22708 36260
rect 22652 36206 22654 36258
rect 22654 36206 22706 36258
rect 22706 36206 22708 36258
rect 22652 36204 22708 36206
rect 22652 35196 22708 35252
rect 22428 34130 22484 34132
rect 22428 34078 22430 34130
rect 22430 34078 22482 34130
rect 22482 34078 22484 34130
rect 22428 34076 22484 34078
rect 23212 49420 23268 49476
rect 23772 49868 23828 49924
rect 24108 51324 24164 51380
rect 23996 50876 24052 50932
rect 23884 50482 23940 50484
rect 23884 50430 23886 50482
rect 23886 50430 23938 50482
rect 23938 50430 23940 50482
rect 23884 50428 23940 50430
rect 23100 48860 23156 48916
rect 22988 48412 23044 48468
rect 23212 48802 23268 48804
rect 23212 48750 23214 48802
rect 23214 48750 23266 48802
rect 23266 48750 23268 48802
rect 23212 48748 23268 48750
rect 23436 48860 23492 48916
rect 23548 48636 23604 48692
rect 23212 48242 23268 48244
rect 23212 48190 23214 48242
rect 23214 48190 23266 48242
rect 23266 48190 23268 48242
rect 23212 48188 23268 48190
rect 23436 48300 23492 48356
rect 23324 47628 23380 47684
rect 24444 54626 24500 54628
rect 24444 54574 24446 54626
rect 24446 54574 24498 54626
rect 24498 54574 24500 54626
rect 24444 54572 24500 54574
rect 24556 54460 24612 54516
rect 24556 53506 24612 53508
rect 24556 53454 24558 53506
rect 24558 53454 24610 53506
rect 24610 53454 24612 53506
rect 24556 53452 24612 53454
rect 24780 52834 24836 52836
rect 24780 52782 24782 52834
rect 24782 52782 24834 52834
rect 24834 52782 24836 52834
rect 24780 52780 24836 52782
rect 24556 52108 24612 52164
rect 24668 52050 24724 52052
rect 24668 51998 24670 52050
rect 24670 51998 24722 52050
rect 24722 51998 24724 52050
rect 24668 51996 24724 51998
rect 25004 54460 25060 54516
rect 25452 54012 25508 54068
rect 25452 53842 25508 53844
rect 25452 53790 25454 53842
rect 25454 53790 25506 53842
rect 25506 53790 25508 53842
rect 25452 53788 25508 53790
rect 25004 53618 25060 53620
rect 25004 53566 25006 53618
rect 25006 53566 25058 53618
rect 25058 53566 25060 53618
rect 25004 53564 25060 53566
rect 25340 53004 25396 53060
rect 25228 52386 25284 52388
rect 25228 52334 25230 52386
rect 25230 52334 25282 52386
rect 25282 52334 25284 52386
rect 25228 52332 25284 52334
rect 25004 52108 25060 52164
rect 24892 52050 24948 52052
rect 24892 51998 24894 52050
rect 24894 51998 24946 52050
rect 24946 51998 24948 52050
rect 24892 51996 24948 51998
rect 25340 51772 25396 51828
rect 25676 53676 25732 53732
rect 24780 51490 24836 51492
rect 24780 51438 24782 51490
rect 24782 51438 24834 51490
rect 24834 51438 24836 51490
rect 24780 51436 24836 51438
rect 24332 49922 24388 49924
rect 24332 49870 24334 49922
rect 24334 49870 24386 49922
rect 24386 49870 24388 49922
rect 24332 49868 24388 49870
rect 24108 49138 24164 49140
rect 24108 49086 24110 49138
rect 24110 49086 24162 49138
rect 24162 49086 24164 49138
rect 24108 49084 24164 49086
rect 23660 48354 23716 48356
rect 23660 48302 23662 48354
rect 23662 48302 23714 48354
rect 23714 48302 23716 48354
rect 23660 48300 23716 48302
rect 23436 47458 23492 47460
rect 23436 47406 23438 47458
rect 23438 47406 23490 47458
rect 23490 47406 23492 47458
rect 23436 47404 23492 47406
rect 22988 47292 23044 47348
rect 23548 47852 23604 47908
rect 23212 46844 23268 46900
rect 23100 45836 23156 45892
rect 23436 45890 23492 45892
rect 23436 45838 23438 45890
rect 23438 45838 23490 45890
rect 23490 45838 23492 45890
rect 23436 45836 23492 45838
rect 23212 44322 23268 44324
rect 23212 44270 23214 44322
rect 23214 44270 23266 44322
rect 23266 44270 23268 44322
rect 23212 44268 23268 44270
rect 23436 44268 23492 44324
rect 23100 44044 23156 44100
rect 23324 43820 23380 43876
rect 23100 42700 23156 42756
rect 23100 42476 23156 42532
rect 23324 42194 23380 42196
rect 23324 42142 23326 42194
rect 23326 42142 23378 42194
rect 23378 42142 23380 42194
rect 23324 42140 23380 42142
rect 23100 41692 23156 41748
rect 23212 41580 23268 41636
rect 23324 41804 23380 41860
rect 22876 41356 22932 41412
rect 22988 39618 23044 39620
rect 22988 39566 22990 39618
rect 22990 39566 23042 39618
rect 23042 39566 23044 39618
rect 22988 39564 23044 39566
rect 23660 47740 23716 47796
rect 24556 49810 24612 49812
rect 24556 49758 24558 49810
rect 24558 49758 24610 49810
rect 24610 49758 24612 49810
rect 24556 49756 24612 49758
rect 24556 49308 24612 49364
rect 24668 49084 24724 49140
rect 24780 50988 24836 51044
rect 24668 48748 24724 48804
rect 25340 50652 25396 50708
rect 24892 50482 24948 50484
rect 24892 50430 24894 50482
rect 24894 50430 24946 50482
rect 24946 50430 24948 50482
rect 24892 50428 24948 50430
rect 24892 49922 24948 49924
rect 24892 49870 24894 49922
rect 24894 49870 24946 49922
rect 24946 49870 24948 49922
rect 24892 49868 24948 49870
rect 25116 49196 25172 49252
rect 25564 52050 25620 52052
rect 25564 51998 25566 52050
rect 25566 51998 25618 52050
rect 25618 51998 25620 52050
rect 25564 51996 25620 51998
rect 26236 55186 26292 55188
rect 26236 55134 26238 55186
rect 26238 55134 26290 55186
rect 26290 55134 26292 55186
rect 26236 55132 26292 55134
rect 26124 53058 26180 53060
rect 26124 53006 26126 53058
rect 26126 53006 26178 53058
rect 26178 53006 26180 53058
rect 26124 53004 26180 53006
rect 27468 56306 27524 56308
rect 27468 56254 27470 56306
rect 27470 56254 27522 56306
rect 27522 56254 27524 56306
rect 27468 56252 27524 56254
rect 33852 58156 33908 58212
rect 33628 56700 33684 56756
rect 32956 56588 33012 56644
rect 31276 56364 31332 56420
rect 28924 56252 28980 56308
rect 30268 56252 30324 56308
rect 26572 56194 26628 56196
rect 26572 56142 26574 56194
rect 26574 56142 26626 56194
rect 26626 56142 26628 56194
rect 26572 56140 26628 56142
rect 26572 55468 26628 55524
rect 27916 54908 27972 54964
rect 27132 54796 27188 54852
rect 27244 54684 27300 54740
rect 26684 54572 26740 54628
rect 26908 54626 26964 54628
rect 26908 54574 26910 54626
rect 26910 54574 26962 54626
rect 26962 54574 26964 54626
rect 26908 54572 26964 54574
rect 26796 54514 26852 54516
rect 26796 54462 26798 54514
rect 26798 54462 26850 54514
rect 26850 54462 26852 54514
rect 26796 54460 26852 54462
rect 26684 54402 26740 54404
rect 26684 54350 26686 54402
rect 26686 54350 26738 54402
rect 26738 54350 26740 54402
rect 26684 54348 26740 54350
rect 26572 53788 26628 53844
rect 27020 53788 27076 53844
rect 26460 52780 26516 52836
rect 26572 53618 26628 53620
rect 26572 53566 26574 53618
rect 26574 53566 26626 53618
rect 26626 53566 26628 53618
rect 26572 53564 26628 53566
rect 25900 52444 25956 52500
rect 25676 51548 25732 51604
rect 25564 51490 25620 51492
rect 25564 51438 25566 51490
rect 25566 51438 25618 51490
rect 25618 51438 25620 51490
rect 25564 51436 25620 51438
rect 25788 50316 25844 50372
rect 26460 52444 26516 52500
rect 26124 52050 26180 52052
rect 26124 51998 26126 52050
rect 26126 51998 26178 52050
rect 26178 51998 26180 52050
rect 26124 51996 26180 51998
rect 26796 53170 26852 53172
rect 26796 53118 26798 53170
rect 26798 53118 26850 53170
rect 26850 53118 26852 53170
rect 26796 53116 26852 53118
rect 26684 52946 26740 52948
rect 26684 52894 26686 52946
rect 26686 52894 26738 52946
rect 26738 52894 26740 52946
rect 26684 52892 26740 52894
rect 26684 52332 26740 52388
rect 26796 52780 26852 52836
rect 26572 52108 26628 52164
rect 25900 50204 25956 50260
rect 26124 51772 26180 51828
rect 26236 51548 26292 51604
rect 26124 50092 26180 50148
rect 25564 49532 25620 49588
rect 24780 48636 24836 48692
rect 25340 48972 25396 49028
rect 24108 47852 24164 47908
rect 23996 47740 24052 47796
rect 23772 47292 23828 47348
rect 23660 45388 23716 45444
rect 23884 45836 23940 45892
rect 23548 43596 23604 43652
rect 24108 45388 24164 45444
rect 24892 48130 24948 48132
rect 24892 48078 24894 48130
rect 24894 48078 24946 48130
rect 24946 48078 24948 48130
rect 24892 48076 24948 48078
rect 25228 47964 25284 48020
rect 24444 47458 24500 47460
rect 24444 47406 24446 47458
rect 24446 47406 24498 47458
rect 24498 47406 24500 47458
rect 24444 47404 24500 47406
rect 24892 47404 24948 47460
rect 24332 46674 24388 46676
rect 24332 46622 24334 46674
rect 24334 46622 24386 46674
rect 24386 46622 24388 46674
rect 24332 46620 24388 46622
rect 24780 46396 24836 46452
rect 24108 44322 24164 44324
rect 24108 44270 24110 44322
rect 24110 44270 24162 44322
rect 24162 44270 24164 44322
rect 24108 44268 24164 44270
rect 23996 43932 24052 43988
rect 24220 44156 24276 44212
rect 23660 42700 23716 42756
rect 23548 42588 23604 42644
rect 23772 42028 23828 42084
rect 23660 41804 23716 41860
rect 23772 41186 23828 41188
rect 23772 41134 23774 41186
rect 23774 41134 23826 41186
rect 23826 41134 23828 41186
rect 23772 41132 23828 41134
rect 23548 40796 23604 40852
rect 23436 40684 23492 40740
rect 23548 40402 23604 40404
rect 23548 40350 23550 40402
rect 23550 40350 23602 40402
rect 23602 40350 23604 40402
rect 23548 40348 23604 40350
rect 23660 40236 23716 40292
rect 23100 39394 23156 39396
rect 23100 39342 23102 39394
rect 23102 39342 23154 39394
rect 23154 39342 23156 39394
rect 23100 39340 23156 39342
rect 23660 39788 23716 39844
rect 23212 38946 23268 38948
rect 23212 38894 23214 38946
rect 23214 38894 23266 38946
rect 23266 38894 23268 38946
rect 23212 38892 23268 38894
rect 23212 38668 23268 38724
rect 23660 38332 23716 38388
rect 23436 38162 23492 38164
rect 23436 38110 23438 38162
rect 23438 38110 23490 38162
rect 23490 38110 23492 38162
rect 23436 38108 23492 38110
rect 23324 37772 23380 37828
rect 23660 37996 23716 38052
rect 23324 37324 23380 37380
rect 23212 36988 23268 37044
rect 22764 34860 22820 34916
rect 22540 33964 22596 34020
rect 22428 31724 22484 31780
rect 22540 31836 22596 31892
rect 23772 37436 23828 37492
rect 24108 41468 24164 41524
rect 24108 40796 24164 40852
rect 24444 45106 24500 45108
rect 24444 45054 24446 45106
rect 24446 45054 24498 45106
rect 24498 45054 24500 45106
rect 24444 45052 24500 45054
rect 24780 44882 24836 44884
rect 24780 44830 24782 44882
rect 24782 44830 24834 44882
rect 24834 44830 24836 44882
rect 24780 44828 24836 44830
rect 24556 44716 24612 44772
rect 24556 44098 24612 44100
rect 24556 44046 24558 44098
rect 24558 44046 24610 44098
rect 24610 44046 24612 44098
rect 24556 44044 24612 44046
rect 24444 42530 24500 42532
rect 24444 42478 24446 42530
rect 24446 42478 24498 42530
rect 24498 42478 24500 42530
rect 24444 42476 24500 42478
rect 24668 41970 24724 41972
rect 24668 41918 24670 41970
rect 24670 41918 24722 41970
rect 24722 41918 24724 41970
rect 24668 41916 24724 41918
rect 24556 41580 24612 41636
rect 25004 47068 25060 47124
rect 25116 46956 25172 47012
rect 25116 45948 25172 46004
rect 25452 47570 25508 47572
rect 25452 47518 25454 47570
rect 25454 47518 25506 47570
rect 25506 47518 25508 47570
rect 25452 47516 25508 47518
rect 25452 46844 25508 46900
rect 25452 45612 25508 45668
rect 25340 44604 25396 44660
rect 25004 43426 25060 43428
rect 25004 43374 25006 43426
rect 25006 43374 25058 43426
rect 25058 43374 25060 43426
rect 25004 43372 25060 43374
rect 25004 42028 25060 42084
rect 25004 41580 25060 41636
rect 24556 39900 24612 39956
rect 25228 42028 25284 42084
rect 25228 41298 25284 41300
rect 25228 41246 25230 41298
rect 25230 41246 25282 41298
rect 25282 41246 25284 41298
rect 25228 41244 25284 41246
rect 25228 41020 25284 41076
rect 24780 39452 24836 39508
rect 24668 38722 24724 38724
rect 24668 38670 24670 38722
rect 24670 38670 24722 38722
rect 24722 38670 24724 38722
rect 24668 38668 24724 38670
rect 23996 37660 24052 37716
rect 24220 37548 24276 37604
rect 23660 36370 23716 36372
rect 23660 36318 23662 36370
rect 23662 36318 23714 36370
rect 23714 36318 23716 36370
rect 23660 36316 23716 36318
rect 23548 35420 23604 35476
rect 23212 34412 23268 34468
rect 23436 35308 23492 35364
rect 23100 34242 23156 34244
rect 23100 34190 23102 34242
rect 23102 34190 23154 34242
rect 23154 34190 23156 34242
rect 23100 34188 23156 34190
rect 23996 35196 24052 35252
rect 23884 34802 23940 34804
rect 23884 34750 23886 34802
rect 23886 34750 23938 34802
rect 23938 34750 23940 34802
rect 23884 34748 23940 34750
rect 23996 34188 24052 34244
rect 23884 34076 23940 34132
rect 24220 33964 24276 34020
rect 22764 33234 22820 33236
rect 22764 33182 22766 33234
rect 22766 33182 22818 33234
rect 22818 33182 22820 33234
rect 22764 33180 22820 33182
rect 22988 32844 23044 32900
rect 22652 32508 22708 32564
rect 22876 32732 22932 32788
rect 22876 31500 22932 31556
rect 22316 31164 22372 31220
rect 22540 31276 22596 31332
rect 21980 30770 22036 30772
rect 21980 30718 21982 30770
rect 21982 30718 22034 30770
rect 22034 30718 22036 30770
rect 21980 30716 22036 30718
rect 21420 29484 21476 29540
rect 21532 29708 21588 29764
rect 21196 24668 21252 24724
rect 20636 24610 20692 24612
rect 20636 24558 20638 24610
rect 20638 24558 20690 24610
rect 20690 24558 20692 24610
rect 20636 24556 20692 24558
rect 20300 23436 20356 23492
rect 20972 24332 21028 24388
rect 21980 30322 22036 30324
rect 21980 30270 21982 30322
rect 21982 30270 22034 30322
rect 22034 30270 22036 30322
rect 21980 30268 22036 30270
rect 22428 29986 22484 29988
rect 22428 29934 22430 29986
rect 22430 29934 22482 29986
rect 22482 29934 22484 29986
rect 22428 29932 22484 29934
rect 22316 29820 22372 29876
rect 22316 29148 22372 29204
rect 22428 29708 22484 29764
rect 22428 28754 22484 28756
rect 22428 28702 22430 28754
rect 22430 28702 22482 28754
rect 22482 28702 22484 28754
rect 22428 28700 22484 28702
rect 21868 28364 21924 28420
rect 21644 27580 21700 27636
rect 21980 26962 22036 26964
rect 21980 26910 21982 26962
rect 21982 26910 22034 26962
rect 22034 26910 22036 26962
rect 21980 26908 22036 26910
rect 21532 25282 21588 25284
rect 21532 25230 21534 25282
rect 21534 25230 21586 25282
rect 21586 25230 21588 25282
rect 21532 25228 21588 25230
rect 21756 26124 21812 26180
rect 21420 24946 21476 24948
rect 21420 24894 21422 24946
rect 21422 24894 21474 24946
rect 21474 24894 21476 24946
rect 21420 24892 21476 24894
rect 21868 25676 21924 25732
rect 21308 23996 21364 24052
rect 17836 22204 17892 22260
rect 18732 22258 18788 22260
rect 18732 22206 18734 22258
rect 18734 22206 18786 22258
rect 18786 22206 18788 22258
rect 18732 22204 18788 22206
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20860 19068 20916 19124
rect 18956 18956 19012 19012
rect 18172 18450 18228 18452
rect 18172 18398 18174 18450
rect 18174 18398 18226 18450
rect 18226 18398 18228 18450
rect 18172 18396 18228 18398
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 17500 17890 17556 17892
rect 17500 17838 17502 17890
rect 17502 17838 17554 17890
rect 17554 17838 17556 17890
rect 17500 17836 17556 17838
rect 17836 17612 17892 17668
rect 17612 17442 17668 17444
rect 17612 17390 17614 17442
rect 17614 17390 17666 17442
rect 17666 17390 17668 17442
rect 17612 17388 17668 17390
rect 17836 17052 17892 17108
rect 18620 17554 18676 17556
rect 18620 17502 18622 17554
rect 18622 17502 18674 17554
rect 18674 17502 18676 17554
rect 18620 17500 18676 17502
rect 18508 17442 18564 17444
rect 18508 17390 18510 17442
rect 18510 17390 18562 17442
rect 18562 17390 18564 17442
rect 18508 17388 18564 17390
rect 18396 16828 18452 16884
rect 17612 15484 17668 15540
rect 19852 17778 19908 17780
rect 19852 17726 19854 17778
rect 19854 17726 19906 17778
rect 19906 17726 19908 17778
rect 19852 17724 19908 17726
rect 20524 17778 20580 17780
rect 20524 17726 20526 17778
rect 20526 17726 20578 17778
rect 20578 17726 20580 17778
rect 20524 17724 20580 17726
rect 20300 17666 20356 17668
rect 20300 17614 20302 17666
rect 20302 17614 20354 17666
rect 20354 17614 20356 17666
rect 20300 17612 20356 17614
rect 20188 17500 20244 17556
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 16828 19684 16884
rect 19964 16882 20020 16884
rect 19964 16830 19966 16882
rect 19966 16830 20018 16882
rect 20018 16830 20020 16882
rect 19964 16828 20020 16830
rect 20188 16828 20244 16884
rect 19180 16210 19236 16212
rect 19180 16158 19182 16210
rect 19182 16158 19234 16210
rect 19234 16158 19236 16210
rect 19180 16156 19236 16158
rect 18956 15820 19012 15876
rect 18844 15708 18900 15764
rect 19964 16210 20020 16212
rect 19964 16158 19966 16210
rect 19966 16158 20018 16210
rect 20018 16158 20020 16210
rect 19964 16156 20020 16158
rect 18956 14700 19012 14756
rect 17948 14306 18004 14308
rect 17948 14254 17950 14306
rect 17950 14254 18002 14306
rect 18002 14254 18004 14306
rect 17948 14252 18004 14254
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20412 15708 20468 15764
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 17948 13692 18004 13748
rect 20524 15036 20580 15092
rect 20524 14700 20580 14756
rect 20300 14642 20356 14644
rect 20300 14590 20302 14642
rect 20302 14590 20354 14642
rect 20354 14590 20356 14642
rect 20300 14588 20356 14590
rect 20636 14530 20692 14532
rect 20636 14478 20638 14530
rect 20638 14478 20690 14530
rect 20690 14478 20692 14530
rect 20636 14476 20692 14478
rect 20860 13634 20916 13636
rect 20860 13582 20862 13634
rect 20862 13582 20914 13634
rect 20914 13582 20916 13634
rect 20860 13580 20916 13582
rect 19852 13020 19908 13076
rect 18508 12738 18564 12740
rect 18508 12686 18510 12738
rect 18510 12686 18562 12738
rect 18562 12686 18564 12738
rect 18508 12684 18564 12686
rect 20860 13074 20916 13076
rect 20860 13022 20862 13074
rect 20862 13022 20914 13074
rect 20914 13022 20916 13074
rect 20860 13020 20916 13022
rect 19964 12850 20020 12852
rect 19964 12798 19966 12850
rect 19966 12798 20018 12850
rect 20018 12798 20020 12850
rect 19964 12796 20020 12798
rect 20524 12796 20580 12852
rect 18956 12012 19012 12068
rect 19068 12738 19124 12740
rect 19068 12686 19070 12738
rect 19070 12686 19122 12738
rect 19122 12686 19124 12738
rect 19068 12684 19124 12686
rect 19068 11900 19124 11956
rect 17276 11228 17332 11284
rect 19404 12066 19460 12068
rect 19404 12014 19406 12066
rect 19406 12014 19458 12066
rect 19458 12014 19460 12066
rect 19404 12012 19460 12014
rect 19516 11900 19572 11956
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20524 12572 20580 12628
rect 20044 12516 20100 12518
rect 20300 12066 20356 12068
rect 20300 12014 20302 12066
rect 20302 12014 20354 12066
rect 20354 12014 20356 12066
rect 20300 12012 20356 12014
rect 20524 11900 20580 11956
rect 19292 11340 19348 11396
rect 16268 10668 16324 10724
rect 16156 10444 16212 10500
rect 16044 9884 16100 9940
rect 15596 9772 15652 9828
rect 16492 10556 16548 10612
rect 16828 10722 16884 10724
rect 16828 10670 16830 10722
rect 16830 10670 16882 10722
rect 16882 10670 16884 10722
rect 16828 10668 16884 10670
rect 16940 10610 16996 10612
rect 16940 10558 16942 10610
rect 16942 10558 16994 10610
rect 16994 10558 16996 10610
rect 16940 10556 16996 10558
rect 17724 10610 17780 10612
rect 17724 10558 17726 10610
rect 17726 10558 17778 10610
rect 17778 10558 17780 10610
rect 17724 10556 17780 10558
rect 16716 10444 16772 10500
rect 17612 10444 17668 10500
rect 17500 10050 17556 10052
rect 17500 9998 17502 10050
rect 17502 9998 17554 10050
rect 17554 9998 17556 10050
rect 17500 9996 17556 9998
rect 9212 4508 9268 4564
rect 13020 9154 13076 9156
rect 13020 9102 13022 9154
rect 13022 9102 13074 9154
rect 13074 9102 13076 9154
rect 13020 9100 13076 9102
rect 13804 9100 13860 9156
rect 16492 9660 16548 9716
rect 17836 10050 17892 10052
rect 17836 9998 17838 10050
rect 17838 9998 17890 10050
rect 17890 9998 17892 10050
rect 17836 9996 17892 9998
rect 17276 8258 17332 8260
rect 17276 8206 17278 8258
rect 17278 8206 17330 8258
rect 17330 8206 17332 8258
rect 17276 8204 17332 8206
rect 18060 10722 18116 10724
rect 18060 10670 18062 10722
rect 18062 10670 18114 10722
rect 18114 10670 18116 10722
rect 18060 10668 18116 10670
rect 18284 10444 18340 10500
rect 18620 9996 18676 10052
rect 18284 9884 18340 9940
rect 18508 8258 18564 8260
rect 18508 8206 18510 8258
rect 18510 8206 18562 8258
rect 18562 8206 18564 8258
rect 18508 8204 18564 8206
rect 19740 11394 19796 11396
rect 19740 11342 19742 11394
rect 19742 11342 19794 11394
rect 19794 11342 19796 11394
rect 19740 11340 19796 11342
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19292 10498 19348 10500
rect 19292 10446 19294 10498
rect 19294 10446 19346 10498
rect 19346 10446 19348 10498
rect 19292 10444 19348 10446
rect 19068 9996 19124 10052
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 20300 8988 20356 9044
rect 19740 8316 19796 8372
rect 19180 8204 19236 8260
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 20412 8370 20468 8372
rect 20412 8318 20414 8370
rect 20414 8318 20466 8370
rect 20466 8318 20468 8370
rect 20412 8316 20468 8318
rect 20636 8258 20692 8260
rect 20636 8206 20638 8258
rect 20638 8206 20690 8258
rect 20690 8206 20692 8258
rect 20636 8204 20692 8206
rect 19404 6972 19460 7028
rect 19292 6690 19348 6692
rect 19292 6638 19294 6690
rect 19294 6638 19346 6690
rect 19346 6638 19348 6690
rect 19292 6636 19348 6638
rect 18844 5068 18900 5124
rect 20748 7474 20804 7476
rect 20748 7422 20750 7474
rect 20750 7422 20802 7474
rect 20802 7422 20804 7474
rect 20748 7420 20804 7422
rect 22652 31218 22708 31220
rect 22652 31166 22654 31218
rect 22654 31166 22706 31218
rect 22706 31166 22708 31218
rect 22652 31164 22708 31166
rect 22764 30268 22820 30324
rect 22652 29932 22708 29988
rect 22876 29986 22932 29988
rect 22876 29934 22878 29986
rect 22878 29934 22930 29986
rect 22930 29934 22932 29986
rect 22876 29932 22932 29934
rect 23548 33122 23604 33124
rect 23548 33070 23550 33122
rect 23550 33070 23602 33122
rect 23602 33070 23604 33122
rect 23548 33068 23604 33070
rect 24108 33122 24164 33124
rect 24108 33070 24110 33122
rect 24110 33070 24162 33122
rect 24162 33070 24164 33122
rect 24108 33068 24164 33070
rect 23660 31778 23716 31780
rect 23660 31726 23662 31778
rect 23662 31726 23714 31778
rect 23714 31726 23716 31778
rect 23660 31724 23716 31726
rect 24444 38050 24500 38052
rect 24444 37998 24446 38050
rect 24446 37998 24498 38050
rect 24498 37998 24500 38050
rect 24444 37996 24500 37998
rect 24892 37826 24948 37828
rect 24892 37774 24894 37826
rect 24894 37774 24946 37826
rect 24946 37774 24948 37826
rect 24892 37772 24948 37774
rect 24556 36370 24612 36372
rect 24556 36318 24558 36370
rect 24558 36318 24610 36370
rect 24610 36318 24612 36370
rect 24556 36316 24612 36318
rect 24668 35420 24724 35476
rect 24780 35196 24836 35252
rect 24668 34914 24724 34916
rect 24668 34862 24670 34914
rect 24670 34862 24722 34914
rect 24722 34862 24724 34914
rect 24668 34860 24724 34862
rect 24556 34748 24612 34804
rect 24444 34412 24500 34468
rect 24556 34188 24612 34244
rect 24668 34300 24724 34356
rect 24108 31554 24164 31556
rect 24108 31502 24110 31554
rect 24110 31502 24162 31554
rect 24162 31502 24164 31554
rect 24108 31500 24164 31502
rect 23772 31218 23828 31220
rect 23772 31166 23774 31218
rect 23774 31166 23826 31218
rect 23826 31166 23828 31218
rect 23772 31164 23828 31166
rect 23324 29932 23380 29988
rect 24220 29820 24276 29876
rect 23324 29148 23380 29204
rect 23996 29148 24052 29204
rect 23548 28924 23604 28980
rect 23996 28700 24052 28756
rect 25004 35420 25060 35476
rect 25452 42140 25508 42196
rect 25452 41916 25508 41972
rect 25340 39004 25396 39060
rect 25452 40684 25508 40740
rect 25676 45948 25732 46004
rect 26124 48748 26180 48804
rect 26236 50316 26292 50372
rect 26012 48412 26068 48468
rect 26012 47964 26068 48020
rect 26012 47346 26068 47348
rect 26012 47294 26014 47346
rect 26014 47294 26066 47346
rect 26066 47294 26068 47346
rect 26012 47292 26068 47294
rect 26124 47180 26180 47236
rect 26796 51548 26852 51604
rect 27020 52780 27076 52836
rect 27132 52444 27188 52500
rect 27692 54626 27748 54628
rect 27692 54574 27694 54626
rect 27694 54574 27746 54626
rect 27746 54574 27748 54626
rect 27692 54572 27748 54574
rect 27356 53618 27412 53620
rect 27356 53566 27358 53618
rect 27358 53566 27410 53618
rect 27410 53566 27412 53618
rect 27356 53564 27412 53566
rect 28252 55298 28308 55300
rect 28252 55246 28254 55298
rect 28254 55246 28306 55298
rect 28306 55246 28308 55298
rect 28252 55244 28308 55246
rect 28028 53842 28084 53844
rect 28028 53790 28030 53842
rect 28030 53790 28082 53842
rect 28082 53790 28084 53842
rect 28028 53788 28084 53790
rect 29260 55970 29316 55972
rect 29260 55918 29262 55970
rect 29262 55918 29314 55970
rect 29314 55918 29316 55970
rect 29260 55916 29316 55918
rect 28476 55410 28532 55412
rect 28476 55358 28478 55410
rect 28478 55358 28530 55410
rect 28530 55358 28532 55410
rect 28476 55356 28532 55358
rect 32172 55970 32228 55972
rect 32172 55918 32174 55970
rect 32174 55918 32226 55970
rect 32226 55918 32228 55970
rect 32172 55916 32228 55918
rect 29932 55298 29988 55300
rect 29932 55246 29934 55298
rect 29934 55246 29986 55298
rect 29986 55246 29988 55298
rect 29932 55244 29988 55246
rect 30156 55186 30212 55188
rect 30156 55134 30158 55186
rect 30158 55134 30210 55186
rect 30210 55134 30212 55186
rect 30156 55132 30212 55134
rect 28476 55020 28532 55076
rect 28588 54908 28644 54964
rect 28364 53676 28420 53732
rect 27916 53228 27972 53284
rect 27916 53058 27972 53060
rect 27916 53006 27918 53058
rect 27918 53006 27970 53058
rect 27970 53006 27972 53058
rect 27916 53004 27972 53006
rect 27804 52946 27860 52948
rect 27804 52894 27806 52946
rect 27806 52894 27858 52946
rect 27858 52894 27860 52946
rect 27804 52892 27860 52894
rect 27468 52444 27524 52500
rect 27020 51772 27076 51828
rect 27132 51996 27188 52052
rect 27244 51772 27300 51828
rect 27132 51324 27188 51380
rect 27692 52108 27748 52164
rect 27580 50652 27636 50708
rect 27356 50540 27412 50596
rect 27020 50428 27076 50484
rect 26460 49868 26516 49924
rect 26348 48802 26404 48804
rect 26348 48750 26350 48802
rect 26350 48750 26402 48802
rect 26402 48750 26404 48802
rect 26348 48748 26404 48750
rect 26236 45612 26292 45668
rect 26348 48188 26404 48244
rect 26012 45164 26068 45220
rect 26124 45106 26180 45108
rect 26124 45054 26126 45106
rect 26126 45054 26178 45106
rect 26178 45054 26180 45106
rect 26124 45052 26180 45054
rect 25900 44604 25956 44660
rect 25900 44434 25956 44436
rect 25900 44382 25902 44434
rect 25902 44382 25954 44434
rect 25954 44382 25956 44434
rect 25900 44380 25956 44382
rect 28476 52834 28532 52836
rect 28476 52782 28478 52834
rect 28478 52782 28530 52834
rect 28530 52782 28532 52834
rect 28476 52780 28532 52782
rect 28140 51436 28196 51492
rect 27804 50482 27860 50484
rect 27804 50430 27806 50482
rect 27806 50430 27858 50482
rect 27858 50430 27860 50482
rect 27804 50428 27860 50430
rect 26684 48076 26740 48132
rect 26572 47964 26628 48020
rect 26572 47516 26628 47572
rect 26460 44604 26516 44660
rect 26460 44156 26516 44212
rect 25900 43426 25956 43428
rect 25900 43374 25902 43426
rect 25902 43374 25954 43426
rect 25954 43374 25956 43426
rect 25900 43372 25956 43374
rect 26348 43372 26404 43428
rect 26012 42866 26068 42868
rect 26012 42814 26014 42866
rect 26014 42814 26066 42866
rect 26066 42814 26068 42866
rect 26012 42812 26068 42814
rect 25676 42700 25732 42756
rect 25676 41970 25732 41972
rect 25676 41918 25678 41970
rect 25678 41918 25730 41970
rect 25730 41918 25732 41970
rect 25676 41916 25732 41918
rect 25788 41244 25844 41300
rect 26460 42140 26516 42196
rect 26012 42082 26068 42084
rect 26012 42030 26014 42082
rect 26014 42030 26066 42082
rect 26066 42030 26068 42082
rect 26012 42028 26068 42030
rect 26908 48076 26964 48132
rect 27804 49922 27860 49924
rect 27804 49870 27806 49922
rect 27806 49870 27858 49922
rect 27858 49870 27860 49922
rect 27804 49868 27860 49870
rect 28700 54348 28756 54404
rect 29148 54348 29204 54404
rect 28700 53900 28756 53956
rect 28924 53954 28980 53956
rect 28924 53902 28926 53954
rect 28926 53902 28978 53954
rect 28978 53902 28980 53954
rect 28924 53900 28980 53902
rect 30044 55074 30100 55076
rect 30044 55022 30046 55074
rect 30046 55022 30098 55074
rect 30098 55022 30100 55074
rect 30044 55020 30100 55022
rect 29708 54908 29764 54964
rect 29932 54402 29988 54404
rect 29932 54350 29934 54402
rect 29934 54350 29986 54402
rect 29986 54350 29988 54402
rect 29932 54348 29988 54350
rect 30156 53730 30212 53732
rect 30156 53678 30158 53730
rect 30158 53678 30210 53730
rect 30210 53678 30212 53730
rect 30156 53676 30212 53678
rect 29372 52834 29428 52836
rect 29372 52782 29374 52834
rect 29374 52782 29426 52834
rect 29426 52782 29428 52834
rect 29372 52780 29428 52782
rect 28924 52556 28980 52612
rect 28364 51378 28420 51380
rect 28364 51326 28366 51378
rect 28366 51326 28418 51378
rect 28418 51326 28420 51378
rect 28364 51324 28420 51326
rect 28812 50652 28868 50708
rect 28476 50482 28532 50484
rect 28476 50430 28478 50482
rect 28478 50430 28530 50482
rect 28530 50430 28532 50482
rect 28476 50428 28532 50430
rect 28252 49980 28308 50036
rect 28364 50316 28420 50372
rect 28364 49756 28420 49812
rect 28252 49420 28308 49476
rect 28924 49420 28980 49476
rect 28252 49138 28308 49140
rect 28252 49086 28254 49138
rect 28254 49086 28306 49138
rect 28306 49086 28308 49138
rect 28252 49084 28308 49086
rect 28924 48972 28980 49028
rect 29036 49084 29092 49140
rect 27468 48860 27524 48916
rect 27132 48188 27188 48244
rect 26684 45276 26740 45332
rect 26684 44380 26740 44436
rect 26684 44210 26740 44212
rect 26684 44158 26686 44210
rect 26686 44158 26738 44210
rect 26738 44158 26740 44210
rect 26684 44156 26740 44158
rect 26684 43596 26740 43652
rect 27244 47404 27300 47460
rect 27356 46732 27412 46788
rect 27020 46396 27076 46452
rect 27244 46284 27300 46340
rect 27020 45666 27076 45668
rect 27020 45614 27022 45666
rect 27022 45614 27074 45666
rect 27074 45614 27076 45666
rect 27020 45612 27076 45614
rect 26908 44994 26964 44996
rect 26908 44942 26910 44994
rect 26910 44942 26962 44994
rect 26962 44942 26964 44994
rect 26908 44940 26964 44942
rect 27132 45106 27188 45108
rect 27132 45054 27134 45106
rect 27134 45054 27186 45106
rect 27186 45054 27188 45106
rect 27132 45052 27188 45054
rect 27132 44604 27188 44660
rect 27356 45218 27412 45220
rect 27356 45166 27358 45218
rect 27358 45166 27410 45218
rect 27410 45166 27412 45218
rect 27356 45164 27412 45166
rect 27020 43596 27076 43652
rect 26796 42252 26852 42308
rect 27020 43260 27076 43316
rect 26684 42082 26740 42084
rect 26684 42030 26686 42082
rect 26686 42030 26738 42082
rect 26738 42030 26740 42082
rect 26684 42028 26740 42030
rect 26908 42082 26964 42084
rect 26908 42030 26910 42082
rect 26910 42030 26962 42082
rect 26962 42030 26964 42082
rect 26908 42028 26964 42030
rect 27020 41916 27076 41972
rect 26348 41298 26404 41300
rect 26348 41246 26350 41298
rect 26350 41246 26402 41298
rect 26402 41246 26404 41298
rect 26348 41244 26404 41246
rect 27020 41356 27076 41412
rect 25788 41074 25844 41076
rect 25788 41022 25790 41074
rect 25790 41022 25842 41074
rect 25842 41022 25844 41074
rect 25788 41020 25844 41022
rect 26124 40684 26180 40740
rect 25900 40572 25956 40628
rect 25900 39452 25956 39508
rect 25676 39004 25732 39060
rect 25564 38668 25620 38724
rect 25788 38834 25844 38836
rect 25788 38782 25790 38834
rect 25790 38782 25842 38834
rect 25842 38782 25844 38834
rect 25788 38780 25844 38782
rect 26348 40626 26404 40628
rect 26348 40574 26350 40626
rect 26350 40574 26402 40626
rect 26402 40574 26404 40626
rect 26348 40572 26404 40574
rect 26012 38892 26068 38948
rect 26460 38780 26516 38836
rect 26012 38332 26068 38388
rect 25788 37826 25844 37828
rect 25788 37774 25790 37826
rect 25790 37774 25842 37826
rect 25842 37774 25844 37826
rect 25788 37772 25844 37774
rect 25676 36540 25732 36596
rect 25452 36258 25508 36260
rect 25452 36206 25454 36258
rect 25454 36206 25506 36258
rect 25506 36206 25508 36258
rect 25452 36204 25508 36206
rect 25564 35420 25620 35476
rect 25228 34300 25284 34356
rect 24892 33068 24948 33124
rect 26012 34972 26068 35028
rect 25564 34354 25620 34356
rect 25564 34302 25566 34354
rect 25566 34302 25618 34354
rect 25618 34302 25620 34354
rect 25564 34300 25620 34302
rect 26012 33740 26068 33796
rect 24556 30716 24612 30772
rect 25004 32284 25060 32340
rect 24332 28700 24388 28756
rect 24892 29932 24948 29988
rect 24780 27634 24836 27636
rect 24780 27582 24782 27634
rect 24782 27582 24834 27634
rect 24834 27582 24836 27634
rect 24780 27580 24836 27582
rect 22540 24892 22596 24948
rect 23772 26908 23828 26964
rect 22540 24220 22596 24276
rect 21980 23714 22036 23716
rect 21980 23662 21982 23714
rect 21982 23662 22034 23714
rect 22034 23662 22036 23714
rect 21980 23660 22036 23662
rect 21756 23548 21812 23604
rect 21308 23436 21364 23492
rect 21756 21474 21812 21476
rect 21756 21422 21758 21474
rect 21758 21422 21810 21474
rect 21810 21422 21812 21474
rect 21756 21420 21812 21422
rect 21644 19122 21700 19124
rect 21644 19070 21646 19122
rect 21646 19070 21698 19122
rect 21698 19070 21700 19122
rect 21644 19068 21700 19070
rect 21308 18844 21364 18900
rect 21196 18450 21252 18452
rect 21196 18398 21198 18450
rect 21198 18398 21250 18450
rect 21250 18398 21252 18450
rect 21196 18396 21252 18398
rect 21420 17612 21476 17668
rect 21308 16882 21364 16884
rect 21308 16830 21310 16882
rect 21310 16830 21362 16882
rect 21362 16830 21364 16882
rect 21308 16828 21364 16830
rect 22764 24220 22820 24276
rect 22652 21644 22708 21700
rect 22428 21586 22484 21588
rect 22428 21534 22430 21586
rect 22430 21534 22482 21586
rect 22482 21534 22484 21586
rect 22428 21532 22484 21534
rect 22316 21420 22372 21476
rect 22204 19852 22260 19908
rect 22092 19010 22148 19012
rect 22092 18958 22094 19010
rect 22094 18958 22146 19010
rect 22146 18958 22148 19010
rect 22092 18956 22148 18958
rect 22204 18396 22260 18452
rect 22092 17388 22148 17444
rect 21868 16828 21924 16884
rect 21532 16210 21588 16212
rect 21532 16158 21534 16210
rect 21534 16158 21586 16210
rect 21586 16158 21588 16210
rect 21532 16156 21588 16158
rect 21532 14588 21588 14644
rect 21980 15708 22036 15764
rect 21980 13580 22036 13636
rect 21196 13020 21252 13076
rect 21196 12572 21252 12628
rect 21868 12572 21924 12628
rect 21980 12178 22036 12180
rect 21980 12126 21982 12178
rect 21982 12126 22034 12178
rect 22034 12126 22036 12178
rect 21980 12124 22036 12126
rect 21084 9884 21140 9940
rect 21532 9938 21588 9940
rect 21532 9886 21534 9938
rect 21534 9886 21586 9938
rect 21586 9886 21588 9938
rect 21532 9884 21588 9886
rect 21756 9884 21812 9940
rect 21084 9042 21140 9044
rect 21084 8990 21086 9042
rect 21086 8990 21138 9042
rect 21138 8990 21140 9042
rect 21084 8988 21140 8990
rect 21644 7420 21700 7476
rect 20972 6972 21028 7028
rect 20412 6636 20468 6692
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19628 6076 19684 6132
rect 20636 6130 20692 6132
rect 20636 6078 20638 6130
rect 20638 6078 20690 6130
rect 20690 6078 20692 6130
rect 20636 6076 20692 6078
rect 22540 21420 22596 21476
rect 23212 24220 23268 24276
rect 22988 23826 23044 23828
rect 22988 23774 22990 23826
rect 22990 23774 23042 23826
rect 23042 23774 23044 23826
rect 22988 23772 23044 23774
rect 23100 23660 23156 23716
rect 24556 26962 24612 26964
rect 24556 26910 24558 26962
rect 24558 26910 24610 26962
rect 24610 26910 24612 26962
rect 24556 26908 24612 26910
rect 24444 26796 24500 26852
rect 25116 28028 25172 28084
rect 24892 26850 24948 26852
rect 24892 26798 24894 26850
rect 24894 26798 24946 26850
rect 24946 26798 24948 26850
rect 24892 26796 24948 26798
rect 25004 26572 25060 26628
rect 24108 25116 24164 25172
rect 24668 25116 24724 25172
rect 24668 24834 24724 24836
rect 24668 24782 24670 24834
rect 24670 24782 24722 24834
rect 24722 24782 24724 24834
rect 24668 24780 24724 24782
rect 24892 24556 24948 24612
rect 24332 24050 24388 24052
rect 24332 23998 24334 24050
rect 24334 23998 24386 24050
rect 24386 23998 24388 24050
rect 24332 23996 24388 23998
rect 24108 23660 24164 23716
rect 24668 23548 24724 23604
rect 23212 22428 23268 22484
rect 23772 22482 23828 22484
rect 23772 22430 23774 22482
rect 23774 22430 23826 22482
rect 23826 22430 23828 22482
rect 23772 22428 23828 22430
rect 25116 24332 25172 24388
rect 25676 32508 25732 32564
rect 26012 32674 26068 32676
rect 26012 32622 26014 32674
rect 26014 32622 26066 32674
rect 26066 32622 26068 32674
rect 26012 32620 26068 32622
rect 25900 31836 25956 31892
rect 27244 43650 27300 43652
rect 27244 43598 27246 43650
rect 27246 43598 27298 43650
rect 27298 43598 27300 43650
rect 27244 43596 27300 43598
rect 27916 47964 27972 48020
rect 28588 47852 28644 47908
rect 28476 47740 28532 47796
rect 28140 47458 28196 47460
rect 28140 47406 28142 47458
rect 28142 47406 28194 47458
rect 28194 47406 28196 47458
rect 28140 47404 28196 47406
rect 27580 47068 27636 47124
rect 28140 46956 28196 47012
rect 28028 46786 28084 46788
rect 28028 46734 28030 46786
rect 28030 46734 28082 46786
rect 28082 46734 28084 46786
rect 28028 46732 28084 46734
rect 28364 46450 28420 46452
rect 28364 46398 28366 46450
rect 28366 46398 28418 46450
rect 28418 46398 28420 46450
rect 28364 46396 28420 46398
rect 28252 45500 28308 45556
rect 28140 45276 28196 45332
rect 28028 45218 28084 45220
rect 28028 45166 28030 45218
rect 28030 45166 28082 45218
rect 28082 45166 28084 45218
rect 28028 45164 28084 45166
rect 28140 45106 28196 45108
rect 28140 45054 28142 45106
rect 28142 45054 28194 45106
rect 28194 45054 28196 45106
rect 28140 45052 28196 45054
rect 27692 44604 27748 44660
rect 27692 43932 27748 43988
rect 28252 43932 28308 43988
rect 26796 40626 26852 40628
rect 26796 40574 26798 40626
rect 26798 40574 26850 40626
rect 26850 40574 26852 40626
rect 26796 40572 26852 40574
rect 26684 38892 26740 38948
rect 26572 38332 26628 38388
rect 26684 38274 26740 38276
rect 26684 38222 26686 38274
rect 26686 38222 26738 38274
rect 26738 38222 26740 38274
rect 26684 38220 26740 38222
rect 26572 38050 26628 38052
rect 26572 37998 26574 38050
rect 26574 37998 26626 38050
rect 26626 37998 26628 38050
rect 26572 37996 26628 37998
rect 26236 37266 26292 37268
rect 26236 37214 26238 37266
rect 26238 37214 26290 37266
rect 26290 37214 26292 37266
rect 26236 37212 26292 37214
rect 26684 37772 26740 37828
rect 26684 37100 26740 37156
rect 26460 36988 26516 37044
rect 26236 36876 26292 36932
rect 26236 36594 26292 36596
rect 26236 36542 26238 36594
rect 26238 36542 26290 36594
rect 26290 36542 26292 36594
rect 26236 36540 26292 36542
rect 26908 36876 26964 36932
rect 26348 35196 26404 35252
rect 27580 42194 27636 42196
rect 27580 42142 27582 42194
rect 27582 42142 27634 42194
rect 27634 42142 27636 42194
rect 27580 42140 27636 42142
rect 28028 42364 28084 42420
rect 27916 41916 27972 41972
rect 26908 35026 26964 35028
rect 26908 34974 26910 35026
rect 26910 34974 26962 35026
rect 26962 34974 26964 35026
rect 26908 34972 26964 34974
rect 26572 33740 26628 33796
rect 26908 34076 26964 34132
rect 27356 40684 27412 40740
rect 27356 38834 27412 38836
rect 27356 38782 27358 38834
rect 27358 38782 27410 38834
rect 27410 38782 27412 38834
rect 27356 38780 27412 38782
rect 27244 38220 27300 38276
rect 27356 38050 27412 38052
rect 27356 37998 27358 38050
rect 27358 37998 27410 38050
rect 27410 37998 27412 38050
rect 27356 37996 27412 37998
rect 27692 39452 27748 39508
rect 27580 38892 27636 38948
rect 27916 41244 27972 41300
rect 28028 40626 28084 40628
rect 28028 40574 28030 40626
rect 28030 40574 28082 40626
rect 28082 40574 28084 40626
rect 28028 40572 28084 40574
rect 28700 43820 28756 43876
rect 30604 55410 30660 55412
rect 30604 55358 30606 55410
rect 30606 55358 30658 55410
rect 30658 55358 30660 55410
rect 30604 55356 30660 55358
rect 32172 55356 32228 55412
rect 33628 56306 33684 56308
rect 33628 56254 33630 56306
rect 33630 56254 33682 56306
rect 33682 56254 33684 56306
rect 33628 56252 33684 56254
rect 33068 55468 33124 55524
rect 33292 55916 33348 55972
rect 30604 55132 30660 55188
rect 31164 55186 31220 55188
rect 31164 55134 31166 55186
rect 31166 55134 31218 55186
rect 31218 55134 31220 55186
rect 31164 55132 31220 55134
rect 30716 55020 30772 55076
rect 31388 55074 31444 55076
rect 31388 55022 31390 55074
rect 31390 55022 31442 55074
rect 31442 55022 31444 55074
rect 31388 55020 31444 55022
rect 31164 54908 31220 54964
rect 30940 54738 30996 54740
rect 30940 54686 30942 54738
rect 30942 54686 30994 54738
rect 30994 54686 30996 54738
rect 30940 54684 30996 54686
rect 30492 54236 30548 54292
rect 31612 54908 31668 54964
rect 30604 53900 30660 53956
rect 30940 54348 30996 54404
rect 30380 53788 30436 53844
rect 30828 53842 30884 53844
rect 30828 53790 30830 53842
rect 30830 53790 30882 53842
rect 30882 53790 30884 53842
rect 30828 53788 30884 53790
rect 30268 52668 30324 52724
rect 30828 53340 30884 53396
rect 30716 52332 30772 52388
rect 29820 52274 29876 52276
rect 29820 52222 29822 52274
rect 29822 52222 29874 52274
rect 29874 52222 29876 52274
rect 29820 52220 29876 52222
rect 29708 51436 29764 51492
rect 29148 44716 29204 44772
rect 28924 43708 28980 43764
rect 28252 41804 28308 41860
rect 28252 40572 28308 40628
rect 28364 41580 28420 41636
rect 28588 41970 28644 41972
rect 28588 41918 28590 41970
rect 28590 41918 28642 41970
rect 28642 41918 28644 41970
rect 28588 41916 28644 41918
rect 28924 41132 28980 41188
rect 28476 41020 28532 41076
rect 28924 40460 28980 40516
rect 28364 39004 28420 39060
rect 28700 38946 28756 38948
rect 28700 38894 28702 38946
rect 28702 38894 28754 38946
rect 28754 38894 28756 38946
rect 28700 38892 28756 38894
rect 28140 38668 28196 38724
rect 28476 38834 28532 38836
rect 28476 38782 28478 38834
rect 28478 38782 28530 38834
rect 28530 38782 28532 38834
rect 28476 38780 28532 38782
rect 28812 38668 28868 38724
rect 28364 38220 28420 38276
rect 28812 38444 28868 38500
rect 28252 37548 28308 37604
rect 27468 37100 27524 37156
rect 27132 33628 27188 33684
rect 27244 36988 27300 37044
rect 26460 32508 26516 32564
rect 26236 29986 26292 29988
rect 26236 29934 26238 29986
rect 26238 29934 26290 29986
rect 26290 29934 26292 29986
rect 26236 29932 26292 29934
rect 25564 29484 25620 29540
rect 25900 28754 25956 28756
rect 25900 28702 25902 28754
rect 25902 28702 25954 28754
rect 25954 28702 25956 28754
rect 25900 28700 25956 28702
rect 25676 28082 25732 28084
rect 25676 28030 25678 28082
rect 25678 28030 25730 28082
rect 25730 28030 25732 28082
rect 25676 28028 25732 28030
rect 27020 31612 27076 31668
rect 28140 37266 28196 37268
rect 28140 37214 28142 37266
rect 28142 37214 28194 37266
rect 28194 37214 28196 37266
rect 28140 37212 28196 37214
rect 27916 36988 27972 37044
rect 27692 36706 27748 36708
rect 27692 36654 27694 36706
rect 27694 36654 27746 36706
rect 27746 36654 27748 36706
rect 27692 36652 27748 36654
rect 28476 37100 28532 37156
rect 28700 36764 28756 36820
rect 28812 36428 28868 36484
rect 29148 37154 29204 37156
rect 29148 37102 29150 37154
rect 29150 37102 29202 37154
rect 29202 37102 29204 37154
rect 29148 37100 29204 37102
rect 29372 50316 29428 50372
rect 29372 48972 29428 49028
rect 30380 51490 30436 51492
rect 30380 51438 30382 51490
rect 30382 51438 30434 51490
rect 30434 51438 30436 51490
rect 30380 51436 30436 51438
rect 29820 51212 29876 51268
rect 29932 50706 29988 50708
rect 29932 50654 29934 50706
rect 29934 50654 29986 50706
rect 29986 50654 29988 50706
rect 29932 50652 29988 50654
rect 29932 48412 29988 48468
rect 29932 48242 29988 48244
rect 29932 48190 29934 48242
rect 29934 48190 29986 48242
rect 29986 48190 29988 48242
rect 29932 48188 29988 48190
rect 29484 47180 29540 47236
rect 30156 51212 30212 51268
rect 31612 54684 31668 54740
rect 32172 54908 32228 54964
rect 32620 54908 32676 54964
rect 31276 54402 31332 54404
rect 31276 54350 31278 54402
rect 31278 54350 31330 54402
rect 31330 54350 31332 54402
rect 31276 54348 31332 54350
rect 31164 53788 31220 53844
rect 31948 53676 32004 53732
rect 31948 53116 32004 53172
rect 31276 51996 31332 52052
rect 31276 51660 31332 51716
rect 31052 51602 31108 51604
rect 31052 51550 31054 51602
rect 31054 51550 31106 51602
rect 31106 51550 31108 51602
rect 31052 51548 31108 51550
rect 32060 52220 32116 52276
rect 31836 52050 31892 52052
rect 31836 51998 31838 52050
rect 31838 51998 31890 52050
rect 31890 51998 31892 52050
rect 31836 51996 31892 51998
rect 31612 51548 31668 51604
rect 31612 51378 31668 51380
rect 31612 51326 31614 51378
rect 31614 51326 31666 51378
rect 31666 51326 31668 51378
rect 31612 51324 31668 51326
rect 31388 51100 31444 51156
rect 30156 50092 30212 50148
rect 30604 50428 30660 50484
rect 30828 49868 30884 49924
rect 29820 47516 29876 47572
rect 30604 49026 30660 49028
rect 30604 48974 30606 49026
rect 30606 48974 30658 49026
rect 30658 48974 30660 49026
rect 30604 48972 30660 48974
rect 30156 47628 30212 47684
rect 30268 47570 30324 47572
rect 30268 47518 30270 47570
rect 30270 47518 30322 47570
rect 30322 47518 30324 47570
rect 30268 47516 30324 47518
rect 30156 47180 30212 47236
rect 29484 46172 29540 46228
rect 29484 45500 29540 45556
rect 30044 45500 30100 45556
rect 29372 44044 29428 44100
rect 29372 43708 29428 43764
rect 29484 42924 29540 42980
rect 29708 44098 29764 44100
rect 29708 44046 29710 44098
rect 29710 44046 29762 44098
rect 29762 44046 29764 44098
rect 29708 44044 29764 44046
rect 29708 43820 29764 43876
rect 30156 43708 30212 43764
rect 29932 42924 29988 42980
rect 29596 42364 29652 42420
rect 29484 42140 29540 42196
rect 30156 42588 30212 42644
rect 29820 42028 29876 42084
rect 29372 40908 29428 40964
rect 29372 40514 29428 40516
rect 29372 40462 29374 40514
rect 29374 40462 29426 40514
rect 29426 40462 29428 40514
rect 29372 40460 29428 40462
rect 29596 40962 29652 40964
rect 29596 40910 29598 40962
rect 29598 40910 29650 40962
rect 29650 40910 29652 40962
rect 29596 40908 29652 40910
rect 30044 40962 30100 40964
rect 30044 40910 30046 40962
rect 30046 40910 30098 40962
rect 30098 40910 30100 40962
rect 30044 40908 30100 40910
rect 29484 38108 29540 38164
rect 30044 39058 30100 39060
rect 30044 39006 30046 39058
rect 30046 39006 30098 39058
rect 30098 39006 30100 39058
rect 30044 39004 30100 39006
rect 29820 38444 29876 38500
rect 29596 38050 29652 38052
rect 29596 37998 29598 38050
rect 29598 37998 29650 38050
rect 29650 37998 29652 38050
rect 29596 37996 29652 37998
rect 30044 38050 30100 38052
rect 30044 37998 30046 38050
rect 30046 37998 30098 38050
rect 30098 37998 30100 38050
rect 30044 37996 30100 37998
rect 29932 37436 29988 37492
rect 29036 36316 29092 36372
rect 28140 36204 28196 36260
rect 28812 36204 28868 36260
rect 27692 35420 27748 35476
rect 28588 35586 28644 35588
rect 28588 35534 28590 35586
rect 28590 35534 28642 35586
rect 28642 35534 28644 35586
rect 28588 35532 28644 35534
rect 28588 35196 28644 35252
rect 28924 35532 28980 35588
rect 28252 34354 28308 34356
rect 28252 34302 28254 34354
rect 28254 34302 28306 34354
rect 28306 34302 28308 34354
rect 28252 34300 28308 34302
rect 27804 34130 27860 34132
rect 27804 34078 27806 34130
rect 27806 34078 27858 34130
rect 27858 34078 27860 34130
rect 27804 34076 27860 34078
rect 27804 33068 27860 33124
rect 27804 32674 27860 32676
rect 27804 32622 27806 32674
rect 27806 32622 27858 32674
rect 27858 32622 27860 32674
rect 27804 32620 27860 32622
rect 28364 34076 28420 34132
rect 28252 32284 28308 32340
rect 28476 32562 28532 32564
rect 28476 32510 28478 32562
rect 28478 32510 28530 32562
rect 28530 32510 28532 32562
rect 28476 32508 28532 32510
rect 28140 31836 28196 31892
rect 28700 34018 28756 34020
rect 28700 33966 28702 34018
rect 28702 33966 28754 34018
rect 28754 33966 28756 34018
rect 28700 33964 28756 33966
rect 28924 33628 28980 33684
rect 28924 32284 28980 32340
rect 28588 31836 28644 31892
rect 27692 31612 27748 31668
rect 27580 31500 27636 31556
rect 27468 30828 27524 30884
rect 26572 29932 26628 29988
rect 27356 29986 27412 29988
rect 27356 29934 27358 29986
rect 27358 29934 27410 29986
rect 27410 29934 27412 29986
rect 27356 29932 27412 29934
rect 27244 29820 27300 29876
rect 27132 29596 27188 29652
rect 26460 29484 26516 29540
rect 26460 28924 26516 28980
rect 27020 28924 27076 28980
rect 26012 27634 26068 27636
rect 26012 27582 26014 27634
rect 26014 27582 26066 27634
rect 26066 27582 26068 27634
rect 26012 27580 26068 27582
rect 26684 27074 26740 27076
rect 26684 27022 26686 27074
rect 26686 27022 26738 27074
rect 26738 27022 26740 27074
rect 26684 27020 26740 27022
rect 26348 26908 26404 26964
rect 25228 24108 25284 24164
rect 25564 26572 25620 26628
rect 25676 26796 25732 26852
rect 25900 24946 25956 24948
rect 25900 24894 25902 24946
rect 25902 24894 25954 24946
rect 25954 24894 25956 24946
rect 25900 24892 25956 24894
rect 25340 23436 25396 23492
rect 25676 24722 25732 24724
rect 25676 24670 25678 24722
rect 25678 24670 25730 24722
rect 25730 24670 25732 24722
rect 25676 24668 25732 24670
rect 25116 22482 25172 22484
rect 25116 22430 25118 22482
rect 25118 22430 25170 22482
rect 25170 22430 25172 22482
rect 25116 22428 25172 22430
rect 22988 21532 23044 21588
rect 23100 21644 23156 21700
rect 23324 21698 23380 21700
rect 23324 21646 23326 21698
rect 23326 21646 23378 21698
rect 23378 21646 23380 21698
rect 23324 21644 23380 21646
rect 22652 18396 22708 18452
rect 22764 18338 22820 18340
rect 22764 18286 22766 18338
rect 22766 18286 22818 18338
rect 22818 18286 22820 18338
rect 22764 18284 22820 18286
rect 23212 18562 23268 18564
rect 23212 18510 23214 18562
rect 23214 18510 23266 18562
rect 23266 18510 23268 18562
rect 23212 18508 23268 18510
rect 22652 17666 22708 17668
rect 22652 17614 22654 17666
rect 22654 17614 22706 17666
rect 22706 17614 22708 17666
rect 22652 17612 22708 17614
rect 22876 17836 22932 17892
rect 23212 17724 23268 17780
rect 22988 17106 23044 17108
rect 22988 17054 22990 17106
rect 22990 17054 23042 17106
rect 23042 17054 23044 17106
rect 22988 17052 23044 17054
rect 23212 16940 23268 16996
rect 22988 16882 23044 16884
rect 22988 16830 22990 16882
rect 22990 16830 23042 16882
rect 23042 16830 23044 16882
rect 22988 16828 23044 16830
rect 23212 16210 23268 16212
rect 23212 16158 23214 16210
rect 23214 16158 23266 16210
rect 23266 16158 23268 16210
rect 23212 16156 23268 16158
rect 22316 14476 22372 14532
rect 22316 13916 22372 13972
rect 22652 14530 22708 14532
rect 22652 14478 22654 14530
rect 22654 14478 22706 14530
rect 22706 14478 22708 14530
rect 22652 14476 22708 14478
rect 22988 13970 23044 13972
rect 22988 13918 22990 13970
rect 22990 13918 23042 13970
rect 23042 13918 23044 13970
rect 22988 13916 23044 13918
rect 23212 11788 23268 11844
rect 22876 11340 22932 11396
rect 22652 10780 22708 10836
rect 22540 9772 22596 9828
rect 22988 9772 23044 9828
rect 22876 9436 22932 9492
rect 23212 9436 23268 9492
rect 21980 8316 22036 8372
rect 22204 8204 22260 8260
rect 22764 8370 22820 8372
rect 22764 8318 22766 8370
rect 22766 8318 22818 8370
rect 22818 8318 22820 8370
rect 22764 8316 22820 8318
rect 22540 7868 22596 7924
rect 22092 7474 22148 7476
rect 22092 7422 22094 7474
rect 22094 7422 22146 7474
rect 22146 7422 22148 7474
rect 22092 7420 22148 7422
rect 23212 7420 23268 7476
rect 22316 7084 22372 7140
rect 22876 7084 22932 7140
rect 21420 6076 21476 6132
rect 20524 5122 20580 5124
rect 20524 5070 20526 5122
rect 20526 5070 20578 5122
rect 20578 5070 20580 5122
rect 20524 5068 20580 5070
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 21868 5122 21924 5124
rect 21868 5070 21870 5122
rect 21870 5070 21922 5122
rect 21922 5070 21924 5122
rect 21868 5068 21924 5070
rect 20636 4284 20692 4340
rect 21980 4732 22036 4788
rect 22428 4956 22484 5012
rect 23212 7196 23268 7252
rect 23436 21474 23492 21476
rect 23436 21422 23438 21474
rect 23438 21422 23490 21474
rect 23490 21422 23492 21474
rect 23436 21420 23492 21422
rect 24780 21698 24836 21700
rect 24780 21646 24782 21698
rect 24782 21646 24834 21698
rect 24834 21646 24836 21698
rect 24780 21644 24836 21646
rect 23436 20578 23492 20580
rect 23436 20526 23438 20578
rect 23438 20526 23490 20578
rect 23490 20526 23492 20578
rect 23436 20524 23492 20526
rect 23996 20578 24052 20580
rect 23996 20526 23998 20578
rect 23998 20526 24050 20578
rect 24050 20526 24052 20578
rect 23996 20524 24052 20526
rect 25788 24610 25844 24612
rect 25788 24558 25790 24610
rect 25790 24558 25842 24610
rect 25842 24558 25844 24610
rect 25788 24556 25844 24558
rect 26012 24332 26068 24388
rect 27356 29596 27412 29652
rect 27916 29372 27972 29428
rect 27692 27804 27748 27860
rect 27468 27074 27524 27076
rect 27468 27022 27470 27074
rect 27470 27022 27522 27074
rect 27522 27022 27524 27074
rect 27468 27020 27524 27022
rect 27580 27132 27636 27188
rect 27244 26962 27300 26964
rect 27244 26910 27246 26962
rect 27246 26910 27298 26962
rect 27298 26910 27300 26962
rect 27244 26908 27300 26910
rect 28140 27970 28196 27972
rect 28140 27918 28142 27970
rect 28142 27918 28194 27970
rect 28194 27918 28196 27970
rect 28140 27916 28196 27918
rect 28252 27132 28308 27188
rect 28028 27074 28084 27076
rect 28028 27022 28030 27074
rect 28030 27022 28082 27074
rect 28082 27022 28084 27074
rect 28364 31500 28420 31556
rect 28028 27020 28084 27022
rect 29596 36764 29652 36820
rect 29708 36370 29764 36372
rect 29708 36318 29710 36370
rect 29710 36318 29762 36370
rect 29762 36318 29764 36370
rect 29708 36316 29764 36318
rect 29596 36204 29652 36260
rect 30044 35586 30100 35588
rect 30044 35534 30046 35586
rect 30046 35534 30098 35586
rect 30098 35534 30100 35586
rect 30044 35532 30100 35534
rect 29932 35308 29988 35364
rect 29932 34130 29988 34132
rect 29932 34078 29934 34130
rect 29934 34078 29986 34130
rect 29986 34078 29988 34130
rect 29932 34076 29988 34078
rect 29372 33964 29428 34020
rect 29372 33628 29428 33684
rect 30492 44268 30548 44324
rect 30716 44098 30772 44100
rect 30716 44046 30718 44098
rect 30718 44046 30770 44098
rect 30770 44046 30772 44098
rect 30716 44044 30772 44046
rect 30604 43426 30660 43428
rect 30604 43374 30606 43426
rect 30606 43374 30658 43426
rect 30658 43374 30660 43426
rect 30604 43372 30660 43374
rect 30492 42642 30548 42644
rect 30492 42590 30494 42642
rect 30494 42590 30546 42642
rect 30546 42590 30548 42642
rect 30492 42588 30548 42590
rect 30716 42924 30772 42980
rect 30604 42028 30660 42084
rect 30380 40908 30436 40964
rect 30604 40962 30660 40964
rect 30604 40910 30606 40962
rect 30606 40910 30658 40962
rect 30658 40910 30660 40962
rect 30604 40908 30660 40910
rect 31164 50316 31220 50372
rect 30940 48972 30996 49028
rect 30940 48412 30996 48468
rect 30940 47964 30996 48020
rect 31276 50092 31332 50148
rect 31164 49196 31220 49252
rect 31164 48188 31220 48244
rect 30380 39004 30436 39060
rect 31052 45612 31108 45668
rect 31948 50764 32004 50820
rect 31724 50316 31780 50372
rect 32172 50428 32228 50484
rect 32060 50092 32116 50148
rect 31836 49698 31892 49700
rect 31836 49646 31838 49698
rect 31838 49646 31890 49698
rect 31890 49646 31892 49698
rect 31836 49644 31892 49646
rect 31836 48972 31892 49028
rect 31500 48914 31556 48916
rect 31500 48862 31502 48914
rect 31502 48862 31554 48914
rect 31554 48862 31556 48914
rect 31500 48860 31556 48862
rect 31836 48300 31892 48356
rect 31948 47570 32004 47572
rect 31948 47518 31950 47570
rect 31950 47518 32002 47570
rect 32002 47518 32004 47570
rect 31948 47516 32004 47518
rect 31500 47234 31556 47236
rect 31500 47182 31502 47234
rect 31502 47182 31554 47234
rect 31554 47182 31556 47234
rect 31500 47180 31556 47182
rect 31388 46844 31444 46900
rect 38220 58492 38276 58548
rect 36540 56364 36596 56420
rect 34412 56082 34468 56084
rect 34412 56030 34414 56082
rect 34414 56030 34466 56082
rect 34466 56030 34468 56082
rect 34412 56028 34468 56030
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 33964 55356 34020 55412
rect 34300 55298 34356 55300
rect 34300 55246 34302 55298
rect 34302 55246 34354 55298
rect 34354 55246 34356 55298
rect 34300 55244 34356 55246
rect 36988 55970 37044 55972
rect 36988 55918 36990 55970
rect 36990 55918 37042 55970
rect 37042 55918 37044 55970
rect 36988 55916 37044 55918
rect 37996 55692 38052 55748
rect 40124 58268 40180 58324
rect 38668 57820 38724 57876
rect 38332 57596 38388 57652
rect 36092 55186 36148 55188
rect 36092 55134 36094 55186
rect 36094 55134 36146 55186
rect 36146 55134 36148 55186
rect 36092 55132 36148 55134
rect 33852 54460 33908 54516
rect 34076 54348 34132 54404
rect 33404 54012 33460 54068
rect 33404 53676 33460 53732
rect 32732 53228 32788 53284
rect 32620 53116 32676 53172
rect 32396 51996 32452 52052
rect 32956 52050 33012 52052
rect 32956 51998 32958 52050
rect 32958 51998 33010 52050
rect 33010 51998 33012 52050
rect 32956 51996 33012 51998
rect 32396 51772 32452 51828
rect 33068 51772 33124 51828
rect 32508 51324 32564 51380
rect 32732 51154 32788 51156
rect 32732 51102 32734 51154
rect 32734 51102 32786 51154
rect 32786 51102 32788 51154
rect 32732 51100 32788 51102
rect 32620 50316 32676 50372
rect 31276 46674 31332 46676
rect 31276 46622 31278 46674
rect 31278 46622 31330 46674
rect 31330 46622 31332 46674
rect 31276 46620 31332 46622
rect 31724 46396 31780 46452
rect 31388 45612 31444 45668
rect 31164 45500 31220 45556
rect 32060 46562 32116 46564
rect 32060 46510 32062 46562
rect 32062 46510 32114 46562
rect 32114 46510 32116 46562
rect 32060 46508 32116 46510
rect 31724 45836 31780 45892
rect 31276 44882 31332 44884
rect 31276 44830 31278 44882
rect 31278 44830 31330 44882
rect 31330 44830 31332 44882
rect 31276 44828 31332 44830
rect 31052 41468 31108 41524
rect 31052 40962 31108 40964
rect 31052 40910 31054 40962
rect 31054 40910 31106 40962
rect 31106 40910 31108 40962
rect 31052 40908 31108 40910
rect 30268 35532 30324 35588
rect 30604 38050 30660 38052
rect 30604 37998 30606 38050
rect 30606 37998 30658 38050
rect 30658 37998 30660 38050
rect 30604 37996 30660 37998
rect 30492 36482 30548 36484
rect 30492 36430 30494 36482
rect 30494 36430 30546 36482
rect 30546 36430 30548 36482
rect 30492 36428 30548 36430
rect 30604 36258 30660 36260
rect 30604 36206 30606 36258
rect 30606 36206 30658 36258
rect 30658 36206 30660 36258
rect 30604 36204 30660 36206
rect 31164 40514 31220 40516
rect 31164 40462 31166 40514
rect 31166 40462 31218 40514
rect 31218 40462 31220 40514
rect 31164 40460 31220 40462
rect 31612 44716 31668 44772
rect 31500 43426 31556 43428
rect 31500 43374 31502 43426
rect 31502 43374 31554 43426
rect 31554 43374 31556 43426
rect 31500 43372 31556 43374
rect 30940 39842 30996 39844
rect 30940 39790 30942 39842
rect 30942 39790 30994 39842
rect 30994 39790 30996 39842
rect 30940 39788 30996 39790
rect 30828 38668 30884 38724
rect 30828 37884 30884 37940
rect 30828 36540 30884 36596
rect 30716 35586 30772 35588
rect 30716 35534 30718 35586
rect 30718 35534 30770 35586
rect 30770 35534 30772 35586
rect 30716 35532 30772 35534
rect 30492 34412 30548 34468
rect 30380 34130 30436 34132
rect 30380 34078 30382 34130
rect 30382 34078 30434 34130
rect 30434 34078 30436 34130
rect 30380 34076 30436 34078
rect 30268 33516 30324 33572
rect 30604 33628 30660 33684
rect 31052 38668 31108 38724
rect 31052 38444 31108 38500
rect 31836 44828 31892 44884
rect 32732 49644 32788 49700
rect 32620 48860 32676 48916
rect 32732 49084 32788 49140
rect 33404 53340 33460 53396
rect 33404 52444 33460 52500
rect 33964 53900 34020 53956
rect 34188 54236 34244 54292
rect 33740 53340 33796 53396
rect 33740 53170 33796 53172
rect 33740 53118 33742 53170
rect 33742 53118 33794 53170
rect 33794 53118 33796 53170
rect 33740 53116 33796 53118
rect 33292 52220 33348 52276
rect 33292 50092 33348 50148
rect 33404 51436 33460 51492
rect 32284 48636 32340 48692
rect 32284 48354 32340 48356
rect 32284 48302 32286 48354
rect 32286 48302 32338 48354
rect 32338 48302 32340 48354
rect 32284 48300 32340 48302
rect 33068 49026 33124 49028
rect 33068 48974 33070 49026
rect 33070 48974 33122 49026
rect 33122 48974 33124 49026
rect 33068 48972 33124 48974
rect 33180 48914 33236 48916
rect 33180 48862 33182 48914
rect 33182 48862 33234 48914
rect 33234 48862 33236 48914
rect 33180 48860 33236 48862
rect 32844 48636 32900 48692
rect 32620 48242 32676 48244
rect 32620 48190 32622 48242
rect 32622 48190 32674 48242
rect 32674 48190 32676 48242
rect 32620 48188 32676 48190
rect 32844 47458 32900 47460
rect 32844 47406 32846 47458
rect 32846 47406 32898 47458
rect 32898 47406 32900 47458
rect 32844 47404 32900 47406
rect 33180 47346 33236 47348
rect 33180 47294 33182 47346
rect 33182 47294 33234 47346
rect 33234 47294 33236 47346
rect 33180 47292 33236 47294
rect 32844 47068 32900 47124
rect 32508 46956 32564 47012
rect 32284 44156 32340 44212
rect 32172 44044 32228 44100
rect 31724 43596 31780 43652
rect 31836 43372 31892 43428
rect 32060 42924 32116 42980
rect 31500 39788 31556 39844
rect 31276 38444 31332 38500
rect 31388 37884 31444 37940
rect 30940 34300 30996 34356
rect 31276 36764 31332 36820
rect 31388 35532 31444 35588
rect 32284 43426 32340 43428
rect 32284 43374 32286 43426
rect 32286 43374 32338 43426
rect 32338 43374 32340 43426
rect 32284 43372 32340 43374
rect 31948 42082 32004 42084
rect 31948 42030 31950 42082
rect 31950 42030 32002 42082
rect 32002 42030 32004 42082
rect 31948 42028 32004 42030
rect 31836 41468 31892 41524
rect 31836 39506 31892 39508
rect 31836 39454 31838 39506
rect 31838 39454 31890 39506
rect 31890 39454 31892 39506
rect 31836 39452 31892 39454
rect 33068 47068 33124 47124
rect 32956 46002 33012 46004
rect 32956 45950 32958 46002
rect 32958 45950 33010 46002
rect 33010 45950 33012 46002
rect 32956 45948 33012 45950
rect 32956 44546 33012 44548
rect 32956 44494 32958 44546
rect 32958 44494 33010 44546
rect 33010 44494 33012 44546
rect 32956 44492 33012 44494
rect 32620 43596 32676 43652
rect 32620 43426 32676 43428
rect 32620 43374 32622 43426
rect 32622 43374 32674 43426
rect 32674 43374 32676 43426
rect 32620 43372 32676 43374
rect 33180 46956 33236 47012
rect 33180 45388 33236 45444
rect 34636 54572 34692 54628
rect 35196 55074 35252 55076
rect 35196 55022 35198 55074
rect 35198 55022 35250 55074
rect 35250 55022 35252 55074
rect 35196 55020 35252 55022
rect 35868 55020 35924 55076
rect 34860 54236 34916 54292
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 34636 53788 34692 53844
rect 34412 53340 34468 53396
rect 34748 53452 34804 53508
rect 33740 51772 33796 51828
rect 33852 51490 33908 51492
rect 33852 51438 33854 51490
rect 33854 51438 33906 51490
rect 33906 51438 33908 51490
rect 33852 51436 33908 51438
rect 33740 51378 33796 51380
rect 33740 51326 33742 51378
rect 33742 51326 33794 51378
rect 33794 51326 33796 51378
rect 33740 51324 33796 51326
rect 34412 52274 34468 52276
rect 34412 52222 34414 52274
rect 34414 52222 34466 52274
rect 34466 52222 34468 52274
rect 34412 52220 34468 52222
rect 36988 55020 37044 55076
rect 36204 54738 36260 54740
rect 36204 54686 36206 54738
rect 36206 54686 36258 54738
rect 36258 54686 36260 54738
rect 36204 54684 36260 54686
rect 35980 54236 36036 54292
rect 35644 53506 35700 53508
rect 35644 53454 35646 53506
rect 35646 53454 35698 53506
rect 35698 53454 35700 53506
rect 35644 53452 35700 53454
rect 35084 53340 35140 53396
rect 36092 53340 36148 53396
rect 36988 54290 37044 54292
rect 36988 54238 36990 54290
rect 36990 54238 37042 54290
rect 37042 54238 37044 54290
rect 36988 54236 37044 54238
rect 36876 53452 36932 53508
rect 36764 53340 36820 53396
rect 36764 53170 36820 53172
rect 36764 53118 36766 53170
rect 36766 53118 36818 53170
rect 36818 53118 36820 53170
rect 36764 53116 36820 53118
rect 36540 53058 36596 53060
rect 36540 53006 36542 53058
rect 36542 53006 36594 53058
rect 36594 53006 36596 53058
rect 36540 53004 36596 53006
rect 35980 52946 36036 52948
rect 35980 52894 35982 52946
rect 35982 52894 36034 52946
rect 36034 52894 36036 52946
rect 35980 52892 36036 52894
rect 34524 51436 34580 51492
rect 34076 51324 34132 51380
rect 33964 51212 34020 51268
rect 34860 51212 34916 51268
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35532 52108 35588 52164
rect 35868 52220 35924 52276
rect 35644 51378 35700 51380
rect 35644 51326 35646 51378
rect 35646 51326 35698 51378
rect 35698 51326 35700 51378
rect 35644 51324 35700 51326
rect 36092 51100 36148 51156
rect 34188 50818 34244 50820
rect 34188 50766 34190 50818
rect 34190 50766 34242 50818
rect 34242 50766 34244 50818
rect 34188 50764 34244 50766
rect 34524 50818 34580 50820
rect 34524 50766 34526 50818
rect 34526 50766 34578 50818
rect 34578 50766 34580 50818
rect 34524 50764 34580 50766
rect 34524 50594 34580 50596
rect 34524 50542 34526 50594
rect 34526 50542 34578 50594
rect 34578 50542 34580 50594
rect 34524 50540 34580 50542
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35532 50652 35588 50708
rect 35196 50540 35252 50596
rect 33964 49698 34020 49700
rect 33964 49646 33966 49698
rect 33966 49646 34018 49698
rect 34018 49646 34020 49698
rect 33964 49644 34020 49646
rect 36764 52162 36820 52164
rect 36764 52110 36766 52162
rect 36766 52110 36818 52162
rect 36818 52110 36820 52162
rect 36764 52108 36820 52110
rect 36652 51212 36708 51268
rect 36540 50764 36596 50820
rect 36428 50652 36484 50708
rect 36204 50594 36260 50596
rect 36204 50542 36206 50594
rect 36206 50542 36258 50594
rect 36258 50542 36260 50594
rect 36204 50540 36260 50542
rect 36540 50482 36596 50484
rect 36540 50430 36542 50482
rect 36542 50430 36594 50482
rect 36594 50430 36596 50482
rect 36540 50428 36596 50430
rect 33852 49138 33908 49140
rect 33852 49086 33854 49138
rect 33854 49086 33906 49138
rect 33906 49086 33908 49138
rect 33852 49084 33908 49086
rect 33516 48972 33572 49028
rect 34188 49026 34244 49028
rect 34188 48974 34190 49026
rect 34190 48974 34242 49026
rect 34242 48974 34244 49026
rect 34188 48972 34244 48974
rect 33852 48636 33908 48692
rect 33628 48242 33684 48244
rect 33628 48190 33630 48242
rect 33630 48190 33682 48242
rect 33682 48190 33684 48242
rect 33628 48188 33684 48190
rect 33964 48524 34020 48580
rect 34972 49084 35028 49140
rect 34860 48524 34916 48580
rect 33852 47458 33908 47460
rect 33852 47406 33854 47458
rect 33854 47406 33906 47458
rect 33906 47406 33908 47458
rect 33852 47404 33908 47406
rect 33628 47292 33684 47348
rect 33628 47068 33684 47124
rect 34300 47628 34356 47684
rect 34076 47346 34132 47348
rect 34076 47294 34078 47346
rect 34078 47294 34130 47346
rect 34130 47294 34132 47346
rect 34076 47292 34132 47294
rect 33404 45948 33460 46004
rect 33404 45388 33460 45444
rect 32508 42364 32564 42420
rect 32172 41468 32228 41524
rect 32396 42028 32452 42084
rect 32284 39452 32340 39508
rect 32844 41970 32900 41972
rect 32844 41918 32846 41970
rect 32846 41918 32898 41970
rect 32898 41918 32900 41970
rect 32844 41916 32900 41918
rect 32172 39004 32228 39060
rect 32060 37938 32116 37940
rect 32060 37886 32062 37938
rect 32062 37886 32114 37938
rect 32114 37886 32116 37938
rect 32060 37884 32116 37886
rect 31948 36594 32004 36596
rect 31948 36542 31950 36594
rect 31950 36542 32002 36594
rect 32002 36542 32004 36594
rect 31948 36540 32004 36542
rect 32060 35644 32116 35700
rect 31276 34300 31332 34356
rect 31164 34018 31220 34020
rect 31164 33966 31166 34018
rect 31166 33966 31218 34018
rect 31218 33966 31220 34018
rect 31164 33964 31220 33966
rect 30828 33292 30884 33348
rect 31052 33516 31108 33572
rect 29148 32060 29204 32116
rect 29260 31836 29316 31892
rect 28476 29650 28532 29652
rect 28476 29598 28478 29650
rect 28478 29598 28530 29650
rect 28530 29598 28532 29650
rect 28476 29596 28532 29598
rect 28588 27186 28644 27188
rect 28588 27134 28590 27186
rect 28590 27134 28642 27186
rect 28642 27134 28644 27186
rect 28588 27132 28644 27134
rect 29036 29932 29092 29988
rect 28812 29484 28868 29540
rect 28700 26460 28756 26516
rect 28476 26236 28532 26292
rect 28364 25900 28420 25956
rect 26460 24892 26516 24948
rect 27020 24892 27076 24948
rect 26908 24834 26964 24836
rect 26908 24782 26910 24834
rect 26910 24782 26962 24834
rect 26962 24782 26964 24834
rect 26908 24780 26964 24782
rect 26124 23996 26180 24052
rect 26236 23548 26292 23604
rect 26124 23436 26180 23492
rect 25676 23154 25732 23156
rect 25676 23102 25678 23154
rect 25678 23102 25730 23154
rect 25730 23102 25732 23154
rect 25676 23100 25732 23102
rect 26012 23100 26068 23156
rect 24108 20412 24164 20468
rect 24444 20524 24500 20580
rect 24332 20130 24388 20132
rect 24332 20078 24334 20130
rect 24334 20078 24386 20130
rect 24386 20078 24388 20130
rect 24332 20076 24388 20078
rect 23548 19906 23604 19908
rect 23548 19854 23550 19906
rect 23550 19854 23602 19906
rect 23602 19854 23604 19906
rect 23548 19852 23604 19854
rect 24444 19292 24500 19348
rect 25004 20690 25060 20692
rect 25004 20638 25006 20690
rect 25006 20638 25058 20690
rect 25058 20638 25060 20690
rect 25004 20636 25060 20638
rect 25564 20690 25620 20692
rect 25564 20638 25566 20690
rect 25566 20638 25618 20690
rect 25618 20638 25620 20690
rect 25564 20636 25620 20638
rect 24220 18508 24276 18564
rect 24780 20412 24836 20468
rect 25564 20130 25620 20132
rect 25564 20078 25566 20130
rect 25566 20078 25618 20130
rect 25618 20078 25620 20130
rect 25564 20076 25620 20078
rect 24332 18284 24388 18340
rect 24332 17724 24388 17780
rect 23884 17666 23940 17668
rect 23884 17614 23886 17666
rect 23886 17614 23938 17666
rect 23938 17614 23940 17666
rect 23884 17612 23940 17614
rect 24556 18172 24612 18228
rect 24892 17724 24948 17780
rect 24668 17500 24724 17556
rect 23996 17442 24052 17444
rect 23996 17390 23998 17442
rect 23998 17390 24050 17442
rect 24050 17390 24052 17442
rect 23996 17388 24052 17390
rect 23660 16940 23716 16996
rect 24220 16994 24276 16996
rect 24220 16942 24222 16994
rect 24222 16942 24274 16994
rect 24274 16942 24276 16994
rect 24220 16940 24276 16942
rect 24892 17164 24948 17220
rect 24668 16604 24724 16660
rect 23548 16044 23604 16100
rect 24108 16098 24164 16100
rect 24108 16046 24110 16098
rect 24110 16046 24162 16098
rect 24162 16046 24164 16098
rect 24108 16044 24164 16046
rect 24892 16156 24948 16212
rect 24108 15596 24164 15652
rect 23772 15484 23828 15540
rect 24444 15202 24500 15204
rect 24444 15150 24446 15202
rect 24446 15150 24498 15202
rect 24498 15150 24500 15202
rect 24444 15148 24500 15150
rect 23436 13916 23492 13972
rect 23436 13634 23492 13636
rect 23436 13582 23438 13634
rect 23438 13582 23490 13634
rect 23490 13582 23492 13634
rect 23436 13580 23492 13582
rect 24220 14530 24276 14532
rect 24220 14478 24222 14530
rect 24222 14478 24274 14530
rect 24274 14478 24276 14530
rect 24220 14476 24276 14478
rect 24108 14418 24164 14420
rect 24108 14366 24110 14418
rect 24110 14366 24162 14418
rect 24162 14366 24164 14418
rect 24108 14364 24164 14366
rect 24780 14028 24836 14084
rect 24556 13970 24612 13972
rect 24556 13918 24558 13970
rect 24558 13918 24610 13970
rect 24610 13918 24612 13970
rect 24556 13916 24612 13918
rect 24892 13580 24948 13636
rect 27804 25228 27860 25284
rect 27580 24946 27636 24948
rect 27580 24894 27582 24946
rect 27582 24894 27634 24946
rect 27634 24894 27636 24946
rect 27580 24892 27636 24894
rect 27804 24780 27860 24836
rect 27916 24722 27972 24724
rect 27916 24670 27918 24722
rect 27918 24670 27970 24722
rect 27970 24670 27972 24722
rect 27916 24668 27972 24670
rect 27804 24332 27860 24388
rect 26124 20636 26180 20692
rect 25900 20076 25956 20132
rect 26012 20524 26068 20580
rect 26460 20636 26516 20692
rect 26684 20636 26740 20692
rect 26684 20018 26740 20020
rect 26684 19966 26686 20018
rect 26686 19966 26738 20018
rect 26738 19966 26740 20018
rect 26684 19964 26740 19966
rect 26572 19628 26628 19684
rect 26572 19346 26628 19348
rect 26572 19294 26574 19346
rect 26574 19294 26626 19346
rect 26626 19294 26628 19346
rect 26572 19292 26628 19294
rect 26460 18844 26516 18900
rect 24668 12962 24724 12964
rect 24668 12910 24670 12962
rect 24670 12910 24722 12962
rect 24722 12910 24724 12962
rect 24668 12908 24724 12910
rect 24892 12908 24948 12964
rect 23772 11788 23828 11844
rect 23436 11676 23492 11732
rect 23996 11394 24052 11396
rect 23996 11342 23998 11394
rect 23998 11342 24050 11394
rect 24050 11342 24052 11394
rect 23996 11340 24052 11342
rect 25116 12962 25172 12964
rect 25116 12910 25118 12962
rect 25118 12910 25170 12962
rect 25170 12910 25172 12962
rect 25116 12908 25172 12910
rect 25340 17052 25396 17108
rect 25788 18226 25844 18228
rect 25788 18174 25790 18226
rect 25790 18174 25842 18226
rect 25842 18174 25844 18226
rect 25788 18172 25844 18174
rect 25900 18060 25956 18116
rect 25900 17612 25956 17668
rect 25452 16604 25508 16660
rect 25564 17164 25620 17220
rect 25900 17106 25956 17108
rect 25900 17054 25902 17106
rect 25902 17054 25954 17106
rect 25954 17054 25956 17106
rect 25900 17052 25956 17054
rect 25788 16828 25844 16884
rect 25676 16658 25732 16660
rect 25676 16606 25678 16658
rect 25678 16606 25730 16658
rect 25730 16606 25732 16658
rect 25676 16604 25732 16606
rect 25676 15036 25732 15092
rect 25564 14924 25620 14980
rect 25788 14530 25844 14532
rect 25788 14478 25790 14530
rect 25790 14478 25842 14530
rect 25842 14478 25844 14530
rect 25788 14476 25844 14478
rect 25340 14028 25396 14084
rect 25564 14028 25620 14084
rect 25452 13916 25508 13972
rect 24108 10780 24164 10836
rect 23996 10722 24052 10724
rect 23996 10670 23998 10722
rect 23998 10670 24050 10722
rect 24050 10670 24052 10722
rect 23996 10668 24052 10670
rect 25004 10556 25060 10612
rect 25228 10220 25284 10276
rect 25676 13580 25732 13636
rect 25676 13356 25732 13412
rect 25564 10332 25620 10388
rect 25452 10108 25508 10164
rect 24108 9826 24164 9828
rect 24108 9774 24110 9826
rect 24110 9774 24162 9826
rect 24162 9774 24164 9826
rect 24108 9772 24164 9774
rect 23772 9436 23828 9492
rect 24892 9436 24948 9492
rect 25228 9826 25284 9828
rect 25228 9774 25230 9826
rect 25230 9774 25282 9826
rect 25282 9774 25284 9826
rect 25228 9772 25284 9774
rect 25564 9772 25620 9828
rect 26572 18732 26628 18788
rect 26460 18562 26516 18564
rect 26460 18510 26462 18562
rect 26462 18510 26514 18562
rect 26514 18510 26516 18562
rect 26460 18508 26516 18510
rect 26124 18396 26180 18452
rect 26124 17836 26180 17892
rect 26124 17276 26180 17332
rect 26908 18620 26964 18676
rect 27132 23548 27188 23604
rect 27132 23324 27188 23380
rect 28028 23324 28084 23380
rect 28140 25228 28196 25284
rect 27244 23154 27300 23156
rect 27244 23102 27246 23154
rect 27246 23102 27298 23154
rect 27298 23102 27300 23154
rect 27244 23100 27300 23102
rect 28588 25282 28644 25284
rect 28588 25230 28590 25282
rect 28590 25230 28642 25282
rect 28642 25230 28644 25282
rect 28588 25228 28644 25230
rect 27244 20578 27300 20580
rect 27244 20526 27246 20578
rect 27246 20526 27298 20578
rect 27298 20526 27300 20578
rect 27244 20524 27300 20526
rect 27132 20188 27188 20244
rect 27692 19628 27748 19684
rect 28476 24444 28532 24500
rect 28924 23714 28980 23716
rect 28924 23662 28926 23714
rect 28926 23662 28978 23714
rect 28978 23662 28980 23714
rect 28924 23660 28980 23662
rect 28924 22370 28980 22372
rect 28924 22318 28926 22370
rect 28926 22318 28978 22370
rect 28978 22318 28980 22370
rect 28924 22316 28980 22318
rect 27916 20578 27972 20580
rect 27916 20526 27918 20578
rect 27918 20526 27970 20578
rect 27970 20526 27972 20578
rect 27916 20524 27972 20526
rect 28252 20412 28308 20468
rect 28140 20130 28196 20132
rect 28140 20078 28142 20130
rect 28142 20078 28194 20130
rect 28194 20078 28196 20130
rect 28140 20076 28196 20078
rect 28028 19740 28084 19796
rect 26796 17612 26852 17668
rect 26684 17442 26740 17444
rect 26684 17390 26686 17442
rect 26686 17390 26738 17442
rect 26738 17390 26740 17442
rect 26684 17388 26740 17390
rect 26460 17106 26516 17108
rect 26460 17054 26462 17106
rect 26462 17054 26514 17106
rect 26514 17054 26516 17106
rect 26460 17052 26516 17054
rect 26236 16940 26292 16996
rect 26236 14924 26292 14980
rect 26124 14252 26180 14308
rect 25900 12908 25956 12964
rect 26012 13970 26068 13972
rect 26012 13918 26014 13970
rect 26014 13918 26066 13970
rect 26066 13918 26068 13970
rect 26012 13916 26068 13918
rect 26236 13970 26292 13972
rect 26236 13918 26238 13970
rect 26238 13918 26290 13970
rect 26290 13918 26292 13970
rect 26236 13916 26292 13918
rect 26908 17276 26964 17332
rect 26348 13356 26404 13412
rect 26796 14530 26852 14532
rect 26796 14478 26798 14530
rect 26798 14478 26850 14530
rect 26850 14478 26852 14530
rect 26796 14476 26852 14478
rect 26684 14306 26740 14308
rect 26684 14254 26686 14306
rect 26686 14254 26738 14306
rect 26738 14254 26740 14306
rect 26684 14252 26740 14254
rect 27244 18620 27300 18676
rect 27580 18674 27636 18676
rect 27580 18622 27582 18674
rect 27582 18622 27634 18674
rect 27634 18622 27636 18674
rect 27580 18620 27636 18622
rect 27692 18562 27748 18564
rect 27692 18510 27694 18562
rect 27694 18510 27746 18562
rect 27746 18510 27748 18562
rect 27692 18508 27748 18510
rect 27804 18450 27860 18452
rect 27804 18398 27806 18450
rect 27806 18398 27858 18450
rect 27858 18398 27860 18450
rect 27804 18396 27860 18398
rect 28028 18284 28084 18340
rect 29484 31890 29540 31892
rect 29484 31838 29486 31890
rect 29486 31838 29538 31890
rect 29538 31838 29540 31890
rect 29484 31836 29540 31838
rect 29372 27804 29428 27860
rect 29372 27244 29428 27300
rect 29708 30098 29764 30100
rect 29708 30046 29710 30098
rect 29710 30046 29762 30098
rect 29762 30046 29764 30098
rect 29708 30044 29764 30046
rect 29596 29708 29652 29764
rect 29596 29036 29652 29092
rect 29820 29148 29876 29204
rect 30044 29650 30100 29652
rect 30044 29598 30046 29650
rect 30046 29598 30098 29650
rect 30098 29598 30100 29650
rect 30044 29596 30100 29598
rect 30044 28588 30100 28644
rect 30716 32956 30772 33012
rect 30380 32674 30436 32676
rect 30380 32622 30382 32674
rect 30382 32622 30434 32674
rect 30434 32622 30436 32674
rect 30380 32620 30436 32622
rect 30940 32620 30996 32676
rect 30380 32284 30436 32340
rect 30268 31612 30324 31668
rect 30268 30044 30324 30100
rect 30268 28924 30324 28980
rect 30492 31106 30548 31108
rect 30492 31054 30494 31106
rect 30494 31054 30546 31106
rect 30546 31054 30548 31106
rect 30492 31052 30548 31054
rect 30716 30044 30772 30100
rect 30828 29708 30884 29764
rect 30716 29650 30772 29652
rect 30716 29598 30718 29650
rect 30718 29598 30770 29650
rect 30770 29598 30772 29650
rect 30716 29596 30772 29598
rect 31388 32956 31444 33012
rect 31276 29986 31332 29988
rect 31276 29934 31278 29986
rect 31278 29934 31330 29986
rect 31330 29934 31332 29986
rect 31276 29932 31332 29934
rect 30492 29202 30548 29204
rect 30492 29150 30494 29202
rect 30494 29150 30546 29202
rect 30546 29150 30548 29202
rect 30492 29148 30548 29150
rect 30268 27916 30324 27972
rect 30380 27356 30436 27412
rect 30604 28754 30660 28756
rect 30604 28702 30606 28754
rect 30606 28702 30658 28754
rect 30658 28702 30660 28754
rect 30604 28700 30660 28702
rect 30492 27244 30548 27300
rect 30604 28476 30660 28532
rect 29148 23266 29204 23268
rect 29148 23214 29150 23266
rect 29150 23214 29202 23266
rect 29202 23214 29204 23266
rect 29148 23212 29204 23214
rect 29932 26290 29988 26292
rect 29932 26238 29934 26290
rect 29934 26238 29986 26290
rect 29986 26238 29988 26290
rect 29932 26236 29988 26238
rect 29708 25116 29764 25172
rect 29820 24892 29876 24948
rect 30044 24892 30100 24948
rect 30268 25116 30324 25172
rect 29708 24498 29764 24500
rect 29708 24446 29710 24498
rect 29710 24446 29762 24498
rect 29762 24446 29764 24498
rect 29708 24444 29764 24446
rect 30044 23714 30100 23716
rect 30044 23662 30046 23714
rect 30046 23662 30098 23714
rect 30098 23662 30100 23714
rect 30044 23660 30100 23662
rect 30604 26852 30660 26908
rect 30604 24892 30660 24948
rect 29596 22652 29652 22708
rect 29820 23212 29876 23268
rect 29260 22316 29316 22372
rect 29708 22370 29764 22372
rect 29708 22318 29710 22370
rect 29710 22318 29762 22370
rect 29762 22318 29764 22370
rect 29708 22316 29764 22318
rect 29484 22092 29540 22148
rect 28700 20076 28756 20132
rect 28364 19964 28420 20020
rect 28700 19852 28756 19908
rect 28700 19010 28756 19012
rect 28700 18958 28702 19010
rect 28702 18958 28754 19010
rect 28754 18958 28756 19010
rect 28700 18956 28756 18958
rect 28476 18732 28532 18788
rect 29932 22146 29988 22148
rect 29932 22094 29934 22146
rect 29934 22094 29986 22146
rect 29986 22094 29988 22146
rect 29932 22092 29988 22094
rect 29820 21868 29876 21924
rect 30156 22092 30212 22148
rect 30380 22540 30436 22596
rect 30044 21644 30100 21700
rect 30156 21868 30212 21924
rect 29932 20802 29988 20804
rect 29932 20750 29934 20802
rect 29934 20750 29986 20802
rect 29986 20750 29988 20802
rect 29932 20748 29988 20750
rect 30044 20300 30100 20356
rect 29932 20130 29988 20132
rect 29932 20078 29934 20130
rect 29934 20078 29986 20130
rect 29986 20078 29988 20130
rect 29932 20076 29988 20078
rect 29820 19852 29876 19908
rect 27580 17724 27636 17780
rect 27468 17500 27524 17556
rect 27132 15596 27188 15652
rect 27132 15372 27188 15428
rect 27020 13692 27076 13748
rect 26348 12460 26404 12516
rect 26124 11564 26180 11620
rect 25900 10610 25956 10612
rect 25900 10558 25902 10610
rect 25902 10558 25954 10610
rect 25954 10558 25956 10610
rect 25900 10556 25956 10558
rect 25788 10220 25844 10276
rect 26124 9996 26180 10052
rect 26236 10332 26292 10388
rect 24444 8428 24500 8484
rect 23548 8370 23604 8372
rect 23548 8318 23550 8370
rect 23550 8318 23602 8370
rect 23602 8318 23604 8370
rect 23548 8316 23604 8318
rect 24220 8316 24276 8372
rect 23436 7474 23492 7476
rect 23436 7422 23438 7474
rect 23438 7422 23490 7474
rect 23490 7422 23492 7474
rect 23436 7420 23492 7422
rect 23884 8092 23940 8148
rect 23660 7420 23716 7476
rect 24892 8316 24948 8372
rect 25004 8258 25060 8260
rect 25004 8206 25006 8258
rect 25006 8206 25058 8258
rect 25058 8206 25060 8258
rect 25004 8204 25060 8206
rect 25116 9548 25172 9604
rect 25116 8428 25172 8484
rect 26012 9826 26068 9828
rect 26012 9774 26014 9826
rect 26014 9774 26066 9826
rect 26066 9774 26068 9826
rect 26012 9772 26068 9774
rect 25676 9548 25732 9604
rect 25340 8370 25396 8372
rect 25340 8318 25342 8370
rect 25342 8318 25394 8370
rect 25394 8318 25396 8370
rect 25340 8316 25396 8318
rect 25676 7980 25732 8036
rect 24556 7474 24612 7476
rect 24556 7422 24558 7474
rect 24558 7422 24610 7474
rect 24610 7422 24612 7474
rect 24556 7420 24612 7422
rect 24668 7308 24724 7364
rect 24556 7250 24612 7252
rect 24556 7198 24558 7250
rect 24558 7198 24610 7250
rect 24610 7198 24612 7250
rect 24556 7196 24612 7198
rect 24556 6188 24612 6244
rect 23324 5516 23380 5572
rect 24108 5122 24164 5124
rect 24108 5070 24110 5122
rect 24110 5070 24162 5122
rect 24162 5070 24164 5122
rect 24108 5068 24164 5070
rect 24556 5068 24612 5124
rect 23100 4956 23156 5012
rect 23772 5010 23828 5012
rect 23772 4958 23774 5010
rect 23774 4958 23826 5010
rect 23826 4958 23828 5010
rect 23772 4956 23828 4958
rect 23996 5010 24052 5012
rect 23996 4958 23998 5010
rect 23998 4958 24050 5010
rect 24050 4958 24052 5010
rect 23996 4956 24052 4958
rect 22540 4898 22596 4900
rect 22540 4846 22542 4898
rect 22542 4846 22594 4898
rect 22594 4846 22596 4898
rect 22540 4844 22596 4846
rect 25452 5010 25508 5012
rect 25452 4958 25454 5010
rect 25454 4958 25506 5010
rect 25506 4958 25508 5010
rect 25452 4956 25508 4958
rect 25116 4844 25172 4900
rect 25340 4898 25396 4900
rect 25340 4846 25342 4898
rect 25342 4846 25394 4898
rect 25394 4846 25396 4898
rect 25340 4844 25396 4846
rect 23884 4732 23940 4788
rect 23660 4396 23716 4452
rect 23100 4338 23156 4340
rect 23100 4286 23102 4338
rect 23102 4286 23154 4338
rect 23154 4286 23156 4338
rect 23100 4284 23156 4286
rect 3164 2604 3220 2660
rect 5068 3442 5124 3444
rect 5068 3390 5070 3442
rect 5070 3390 5122 3442
rect 5122 3390 5124 3442
rect 5068 3388 5124 3390
rect 5852 3442 5908 3444
rect 5852 3390 5854 3442
rect 5854 3390 5906 3442
rect 5906 3390 5908 3442
rect 5852 3388 5908 3390
rect 1932 1820 1988 1876
rect 16828 3388 16884 3444
rect 17612 3442 17668 3444
rect 17612 3390 17614 3442
rect 17614 3390 17666 3442
rect 17666 3390 17668 3442
rect 17612 3388 17668 3390
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 25676 7474 25732 7476
rect 25676 7422 25678 7474
rect 25678 7422 25730 7474
rect 25730 7422 25732 7474
rect 25676 7420 25732 7422
rect 25900 8258 25956 8260
rect 25900 8206 25902 8258
rect 25902 8206 25954 8258
rect 25954 8206 25956 8258
rect 25900 8204 25956 8206
rect 26572 12460 26628 12516
rect 27580 17388 27636 17444
rect 27468 15484 27524 15540
rect 28028 17276 28084 17332
rect 27916 15538 27972 15540
rect 27916 15486 27918 15538
rect 27918 15486 27970 15538
rect 27970 15486 27972 15538
rect 27916 15484 27972 15486
rect 28252 17554 28308 17556
rect 28252 17502 28254 17554
rect 28254 17502 28306 17554
rect 28306 17502 28308 17554
rect 28252 17500 28308 17502
rect 28476 17554 28532 17556
rect 28476 17502 28478 17554
rect 28478 17502 28530 17554
rect 28530 17502 28532 17554
rect 28476 17500 28532 17502
rect 29260 18450 29316 18452
rect 29260 18398 29262 18450
rect 29262 18398 29314 18450
rect 29314 18398 29316 18450
rect 29260 18396 29316 18398
rect 28812 18338 28868 18340
rect 28812 18286 28814 18338
rect 28814 18286 28866 18338
rect 28866 18286 28868 18338
rect 28812 18284 28868 18286
rect 28812 17442 28868 17444
rect 28812 17390 28814 17442
rect 28814 17390 28866 17442
rect 28866 17390 28868 17442
rect 28812 17388 28868 17390
rect 28700 16828 28756 16884
rect 28364 15986 28420 15988
rect 28364 15934 28366 15986
rect 28366 15934 28418 15986
rect 28418 15934 28420 15986
rect 28364 15932 28420 15934
rect 28476 15596 28532 15652
rect 28252 15538 28308 15540
rect 28252 15486 28254 15538
rect 28254 15486 28306 15538
rect 28306 15486 28308 15538
rect 28252 15484 28308 15486
rect 27356 14530 27412 14532
rect 27356 14478 27358 14530
rect 27358 14478 27410 14530
rect 27410 14478 27412 14530
rect 27356 14476 27412 14478
rect 27468 14252 27524 14308
rect 28364 15260 28420 15316
rect 26460 10668 26516 10724
rect 26460 9772 26516 9828
rect 26124 8204 26180 8260
rect 26684 10556 26740 10612
rect 26684 9996 26740 10052
rect 27356 11900 27412 11956
rect 26796 9772 26852 9828
rect 27244 10386 27300 10388
rect 27244 10334 27246 10386
rect 27246 10334 27298 10386
rect 27298 10334 27300 10386
rect 27244 10332 27300 10334
rect 26684 9324 26740 9380
rect 27132 9324 27188 9380
rect 26908 9154 26964 9156
rect 26908 9102 26910 9154
rect 26910 9102 26962 9154
rect 26962 9102 26964 9154
rect 26908 9100 26964 9102
rect 26908 8258 26964 8260
rect 26908 8206 26910 8258
rect 26910 8206 26962 8258
rect 26962 8206 26964 8258
rect 26908 8204 26964 8206
rect 26796 8092 26852 8148
rect 25788 7362 25844 7364
rect 25788 7310 25790 7362
rect 25790 7310 25842 7362
rect 25842 7310 25844 7362
rect 25788 7308 25844 7310
rect 27132 6578 27188 6580
rect 27132 6526 27134 6578
rect 27134 6526 27186 6578
rect 27186 6526 27188 6578
rect 27132 6524 27188 6526
rect 27580 10668 27636 10724
rect 27468 9548 27524 9604
rect 27356 9100 27412 9156
rect 27804 13916 27860 13972
rect 27804 13746 27860 13748
rect 27804 13694 27806 13746
rect 27806 13694 27858 13746
rect 27858 13694 27860 13746
rect 27804 13692 27860 13694
rect 28252 14588 28308 14644
rect 28476 13746 28532 13748
rect 28476 13694 28478 13746
rect 28478 13694 28530 13746
rect 28530 13694 28532 13746
rect 28476 13692 28532 13694
rect 28700 15484 28756 15540
rect 28700 14642 28756 14644
rect 28700 14590 28702 14642
rect 28702 14590 28754 14642
rect 28754 14590 28756 14642
rect 28700 14588 28756 14590
rect 28812 15090 28868 15092
rect 28812 15038 28814 15090
rect 28814 15038 28866 15090
rect 28866 15038 28868 15090
rect 28812 15036 28868 15038
rect 28812 13692 28868 13748
rect 28028 9884 28084 9940
rect 28700 13580 28756 13636
rect 28588 13074 28644 13076
rect 28588 13022 28590 13074
rect 28590 13022 28642 13074
rect 28642 13022 28644 13074
rect 28588 13020 28644 13022
rect 28588 12684 28644 12740
rect 28812 12850 28868 12852
rect 28812 12798 28814 12850
rect 28814 12798 28866 12850
rect 28866 12798 28868 12850
rect 28812 12796 28868 12798
rect 28364 10834 28420 10836
rect 28364 10782 28366 10834
rect 28366 10782 28418 10834
rect 28418 10782 28420 10834
rect 28364 10780 28420 10782
rect 28140 9772 28196 9828
rect 29820 18620 29876 18676
rect 29596 18172 29652 18228
rect 29484 17554 29540 17556
rect 29484 17502 29486 17554
rect 29486 17502 29538 17554
rect 29538 17502 29540 17554
rect 29484 17500 29540 17502
rect 29708 17554 29764 17556
rect 29708 17502 29710 17554
rect 29710 17502 29762 17554
rect 29762 17502 29764 17554
rect 29708 17500 29764 17502
rect 29932 17500 29988 17556
rect 29484 16828 29540 16884
rect 29148 15932 29204 15988
rect 30828 28924 30884 28980
rect 30940 28642 30996 28644
rect 30940 28590 30942 28642
rect 30942 28590 30994 28642
rect 30994 28590 30996 28642
rect 30940 28588 30996 28590
rect 31724 34636 31780 34692
rect 31836 34076 31892 34132
rect 31612 33628 31668 33684
rect 31724 33180 31780 33236
rect 31612 32508 31668 32564
rect 32508 39116 32564 39172
rect 32620 39788 32676 39844
rect 32508 38946 32564 38948
rect 32508 38894 32510 38946
rect 32510 38894 32562 38946
rect 32562 38894 32564 38946
rect 32508 38892 32564 38894
rect 32844 41468 32900 41524
rect 32956 39452 33012 39508
rect 32284 38444 32340 38500
rect 33068 38050 33124 38052
rect 33068 37998 33070 38050
rect 33070 37998 33122 38050
rect 33122 37998 33124 38050
rect 33068 37996 33124 37998
rect 32844 36428 32900 36484
rect 33292 44156 33348 44212
rect 33180 36370 33236 36372
rect 33180 36318 33182 36370
rect 33182 36318 33234 36370
rect 33234 36318 33236 36370
rect 33180 36316 33236 36318
rect 33068 36092 33124 36148
rect 32732 35810 32788 35812
rect 32732 35758 32734 35810
rect 32734 35758 32786 35810
rect 32786 35758 32788 35810
rect 32732 35756 32788 35758
rect 32620 35698 32676 35700
rect 32620 35646 32622 35698
rect 32622 35646 32674 35698
rect 32674 35646 32676 35698
rect 32620 35644 32676 35646
rect 32508 34914 32564 34916
rect 32508 34862 32510 34914
rect 32510 34862 32562 34914
rect 32562 34862 32564 34914
rect 32508 34860 32564 34862
rect 32732 34636 32788 34692
rect 32732 34354 32788 34356
rect 32732 34302 32734 34354
rect 32734 34302 32786 34354
rect 32786 34302 32788 34354
rect 32732 34300 32788 34302
rect 32396 33122 32452 33124
rect 32396 33070 32398 33122
rect 32398 33070 32450 33122
rect 32450 33070 32452 33122
rect 32396 33068 32452 33070
rect 32284 32956 32340 33012
rect 32172 31164 32228 31220
rect 31724 31052 31780 31108
rect 32060 31106 32116 31108
rect 32060 31054 32062 31106
rect 32062 31054 32114 31106
rect 32114 31054 32116 31106
rect 32060 31052 32116 31054
rect 31612 30882 31668 30884
rect 31612 30830 31614 30882
rect 31614 30830 31666 30882
rect 31666 30830 31668 30882
rect 31612 30828 31668 30830
rect 31948 30268 32004 30324
rect 31836 29932 31892 29988
rect 31724 28700 31780 28756
rect 31164 27356 31220 27412
rect 31164 27132 31220 27188
rect 30828 26908 30884 26964
rect 32172 28476 32228 28532
rect 32284 28588 32340 28644
rect 32060 28418 32116 28420
rect 32060 28366 32062 28418
rect 32062 28366 32114 28418
rect 32114 28366 32116 28418
rect 32060 28364 32116 28366
rect 31948 27468 32004 27524
rect 31388 27244 31444 27300
rect 32956 31948 33012 32004
rect 33628 45106 33684 45108
rect 33628 45054 33630 45106
rect 33630 45054 33682 45106
rect 33682 45054 33684 45106
rect 33628 45052 33684 45054
rect 33516 44492 33572 44548
rect 33516 44098 33572 44100
rect 33516 44046 33518 44098
rect 33518 44046 33570 44098
rect 33570 44046 33572 44098
rect 33516 44044 33572 44046
rect 33516 42924 33572 42980
rect 33852 45666 33908 45668
rect 33852 45614 33854 45666
rect 33854 45614 33906 45666
rect 33906 45614 33908 45666
rect 33852 45612 33908 45614
rect 33740 41916 33796 41972
rect 33852 45388 33908 45444
rect 33964 45052 34020 45108
rect 33964 42082 34020 42084
rect 33964 42030 33966 42082
rect 33966 42030 34018 42082
rect 34018 42030 34020 42082
rect 33964 42028 34020 42030
rect 33852 40684 33908 40740
rect 33964 40514 34020 40516
rect 33964 40462 33966 40514
rect 33966 40462 34018 40514
rect 34018 40462 34020 40514
rect 33964 40460 34020 40462
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35084 48972 35140 49028
rect 34860 47628 34916 47684
rect 34300 47068 34356 47124
rect 35308 48130 35364 48132
rect 35308 48078 35310 48130
rect 35310 48078 35362 48130
rect 35362 48078 35364 48130
rect 35308 48076 35364 48078
rect 35532 48802 35588 48804
rect 35532 48750 35534 48802
rect 35534 48750 35586 48802
rect 35586 48750 35588 48802
rect 35532 48748 35588 48750
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35196 47458 35252 47460
rect 35196 47406 35198 47458
rect 35198 47406 35250 47458
rect 35250 47406 35252 47458
rect 35196 47404 35252 47406
rect 35532 47458 35588 47460
rect 35532 47406 35534 47458
rect 35534 47406 35586 47458
rect 35586 47406 35588 47458
rect 35532 47404 35588 47406
rect 35420 47180 35476 47236
rect 35084 46956 35140 47012
rect 34412 46898 34468 46900
rect 34412 46846 34414 46898
rect 34414 46846 34466 46898
rect 34466 46846 34468 46898
rect 34412 46844 34468 46846
rect 34636 46844 34692 46900
rect 35308 46562 35364 46564
rect 35308 46510 35310 46562
rect 35310 46510 35362 46562
rect 35362 46510 35364 46562
rect 35308 46508 35364 46510
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 34860 45948 34916 46004
rect 34636 45388 34692 45444
rect 34524 45276 34580 45332
rect 35308 45778 35364 45780
rect 35308 45726 35310 45778
rect 35310 45726 35362 45778
rect 35362 45726 35364 45778
rect 35308 45724 35364 45726
rect 34860 45164 34916 45220
rect 34524 45106 34580 45108
rect 34524 45054 34526 45106
rect 34526 45054 34578 45106
rect 34578 45054 34580 45106
rect 34524 45052 34580 45054
rect 34972 45106 35028 45108
rect 34972 45054 34974 45106
rect 34974 45054 35026 45106
rect 35026 45054 35028 45106
rect 34972 45052 35028 45054
rect 35532 45106 35588 45108
rect 35532 45054 35534 45106
rect 35534 45054 35586 45106
rect 35586 45054 35588 45106
rect 35532 45052 35588 45054
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 36316 49868 36372 49924
rect 36316 48972 36372 49028
rect 35868 48466 35924 48468
rect 35868 48414 35870 48466
rect 35870 48414 35922 48466
rect 35922 48414 35924 48466
rect 35868 48412 35924 48414
rect 36428 48412 36484 48468
rect 36876 51154 36932 51156
rect 36876 51102 36878 51154
rect 36878 51102 36930 51154
rect 36930 51102 36932 51154
rect 36876 51100 36932 51102
rect 36764 49420 36820 49476
rect 37772 54626 37828 54628
rect 37772 54574 37774 54626
rect 37774 54574 37826 54626
rect 37826 54574 37828 54626
rect 37772 54572 37828 54574
rect 37324 53676 37380 53732
rect 37436 53788 37492 53844
rect 37324 53340 37380 53396
rect 37660 53340 37716 53396
rect 37772 53116 37828 53172
rect 38220 53058 38276 53060
rect 38220 53006 38222 53058
rect 38222 53006 38274 53058
rect 38274 53006 38276 53058
rect 38220 53004 38276 53006
rect 37436 52780 37492 52836
rect 37548 52332 37604 52388
rect 37660 51996 37716 52052
rect 37212 51548 37268 51604
rect 38108 51884 38164 51940
rect 37436 50706 37492 50708
rect 37436 50654 37438 50706
rect 37438 50654 37490 50706
rect 37490 50654 37492 50706
rect 37436 50652 37492 50654
rect 37324 50540 37380 50596
rect 38220 51324 38276 51380
rect 38444 55020 38500 55076
rect 39228 57708 39284 57764
rect 38780 56364 38836 56420
rect 39116 55468 39172 55524
rect 38892 55244 38948 55300
rect 38780 54572 38836 54628
rect 39452 56306 39508 56308
rect 39452 56254 39454 56306
rect 39454 56254 39506 56306
rect 39506 56254 39508 56306
rect 39452 56252 39508 56254
rect 39788 55916 39844 55972
rect 42812 57932 42868 57988
rect 40684 57260 40740 57316
rect 40236 55970 40292 55972
rect 40236 55918 40238 55970
rect 40238 55918 40290 55970
rect 40290 55918 40292 55970
rect 40236 55916 40292 55918
rect 39564 55244 39620 55300
rect 39340 54684 39396 54740
rect 39340 54514 39396 54516
rect 39340 54462 39342 54514
rect 39342 54462 39394 54514
rect 39394 54462 39396 54514
rect 39340 54460 39396 54462
rect 40012 55298 40068 55300
rect 40012 55246 40014 55298
rect 40014 55246 40066 55298
rect 40066 55246 40068 55298
rect 40012 55244 40068 55246
rect 39900 55074 39956 55076
rect 39900 55022 39902 55074
rect 39902 55022 39954 55074
rect 39954 55022 39956 55074
rect 39900 55020 39956 55022
rect 39788 53842 39844 53844
rect 39788 53790 39790 53842
rect 39790 53790 39842 53842
rect 39842 53790 39844 53842
rect 39788 53788 39844 53790
rect 40124 54236 40180 54292
rect 40012 53676 40068 53732
rect 39900 53618 39956 53620
rect 39900 53566 39902 53618
rect 39902 53566 39954 53618
rect 39954 53566 39956 53618
rect 39900 53564 39956 53566
rect 38668 52834 38724 52836
rect 38668 52782 38670 52834
rect 38670 52782 38722 52834
rect 38722 52782 38724 52834
rect 38668 52780 38724 52782
rect 38444 52050 38500 52052
rect 38444 51998 38446 52050
rect 38446 51998 38498 52050
rect 38498 51998 38500 52050
rect 38444 51996 38500 51998
rect 38556 51938 38612 51940
rect 38556 51886 38558 51938
rect 38558 51886 38610 51938
rect 38610 51886 38612 51938
rect 38556 51884 38612 51886
rect 38108 50876 38164 50932
rect 37100 49084 37156 49140
rect 37884 50034 37940 50036
rect 37884 49982 37886 50034
rect 37886 49982 37938 50034
rect 37938 49982 37940 50034
rect 37884 49980 37940 49982
rect 38332 50482 38388 50484
rect 38332 50430 38334 50482
rect 38334 50430 38386 50482
rect 38386 50430 38388 50482
rect 38332 50428 38388 50430
rect 38780 50204 38836 50260
rect 38220 49980 38276 50036
rect 39228 50204 39284 50260
rect 36988 48860 37044 48916
rect 36876 48524 36932 48580
rect 35756 46732 35812 46788
rect 35980 47180 36036 47236
rect 38220 49698 38276 49700
rect 38220 49646 38222 49698
rect 38222 49646 38274 49698
rect 38274 49646 38276 49698
rect 38220 49644 38276 49646
rect 38668 49420 38724 49476
rect 37772 49026 37828 49028
rect 37772 48974 37774 49026
rect 37774 48974 37826 49026
rect 37826 48974 37828 49026
rect 37772 48972 37828 48974
rect 38108 48972 38164 49028
rect 37884 48636 37940 48692
rect 38108 48412 38164 48468
rect 36988 48076 37044 48132
rect 36540 47516 36596 47572
rect 35756 45276 35812 45332
rect 35644 44604 35700 44660
rect 35644 44434 35700 44436
rect 35644 44382 35646 44434
rect 35646 44382 35698 44434
rect 35698 44382 35700 44434
rect 35644 44380 35700 44382
rect 36652 47404 36708 47460
rect 36764 47852 36820 47908
rect 36652 47068 36708 47124
rect 36428 45890 36484 45892
rect 36428 45838 36430 45890
rect 36430 45838 36482 45890
rect 36482 45838 36484 45890
rect 36428 45836 36484 45838
rect 36540 45666 36596 45668
rect 36540 45614 36542 45666
rect 36542 45614 36594 45666
rect 36594 45614 36596 45666
rect 36540 45612 36596 45614
rect 36988 47068 37044 47124
rect 36876 46732 36932 46788
rect 36092 44882 36148 44884
rect 36092 44830 36094 44882
rect 36094 44830 36146 44882
rect 36146 44830 36148 44882
rect 36092 44828 36148 44830
rect 34412 43596 34468 43652
rect 34188 43372 34244 43428
rect 34636 43538 34692 43540
rect 34636 43486 34638 43538
rect 34638 43486 34690 43538
rect 34690 43486 34692 43538
rect 34636 43484 34692 43486
rect 34972 43484 35028 43540
rect 34524 43372 34580 43428
rect 34860 43260 34916 43316
rect 34636 42754 34692 42756
rect 34636 42702 34638 42754
rect 34638 42702 34690 42754
rect 34690 42702 34692 42754
rect 34636 42700 34692 42702
rect 34412 42642 34468 42644
rect 34412 42590 34414 42642
rect 34414 42590 34466 42642
rect 34466 42590 34468 42642
rect 34412 42588 34468 42590
rect 35868 43314 35924 43316
rect 35868 43262 35870 43314
rect 35870 43262 35922 43314
rect 35922 43262 35924 43314
rect 35868 43260 35924 43262
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 34860 42476 34916 42532
rect 34188 42252 34244 42308
rect 34972 42364 35028 42420
rect 35196 42924 35252 42980
rect 36204 43314 36260 43316
rect 36204 43262 36206 43314
rect 36206 43262 36258 43314
rect 36258 43262 36260 43314
rect 36204 43260 36260 43262
rect 36092 43148 36148 43204
rect 36652 45388 36708 45444
rect 36764 44322 36820 44324
rect 36764 44270 36766 44322
rect 36766 44270 36818 44322
rect 36818 44270 36820 44322
rect 36764 44268 36820 44270
rect 36652 43820 36708 43876
rect 36652 43148 36708 43204
rect 36316 42924 36372 42980
rect 34300 42082 34356 42084
rect 34300 42030 34302 42082
rect 34302 42030 34354 42082
rect 34354 42030 34356 42082
rect 34300 42028 34356 42030
rect 34860 40572 34916 40628
rect 34636 40514 34692 40516
rect 34636 40462 34638 40514
rect 34638 40462 34690 40514
rect 34690 40462 34692 40514
rect 34636 40460 34692 40462
rect 34188 40236 34244 40292
rect 33740 38892 33796 38948
rect 33516 38444 33572 38500
rect 33964 38050 34020 38052
rect 33964 37998 33966 38050
rect 33966 37998 34018 38050
rect 34018 37998 34020 38050
rect 33964 37996 34020 37998
rect 33964 36652 34020 36708
rect 33628 36482 33684 36484
rect 33628 36430 33630 36482
rect 33630 36430 33682 36482
rect 33682 36430 33684 36482
rect 33628 36428 33684 36430
rect 33740 36370 33796 36372
rect 33740 36318 33742 36370
rect 33742 36318 33794 36370
rect 33794 36318 33796 36370
rect 33740 36316 33796 36318
rect 33740 36092 33796 36148
rect 33628 35756 33684 35812
rect 33964 36092 34020 36148
rect 35756 42642 35812 42644
rect 35756 42590 35758 42642
rect 35758 42590 35810 42642
rect 35810 42590 35812 42642
rect 35756 42588 35812 42590
rect 35980 42642 36036 42644
rect 35980 42590 35982 42642
rect 35982 42590 36034 42642
rect 36034 42590 36036 42642
rect 35980 42588 36036 42590
rect 35756 42140 35812 42196
rect 35420 42028 35476 42084
rect 35644 42028 35700 42084
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35868 42082 35924 42084
rect 35868 42030 35870 42082
rect 35870 42030 35922 42082
rect 35922 42030 35924 42082
rect 35868 42028 35924 42030
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 34972 38892 35028 38948
rect 35532 38892 35588 38948
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 33852 35698 33908 35700
rect 33852 35646 33854 35698
rect 33854 35646 33906 35698
rect 33906 35646 33908 35698
rect 33852 35644 33908 35646
rect 33964 35532 34020 35588
rect 33404 33346 33460 33348
rect 33404 33294 33406 33346
rect 33406 33294 33458 33346
rect 33458 33294 33460 33346
rect 33404 33292 33460 33294
rect 33516 32562 33572 32564
rect 33516 32510 33518 32562
rect 33518 32510 33570 32562
rect 33570 32510 33572 32562
rect 33516 32508 33572 32510
rect 33180 31164 33236 31220
rect 33404 32284 33460 32340
rect 33180 30828 33236 30884
rect 32844 29372 32900 29428
rect 32732 28642 32788 28644
rect 32732 28590 32734 28642
rect 32734 28590 32786 28642
rect 32786 28590 32788 28642
rect 32732 28588 32788 28590
rect 32172 26850 32228 26852
rect 32172 26798 32174 26850
rect 32174 26798 32226 26850
rect 32226 26798 32228 26850
rect 32172 26796 32228 26798
rect 32508 28364 32564 28420
rect 31276 26012 31332 26068
rect 32060 26402 32116 26404
rect 32060 26350 32062 26402
rect 32062 26350 32114 26402
rect 32114 26350 32116 26402
rect 32060 26348 32116 26350
rect 31500 25452 31556 25508
rect 32508 26290 32564 26292
rect 32508 26238 32510 26290
rect 32510 26238 32562 26290
rect 32562 26238 32564 26290
rect 32508 26236 32564 26238
rect 32284 25788 32340 25844
rect 32732 25788 32788 25844
rect 32844 26796 32900 26852
rect 32620 25676 32676 25732
rect 31836 25394 31892 25396
rect 31836 25342 31838 25394
rect 31838 25342 31890 25394
rect 31890 25342 31892 25394
rect 31836 25340 31892 25342
rect 32396 25394 32452 25396
rect 32396 25342 32398 25394
rect 32398 25342 32450 25394
rect 32450 25342 32452 25394
rect 32396 25340 32452 25342
rect 32732 25394 32788 25396
rect 32732 25342 32734 25394
rect 32734 25342 32786 25394
rect 32786 25342 32788 25394
rect 32732 25340 32788 25342
rect 35084 37212 35140 37268
rect 34748 36316 34804 36372
rect 34860 36652 34916 36708
rect 34636 36092 34692 36148
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35420 36428 35476 36484
rect 35420 35868 35476 35924
rect 35644 37266 35700 37268
rect 35644 37214 35646 37266
rect 35646 37214 35698 37266
rect 35698 37214 35700 37266
rect 35644 37212 35700 37214
rect 36316 42028 36372 42084
rect 36988 45836 37044 45892
rect 36988 44380 37044 44436
rect 36540 42082 36596 42084
rect 36540 42030 36542 42082
rect 36542 42030 36594 42082
rect 36594 42030 36596 42082
rect 36540 42028 36596 42030
rect 37548 48130 37604 48132
rect 37548 48078 37550 48130
rect 37550 48078 37602 48130
rect 37602 48078 37604 48130
rect 37548 48076 37604 48078
rect 38556 48354 38612 48356
rect 38556 48302 38558 48354
rect 38558 48302 38610 48354
rect 38610 48302 38612 48354
rect 38556 48300 38612 48302
rect 37212 47404 37268 47460
rect 37436 46956 37492 47012
rect 37884 47570 37940 47572
rect 37884 47518 37886 47570
rect 37886 47518 37938 47570
rect 37938 47518 37940 47570
rect 37884 47516 37940 47518
rect 37884 47068 37940 47124
rect 37772 46956 37828 47012
rect 37548 45666 37604 45668
rect 37548 45614 37550 45666
rect 37550 45614 37602 45666
rect 37602 45614 37604 45666
rect 37548 45612 37604 45614
rect 37324 44268 37380 44324
rect 37212 43762 37268 43764
rect 37212 43710 37214 43762
rect 37214 43710 37266 43762
rect 37266 43710 37268 43762
rect 37212 43708 37268 43710
rect 37436 42252 37492 42308
rect 36876 41804 36932 41860
rect 36540 40626 36596 40628
rect 36540 40574 36542 40626
rect 36542 40574 36594 40626
rect 36594 40574 36596 40626
rect 36540 40572 36596 40574
rect 37100 40908 37156 40964
rect 36876 40402 36932 40404
rect 36876 40350 36878 40402
rect 36878 40350 36930 40402
rect 36930 40350 36932 40402
rect 36876 40348 36932 40350
rect 36876 39788 36932 39844
rect 36876 39004 36932 39060
rect 36988 39116 37044 39172
rect 35756 36540 35812 36596
rect 34412 35532 34468 35588
rect 36092 35922 36148 35924
rect 36092 35870 36094 35922
rect 36094 35870 36146 35922
rect 36146 35870 36148 35922
rect 36092 35868 36148 35870
rect 34972 35532 35028 35588
rect 35868 35532 35924 35588
rect 34860 35420 34916 35476
rect 35644 35420 35700 35476
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 34188 34636 34244 34692
rect 33740 33068 33796 33124
rect 33628 31724 33684 31780
rect 33852 31948 33908 32004
rect 34076 33068 34132 33124
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 36764 38162 36820 38164
rect 36764 38110 36766 38162
rect 36766 38110 36818 38162
rect 36818 38110 36820 38162
rect 36764 38108 36820 38110
rect 36988 36652 37044 36708
rect 36764 36370 36820 36372
rect 36764 36318 36766 36370
rect 36766 36318 36818 36370
rect 36818 36318 36820 36370
rect 36764 36316 36820 36318
rect 38108 47458 38164 47460
rect 38108 47406 38110 47458
rect 38110 47406 38162 47458
rect 38162 47406 38164 47458
rect 38108 47404 38164 47406
rect 38220 47068 38276 47124
rect 38108 46396 38164 46452
rect 37660 43538 37716 43540
rect 37660 43486 37662 43538
rect 37662 43486 37714 43538
rect 37714 43486 37716 43538
rect 37660 43484 37716 43486
rect 37996 43762 38052 43764
rect 37996 43710 37998 43762
rect 37998 43710 38050 43762
rect 38050 43710 38052 43762
rect 37996 43708 38052 43710
rect 37884 43484 37940 43540
rect 37772 42252 37828 42308
rect 37660 42140 37716 42196
rect 38108 42700 38164 42756
rect 38556 47068 38612 47124
rect 38332 46956 38388 47012
rect 38668 46844 38724 46900
rect 39788 51602 39844 51604
rect 39788 51550 39790 51602
rect 39790 51550 39842 51602
rect 39842 51550 39844 51602
rect 39788 51548 39844 51550
rect 40348 54684 40404 54740
rect 40460 52162 40516 52164
rect 40460 52110 40462 52162
rect 40462 52110 40514 52162
rect 40514 52110 40516 52162
rect 40460 52108 40516 52110
rect 41804 55692 41860 55748
rect 41244 55074 41300 55076
rect 41244 55022 41246 55074
rect 41246 55022 41298 55074
rect 41298 55022 41300 55074
rect 41244 55020 41300 55022
rect 41132 54236 41188 54292
rect 40908 53618 40964 53620
rect 40908 53566 40910 53618
rect 40910 53566 40962 53618
rect 40962 53566 40964 53618
rect 40908 53564 40964 53566
rect 41468 54124 41524 54180
rect 42252 54684 42308 54740
rect 42364 55916 42420 55972
rect 42140 54572 42196 54628
rect 42028 54514 42084 54516
rect 42028 54462 42030 54514
rect 42030 54462 42082 54514
rect 42082 54462 42084 54514
rect 42028 54460 42084 54462
rect 42140 53900 42196 53956
rect 43596 56194 43652 56196
rect 43596 56142 43598 56194
rect 43598 56142 43650 56194
rect 43650 56142 43652 56194
rect 43596 56140 43652 56142
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 46396 56140 46452 56196
rect 47292 56140 47348 56196
rect 42812 55580 42868 55636
rect 43484 55804 43540 55860
rect 43148 55298 43204 55300
rect 43148 55246 43150 55298
rect 43150 55246 43202 55298
rect 43202 55246 43204 55298
rect 43148 55244 43204 55246
rect 42476 55186 42532 55188
rect 42476 55134 42478 55186
rect 42478 55134 42530 55186
rect 42530 55134 42532 55186
rect 42476 55132 42532 55134
rect 43036 55020 43092 55076
rect 43148 54124 43204 54180
rect 40796 53058 40852 53060
rect 40796 53006 40798 53058
rect 40798 53006 40850 53058
rect 40850 53006 40852 53058
rect 40796 53004 40852 53006
rect 40572 51660 40628 51716
rect 39676 51378 39732 51380
rect 39676 51326 39678 51378
rect 39678 51326 39730 51378
rect 39730 51326 39732 51378
rect 39676 51324 39732 51326
rect 39564 50204 39620 50260
rect 39564 50034 39620 50036
rect 39564 49982 39566 50034
rect 39566 49982 39618 50034
rect 39618 49982 39620 50034
rect 39564 49980 39620 49982
rect 39452 49532 39508 49588
rect 39788 48972 39844 49028
rect 38892 48466 38948 48468
rect 38892 48414 38894 48466
rect 38894 48414 38946 48466
rect 38946 48414 38948 48466
rect 38892 48412 38948 48414
rect 40236 49698 40292 49700
rect 40236 49646 40238 49698
rect 40238 49646 40290 49698
rect 40290 49646 40292 49698
rect 40236 49644 40292 49646
rect 40124 48972 40180 49028
rect 40908 49868 40964 49924
rect 40684 49420 40740 49476
rect 40460 49026 40516 49028
rect 40460 48974 40462 49026
rect 40462 48974 40514 49026
rect 40514 48974 40516 49026
rect 40460 48972 40516 48974
rect 40236 48860 40292 48916
rect 41132 48914 41188 48916
rect 41132 48862 41134 48914
rect 41134 48862 41186 48914
rect 41186 48862 41188 48914
rect 41132 48860 41188 48862
rect 39788 48354 39844 48356
rect 39788 48302 39790 48354
rect 39790 48302 39842 48354
rect 39842 48302 39844 48354
rect 39788 48300 39844 48302
rect 40012 48636 40068 48692
rect 40348 48130 40404 48132
rect 40348 48078 40350 48130
rect 40350 48078 40402 48130
rect 40402 48078 40404 48130
rect 40348 48076 40404 48078
rect 39228 47964 39284 48020
rect 39004 47570 39060 47572
rect 39004 47518 39006 47570
rect 39006 47518 39058 47570
rect 39058 47518 39060 47570
rect 39004 47516 39060 47518
rect 41020 47740 41076 47796
rect 39676 47346 39732 47348
rect 39676 47294 39678 47346
rect 39678 47294 39730 47346
rect 39730 47294 39732 47346
rect 39676 47292 39732 47294
rect 39228 47068 39284 47124
rect 38780 46620 38836 46676
rect 40124 47068 40180 47124
rect 39676 46002 39732 46004
rect 39676 45950 39678 46002
rect 39678 45950 39730 46002
rect 39730 45950 39732 46002
rect 39676 45948 39732 45950
rect 39452 45500 39508 45556
rect 39788 45500 39844 45556
rect 38332 45276 38388 45332
rect 38892 45330 38948 45332
rect 38892 45278 38894 45330
rect 38894 45278 38946 45330
rect 38946 45278 38948 45330
rect 38892 45276 38948 45278
rect 39228 45052 39284 45108
rect 39004 44994 39060 44996
rect 39004 44942 39006 44994
rect 39006 44942 39058 44994
rect 39058 44942 39060 44994
rect 39004 44940 39060 44942
rect 38332 44828 38388 44884
rect 38556 44380 38612 44436
rect 38556 44156 38612 44212
rect 37436 40402 37492 40404
rect 37436 40350 37438 40402
rect 37438 40350 37490 40402
rect 37490 40350 37492 40402
rect 37436 40348 37492 40350
rect 37660 39788 37716 39844
rect 38220 41916 38276 41972
rect 38444 43484 38500 43540
rect 39004 44546 39060 44548
rect 39004 44494 39006 44546
rect 39006 44494 39058 44546
rect 39058 44494 39060 44546
rect 39004 44492 39060 44494
rect 40572 47292 40628 47348
rect 40348 45948 40404 46004
rect 40012 45052 40068 45108
rect 39228 43708 39284 43764
rect 39452 44380 39508 44436
rect 39676 44322 39732 44324
rect 39676 44270 39678 44322
rect 39678 44270 39730 44322
rect 39730 44270 39732 44322
rect 39676 44268 39732 44270
rect 40124 43596 40180 43652
rect 40460 43708 40516 43764
rect 39340 43372 39396 43428
rect 38892 42700 38948 42756
rect 39116 43148 39172 43204
rect 38444 42476 38500 42532
rect 39004 42530 39060 42532
rect 39004 42478 39006 42530
rect 39006 42478 39058 42530
rect 39058 42478 39060 42530
rect 39004 42476 39060 42478
rect 38892 42140 38948 42196
rect 38668 41970 38724 41972
rect 38668 41918 38670 41970
rect 38670 41918 38722 41970
rect 38722 41918 38724 41970
rect 38668 41916 38724 41918
rect 39564 42700 39620 42756
rect 39228 41916 39284 41972
rect 38668 41244 38724 41300
rect 39004 41298 39060 41300
rect 39004 41246 39006 41298
rect 39006 41246 39058 41298
rect 39058 41246 39060 41298
rect 39004 41244 39060 41246
rect 39340 41244 39396 41300
rect 39900 43260 39956 43316
rect 39788 41746 39844 41748
rect 39788 41694 39790 41746
rect 39790 41694 39842 41746
rect 39842 41694 39844 41746
rect 39788 41692 39844 41694
rect 41132 45724 41188 45780
rect 41580 52946 41636 52948
rect 41580 52894 41582 52946
rect 41582 52894 41634 52946
rect 41634 52894 41636 52946
rect 41580 52892 41636 52894
rect 41580 52668 41636 52724
rect 41244 45276 41300 45332
rect 41356 52108 41412 52164
rect 40796 43650 40852 43652
rect 40796 43598 40798 43650
rect 40798 43598 40850 43650
rect 40850 43598 40852 43650
rect 40796 43596 40852 43598
rect 40572 43484 40628 43540
rect 40124 42754 40180 42756
rect 40124 42702 40126 42754
rect 40126 42702 40178 42754
rect 40178 42702 40180 42754
rect 40124 42700 40180 42702
rect 40684 42082 40740 42084
rect 40684 42030 40686 42082
rect 40686 42030 40738 42082
rect 40738 42030 40740 42082
rect 40684 42028 40740 42030
rect 40460 41970 40516 41972
rect 40460 41918 40462 41970
rect 40462 41918 40514 41970
rect 40514 41918 40516 41970
rect 40460 41916 40516 41918
rect 39676 41244 39732 41300
rect 40012 41020 40068 41076
rect 39900 40962 39956 40964
rect 39900 40910 39902 40962
rect 39902 40910 39954 40962
rect 39954 40910 39956 40962
rect 39900 40908 39956 40910
rect 40572 41692 40628 41748
rect 40348 41020 40404 41076
rect 40460 40908 40516 40964
rect 40684 40908 40740 40964
rect 40012 40626 40068 40628
rect 40012 40574 40014 40626
rect 40014 40574 40066 40626
rect 40066 40574 40068 40626
rect 40012 40572 40068 40574
rect 40796 40626 40852 40628
rect 40796 40574 40798 40626
rect 40798 40574 40850 40626
rect 40850 40574 40852 40626
rect 40796 40572 40852 40574
rect 37884 39788 37940 39844
rect 40908 40236 40964 40292
rect 40796 39788 40852 39844
rect 37772 39116 37828 39172
rect 38108 39116 38164 39172
rect 39340 39618 39396 39620
rect 39340 39566 39342 39618
rect 39342 39566 39394 39618
rect 39394 39566 39396 39618
rect 39340 39564 39396 39566
rect 40572 39618 40628 39620
rect 40572 39566 40574 39618
rect 40574 39566 40626 39618
rect 40626 39566 40628 39618
rect 40572 39564 40628 39566
rect 37772 38668 37828 38724
rect 37548 37548 37604 37604
rect 36316 35420 36372 35476
rect 36764 34412 36820 34468
rect 36316 33292 36372 33348
rect 36764 33964 36820 34020
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 36204 31106 36260 31108
rect 36204 31054 36206 31106
rect 36206 31054 36258 31106
rect 36258 31054 36260 31106
rect 36204 31052 36260 31054
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 33740 30322 33796 30324
rect 33740 30270 33742 30322
rect 33742 30270 33794 30322
rect 33794 30270 33796 30322
rect 33740 30268 33796 30270
rect 35308 30268 35364 30324
rect 33516 29426 33572 29428
rect 33516 29374 33518 29426
rect 33518 29374 33570 29426
rect 33570 29374 33572 29426
rect 33516 29372 33572 29374
rect 34524 29820 34580 29876
rect 35084 29820 35140 29876
rect 36204 30268 36260 30324
rect 35980 29820 36036 29876
rect 33964 29372 34020 29428
rect 35532 29708 35588 29764
rect 33516 29036 33572 29092
rect 33404 28588 33460 28644
rect 33292 27020 33348 27076
rect 33628 28364 33684 28420
rect 33740 27916 33796 27972
rect 34636 28812 34692 28868
rect 34076 27916 34132 27972
rect 33964 27692 34020 27748
rect 34076 27580 34132 27636
rect 35420 29372 35476 29428
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35084 28700 35140 28756
rect 35756 28812 35812 28868
rect 35868 28700 35924 28756
rect 35644 28588 35700 28644
rect 35084 28530 35140 28532
rect 35084 28478 35086 28530
rect 35086 28478 35138 28530
rect 35138 28478 35140 28530
rect 35084 28476 35140 28478
rect 34972 28418 35028 28420
rect 34972 28366 34974 28418
rect 34974 28366 35026 28418
rect 35026 28366 35028 28418
rect 34972 28364 35028 28366
rect 35196 27692 35252 27748
rect 34748 27634 34804 27636
rect 34748 27582 34750 27634
rect 34750 27582 34802 27634
rect 34802 27582 34804 27634
rect 34748 27580 34804 27582
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 33180 26236 33236 26292
rect 33516 26124 33572 26180
rect 32956 25564 33012 25620
rect 33292 25788 33348 25844
rect 31052 23660 31108 23716
rect 30716 22876 30772 22932
rect 30828 23548 30884 23604
rect 30716 21980 30772 22036
rect 31612 23548 31668 23604
rect 32172 24050 32228 24052
rect 32172 23998 32174 24050
rect 32174 23998 32226 24050
rect 32226 23998 32228 24050
rect 32172 23996 32228 23998
rect 31836 23660 31892 23716
rect 31724 23212 31780 23268
rect 31724 22764 31780 22820
rect 31612 22652 31668 22708
rect 30604 21196 30660 21252
rect 31388 22092 31444 22148
rect 30940 21698 30996 21700
rect 30940 21646 30942 21698
rect 30942 21646 30994 21698
rect 30994 21646 30996 21698
rect 30940 21644 30996 21646
rect 31724 21980 31780 22036
rect 30716 20802 30772 20804
rect 30716 20750 30718 20802
rect 30718 20750 30770 20802
rect 30770 20750 30772 20802
rect 30716 20748 30772 20750
rect 30716 20018 30772 20020
rect 30716 19966 30718 20018
rect 30718 19966 30770 20018
rect 30770 19966 30772 20018
rect 30716 19964 30772 19966
rect 30380 19628 30436 19684
rect 30156 19068 30212 19124
rect 30604 19068 30660 19124
rect 30044 15596 30100 15652
rect 29148 15314 29204 15316
rect 29148 15262 29150 15314
rect 29150 15262 29202 15314
rect 29202 15262 29204 15314
rect 29148 15260 29204 15262
rect 29596 15538 29652 15540
rect 29596 15486 29598 15538
rect 29598 15486 29650 15538
rect 29650 15486 29652 15538
rect 29596 15484 29652 15486
rect 30380 17500 30436 17556
rect 30492 18060 30548 18116
rect 30828 19122 30884 19124
rect 30828 19070 30830 19122
rect 30830 19070 30882 19122
rect 30882 19070 30884 19122
rect 30828 19068 30884 19070
rect 30828 17890 30884 17892
rect 30828 17838 30830 17890
rect 30830 17838 30882 17890
rect 30882 17838 30884 17890
rect 30828 17836 30884 17838
rect 30828 17276 30884 17332
rect 30828 16882 30884 16884
rect 30828 16830 30830 16882
rect 30830 16830 30882 16882
rect 30882 16830 30884 16882
rect 30828 16828 30884 16830
rect 30380 15596 30436 15652
rect 29596 15036 29652 15092
rect 30380 15260 30436 15316
rect 29484 14530 29540 14532
rect 29484 14478 29486 14530
rect 29486 14478 29538 14530
rect 29538 14478 29540 14530
rect 29484 14476 29540 14478
rect 29260 13580 29316 13636
rect 29708 13468 29764 13524
rect 29596 13074 29652 13076
rect 29596 13022 29598 13074
rect 29598 13022 29650 13074
rect 29650 13022 29652 13074
rect 29596 13020 29652 13022
rect 29820 14252 29876 14308
rect 30268 14306 30324 14308
rect 30268 14254 30270 14306
rect 30270 14254 30322 14306
rect 30322 14254 30324 14306
rect 30268 14252 30324 14254
rect 30268 13746 30324 13748
rect 30268 13694 30270 13746
rect 30270 13694 30322 13746
rect 30322 13694 30324 13746
rect 30268 13692 30324 13694
rect 29708 12908 29764 12964
rect 29260 12684 29316 12740
rect 29708 12738 29764 12740
rect 29708 12686 29710 12738
rect 29710 12686 29762 12738
rect 29762 12686 29764 12738
rect 29708 12684 29764 12686
rect 31052 20914 31108 20916
rect 31052 20862 31054 20914
rect 31054 20862 31106 20914
rect 31106 20862 31108 20914
rect 31052 20860 31108 20862
rect 31276 20914 31332 20916
rect 31276 20862 31278 20914
rect 31278 20862 31330 20914
rect 31330 20862 31332 20914
rect 31276 20860 31332 20862
rect 32732 24668 32788 24724
rect 32956 24556 33012 24612
rect 32172 22876 32228 22932
rect 32172 22316 32228 22372
rect 31948 21698 32004 21700
rect 31948 21646 31950 21698
rect 31950 21646 32002 21698
rect 32002 21646 32004 21698
rect 31948 21644 32004 21646
rect 31164 20524 31220 20580
rect 30940 14812 30996 14868
rect 31836 20578 31892 20580
rect 31836 20526 31838 20578
rect 31838 20526 31890 20578
rect 31890 20526 31892 20578
rect 31836 20524 31892 20526
rect 31052 19292 31108 19348
rect 31164 17836 31220 17892
rect 31276 19180 31332 19236
rect 31388 19122 31444 19124
rect 31388 19070 31390 19122
rect 31390 19070 31442 19122
rect 31442 19070 31444 19122
rect 31388 19068 31444 19070
rect 31836 19292 31892 19348
rect 31948 19180 32004 19236
rect 32620 21196 32676 21252
rect 32172 20972 32228 21028
rect 32620 20972 32676 21028
rect 31724 18956 31780 19012
rect 31612 18562 31668 18564
rect 31612 18510 31614 18562
rect 31614 18510 31666 18562
rect 31666 18510 31668 18562
rect 31612 18508 31668 18510
rect 31500 17724 31556 17780
rect 32396 19346 32452 19348
rect 32396 19294 32398 19346
rect 32398 19294 32450 19346
rect 32450 19294 32452 19346
rect 32396 19292 32452 19294
rect 31948 18396 32004 18452
rect 31836 18284 31892 18340
rect 31164 17164 31220 17220
rect 31276 17106 31332 17108
rect 31276 17054 31278 17106
rect 31278 17054 31330 17106
rect 31330 17054 31332 17106
rect 31276 17052 31332 17054
rect 31612 17052 31668 17108
rect 32396 18338 32452 18340
rect 32396 18286 32398 18338
rect 32398 18286 32450 18338
rect 32450 18286 32452 18338
rect 32396 18284 32452 18286
rect 32732 19292 32788 19348
rect 32844 20972 32900 21028
rect 33068 23212 33124 23268
rect 33180 22428 33236 22484
rect 33852 25676 33908 25732
rect 33516 25340 33572 25396
rect 33404 24556 33460 24612
rect 33404 22764 33460 22820
rect 33740 25004 33796 25060
rect 33628 24722 33684 24724
rect 33628 24670 33630 24722
rect 33630 24670 33682 24722
rect 33682 24670 33684 24722
rect 33628 24668 33684 24670
rect 34636 26962 34692 26964
rect 34636 26910 34638 26962
rect 34638 26910 34690 26962
rect 34690 26910 34692 26962
rect 34636 26908 34692 26910
rect 34524 26572 34580 26628
rect 34860 27074 34916 27076
rect 34860 27022 34862 27074
rect 34862 27022 34914 27074
rect 34914 27022 34916 27074
rect 34860 27020 34916 27022
rect 34972 26908 35028 26964
rect 33964 25506 34020 25508
rect 33964 25454 33966 25506
rect 33966 25454 34018 25506
rect 34018 25454 34020 25506
rect 33964 25452 34020 25454
rect 34300 25394 34356 25396
rect 34300 25342 34302 25394
rect 34302 25342 34354 25394
rect 34354 25342 34356 25394
rect 34300 25340 34356 25342
rect 34076 24556 34132 24612
rect 34188 24332 34244 24388
rect 34300 24444 34356 24500
rect 33964 24108 34020 24164
rect 33964 23772 34020 23828
rect 34188 23548 34244 23604
rect 33292 22204 33348 22260
rect 33180 21196 33236 21252
rect 33068 18508 33124 18564
rect 32508 17836 32564 17892
rect 32620 18396 32676 18452
rect 32396 17666 32452 17668
rect 32396 17614 32398 17666
rect 32398 17614 32450 17666
rect 32450 17614 32452 17666
rect 32396 17612 32452 17614
rect 31948 17276 32004 17332
rect 32060 16882 32116 16884
rect 32060 16830 32062 16882
rect 32062 16830 32114 16882
rect 32114 16830 32116 16882
rect 32060 16828 32116 16830
rect 31948 16044 32004 16100
rect 32396 17052 32452 17108
rect 31948 15260 32004 15316
rect 31836 15148 31892 15204
rect 30492 14252 30548 14308
rect 30380 12124 30436 12180
rect 29932 12066 29988 12068
rect 29932 12014 29934 12066
rect 29934 12014 29986 12066
rect 29986 12014 29988 12066
rect 29932 12012 29988 12014
rect 30492 12066 30548 12068
rect 30492 12014 30494 12066
rect 30494 12014 30546 12066
rect 30546 12014 30548 12066
rect 30492 12012 30548 12014
rect 27468 8204 27524 8260
rect 27356 8092 27412 8148
rect 27804 8146 27860 8148
rect 27804 8094 27806 8146
rect 27806 8094 27858 8146
rect 27858 8094 27860 8146
rect 27804 8092 27860 8094
rect 27468 7362 27524 7364
rect 27468 7310 27470 7362
rect 27470 7310 27522 7362
rect 27522 7310 27524 7362
rect 27468 7308 27524 7310
rect 27468 6690 27524 6692
rect 27468 6638 27470 6690
rect 27470 6638 27522 6690
rect 27522 6638 27524 6690
rect 27468 6636 27524 6638
rect 26348 4450 26404 4452
rect 26348 4398 26350 4450
rect 26350 4398 26402 4450
rect 26402 4398 26404 4450
rect 26348 4396 26404 4398
rect 26684 4338 26740 4340
rect 26684 4286 26686 4338
rect 26686 4286 26738 4338
rect 26738 4286 26740 4338
rect 26684 4284 26740 4286
rect 25564 4172 25620 4228
rect 26796 3554 26852 3556
rect 26796 3502 26798 3554
rect 26798 3502 26850 3554
rect 26850 3502 26852 3554
rect 26796 3500 26852 3502
rect 27356 3500 27412 3556
rect 23884 2716 23940 2772
rect 28028 9100 28084 9156
rect 29932 10668 29988 10724
rect 30380 11228 30436 11284
rect 29484 9826 29540 9828
rect 29484 9774 29486 9826
rect 29486 9774 29538 9826
rect 29538 9774 29540 9826
rect 29484 9772 29540 9774
rect 29148 9660 29204 9716
rect 29820 8428 29876 8484
rect 28476 8092 28532 8148
rect 28476 7756 28532 7812
rect 28476 7586 28532 7588
rect 28476 7534 28478 7586
rect 28478 7534 28530 7586
rect 28530 7534 28532 7586
rect 28476 7532 28532 7534
rect 28140 7474 28196 7476
rect 28140 7422 28142 7474
rect 28142 7422 28194 7474
rect 28194 7422 28196 7474
rect 28140 7420 28196 7422
rect 28700 7420 28756 7476
rect 28028 6690 28084 6692
rect 28028 6638 28030 6690
rect 28030 6638 28082 6690
rect 28082 6638 28084 6690
rect 28028 6636 28084 6638
rect 28140 6300 28196 6356
rect 28252 6188 28308 6244
rect 28364 7308 28420 7364
rect 29036 7474 29092 7476
rect 29036 7422 29038 7474
rect 29038 7422 29090 7474
rect 29090 7422 29092 7474
rect 29036 7420 29092 7422
rect 30156 9042 30212 9044
rect 30156 8990 30158 9042
rect 30158 8990 30210 9042
rect 30210 8990 30212 9042
rect 30156 8988 30212 8990
rect 30044 7532 30100 7588
rect 29820 7420 29876 7476
rect 29036 7084 29092 7140
rect 29484 6300 29540 6356
rect 29820 6188 29876 6244
rect 28364 5180 28420 5236
rect 28588 4226 28644 4228
rect 28588 4174 28590 4226
rect 28590 4174 28642 4226
rect 28642 4174 28644 4226
rect 28588 4172 28644 4174
rect 29372 4508 29428 4564
rect 29820 4508 29876 4564
rect 27916 3052 27972 3108
rect 28476 3554 28532 3556
rect 28476 3502 28478 3554
rect 28478 3502 28530 3554
rect 28530 3502 28532 3554
rect 28476 3500 28532 3502
rect 31052 14418 31108 14420
rect 31052 14366 31054 14418
rect 31054 14366 31106 14418
rect 31106 14366 31108 14418
rect 31052 14364 31108 14366
rect 32060 14588 32116 14644
rect 31948 14530 32004 14532
rect 31948 14478 31950 14530
rect 31950 14478 32002 14530
rect 32002 14478 32004 14530
rect 31948 14476 32004 14478
rect 30940 12738 30996 12740
rect 30940 12686 30942 12738
rect 30942 12686 30994 12738
rect 30994 12686 30996 12738
rect 30940 12684 30996 12686
rect 31164 12460 31220 12516
rect 31500 13522 31556 13524
rect 31500 13470 31502 13522
rect 31502 13470 31554 13522
rect 31554 13470 31556 13522
rect 31500 13468 31556 13470
rect 31836 13356 31892 13412
rect 31500 12850 31556 12852
rect 31500 12798 31502 12850
rect 31502 12798 31554 12850
rect 31554 12798 31556 12850
rect 31500 12796 31556 12798
rect 31276 12178 31332 12180
rect 31276 12126 31278 12178
rect 31278 12126 31330 12178
rect 31330 12126 31332 12178
rect 31276 12124 31332 12126
rect 31052 12012 31108 12068
rect 30940 11900 30996 11956
rect 30604 11394 30660 11396
rect 30604 11342 30606 11394
rect 30606 11342 30658 11394
rect 30658 11342 30660 11394
rect 30604 11340 30660 11342
rect 30492 11116 30548 11172
rect 30492 10722 30548 10724
rect 30492 10670 30494 10722
rect 30494 10670 30546 10722
rect 30546 10670 30548 10722
rect 30492 10668 30548 10670
rect 30604 9660 30660 9716
rect 30604 8428 30660 8484
rect 30492 8370 30548 8372
rect 30492 8318 30494 8370
rect 30494 8318 30546 8370
rect 30546 8318 30548 8370
rect 30492 8316 30548 8318
rect 31052 11394 31108 11396
rect 31052 11342 31054 11394
rect 31054 11342 31106 11394
rect 31106 11342 31108 11394
rect 31052 11340 31108 11342
rect 31276 11170 31332 11172
rect 31276 11118 31278 11170
rect 31278 11118 31330 11170
rect 31330 11118 31332 11170
rect 31276 11116 31332 11118
rect 31164 10610 31220 10612
rect 31164 10558 31166 10610
rect 31166 10558 31218 10610
rect 31218 10558 31220 10610
rect 31164 10556 31220 10558
rect 32620 16940 32676 16996
rect 32508 16604 32564 16660
rect 32956 17836 33012 17892
rect 32732 15874 32788 15876
rect 32732 15822 32734 15874
rect 32734 15822 32786 15874
rect 32786 15822 32788 15874
rect 32732 15820 32788 15822
rect 32620 15484 32676 15540
rect 32284 15202 32340 15204
rect 32284 15150 32286 15202
rect 32286 15150 32338 15202
rect 32338 15150 32340 15202
rect 32284 15148 32340 15150
rect 32844 15148 32900 15204
rect 32732 14588 32788 14644
rect 32732 14252 32788 14308
rect 32396 13356 32452 13412
rect 32620 12850 32676 12852
rect 32620 12798 32622 12850
rect 32622 12798 32674 12850
rect 32674 12798 32676 12850
rect 32620 12796 32676 12798
rect 31836 12178 31892 12180
rect 31836 12126 31838 12178
rect 31838 12126 31890 12178
rect 31890 12126 31892 12178
rect 31836 12124 31892 12126
rect 31724 11116 31780 11172
rect 31836 11676 31892 11732
rect 31164 8370 31220 8372
rect 31164 8318 31166 8370
rect 31166 8318 31218 8370
rect 31218 8318 31220 8370
rect 31164 8316 31220 8318
rect 30940 7756 30996 7812
rect 30940 7362 30996 7364
rect 30940 7310 30942 7362
rect 30942 7310 30994 7362
rect 30994 7310 30996 7362
rect 30940 7308 30996 7310
rect 32060 11564 32116 11620
rect 31948 11394 32004 11396
rect 31948 11342 31950 11394
rect 31950 11342 32002 11394
rect 32002 11342 32004 11394
rect 31948 11340 32004 11342
rect 32172 11282 32228 11284
rect 32172 11230 32174 11282
rect 32174 11230 32226 11282
rect 32226 11230 32228 11282
rect 32172 11228 32228 11230
rect 32060 10556 32116 10612
rect 31836 8764 31892 8820
rect 32172 8988 32228 9044
rect 32508 12178 32564 12180
rect 32508 12126 32510 12178
rect 32510 12126 32562 12178
rect 32562 12126 32564 12178
rect 32508 12124 32564 12126
rect 32620 11900 32676 11956
rect 32508 11788 32564 11844
rect 32396 11228 32452 11284
rect 32508 9212 32564 9268
rect 32284 8316 32340 8372
rect 32172 7756 32228 7812
rect 31276 7196 31332 7252
rect 30828 6690 30884 6692
rect 30828 6638 30830 6690
rect 30830 6638 30882 6690
rect 30882 6638 30884 6690
rect 30828 6636 30884 6638
rect 30716 6578 30772 6580
rect 30716 6526 30718 6578
rect 30718 6526 30770 6578
rect 30770 6526 30772 6578
rect 30716 6524 30772 6526
rect 31164 6076 31220 6132
rect 30604 4450 30660 4452
rect 30604 4398 30606 4450
rect 30606 4398 30658 4450
rect 30658 4398 30660 4450
rect 30604 4396 30660 4398
rect 30380 3500 30436 3556
rect 31164 5234 31220 5236
rect 31164 5182 31166 5234
rect 31166 5182 31218 5234
rect 31218 5182 31220 5234
rect 31164 5180 31220 5182
rect 31388 6524 31444 6580
rect 31724 7308 31780 7364
rect 31612 6690 31668 6692
rect 31612 6638 31614 6690
rect 31614 6638 31666 6690
rect 31666 6638 31668 6690
rect 31612 6636 31668 6638
rect 31836 6636 31892 6692
rect 32172 5852 32228 5908
rect 32396 6466 32452 6468
rect 32396 6414 32398 6466
rect 32398 6414 32450 6466
rect 32450 6414 32452 6466
rect 32396 6412 32452 6414
rect 31724 5740 31780 5796
rect 31500 5346 31556 5348
rect 31500 5294 31502 5346
rect 31502 5294 31554 5346
rect 31554 5294 31556 5346
rect 31500 5292 31556 5294
rect 32396 5292 32452 5348
rect 32620 6018 32676 6020
rect 32620 5966 32622 6018
rect 32622 5966 32674 6018
rect 32674 5966 32676 6018
rect 32620 5964 32676 5966
rect 32396 4620 32452 4676
rect 31836 4338 31892 4340
rect 31836 4286 31838 4338
rect 31838 4286 31890 4338
rect 31890 4286 31892 4338
rect 31836 4284 31892 4286
rect 30940 2940 30996 2996
rect 32956 12962 33012 12964
rect 32956 12910 32958 12962
rect 32958 12910 33010 12962
rect 33010 12910 33012 12962
rect 32956 12908 33012 12910
rect 33516 22316 33572 22372
rect 33516 22092 33572 22148
rect 33740 22988 33796 23044
rect 33740 21756 33796 21812
rect 33628 21308 33684 21364
rect 33404 18620 33460 18676
rect 33516 19852 33572 19908
rect 33628 19234 33684 19236
rect 33628 19182 33630 19234
rect 33630 19182 33682 19234
rect 33682 19182 33684 19234
rect 33628 19180 33684 19182
rect 33516 19122 33572 19124
rect 33516 19070 33518 19122
rect 33518 19070 33570 19122
rect 33570 19070 33572 19122
rect 33516 19068 33572 19070
rect 33292 17276 33348 17332
rect 33404 17052 33460 17108
rect 33180 16828 33236 16884
rect 34076 22258 34132 22260
rect 34076 22206 34078 22258
rect 34078 22206 34130 22258
rect 34130 22206 34132 22258
rect 34076 22204 34132 22206
rect 34524 25116 34580 25172
rect 34412 22540 34468 22596
rect 34524 24108 34580 24164
rect 34412 22204 34468 22260
rect 35420 26514 35476 26516
rect 35420 26462 35422 26514
rect 35422 26462 35474 26514
rect 35474 26462 35476 26514
rect 35420 26460 35476 26462
rect 35756 27580 35812 27636
rect 35756 27244 35812 27300
rect 35644 27132 35700 27188
rect 35644 26796 35700 26852
rect 36092 28754 36148 28756
rect 36092 28702 36094 28754
rect 36094 28702 36146 28754
rect 36146 28702 36148 28754
rect 36092 28700 36148 28702
rect 35980 27858 36036 27860
rect 35980 27806 35982 27858
rect 35982 27806 36034 27858
rect 36034 27806 36036 27858
rect 35980 27804 36036 27806
rect 35980 27132 36036 27188
rect 35644 26236 35700 26292
rect 35420 26124 35476 26180
rect 35532 26012 35588 26068
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35084 25676 35140 25732
rect 35420 25506 35476 25508
rect 35420 25454 35422 25506
rect 35422 25454 35474 25506
rect 35474 25454 35476 25506
rect 35420 25452 35476 25454
rect 34972 24444 35028 24500
rect 34972 23884 35028 23940
rect 35196 25282 35252 25284
rect 35196 25230 35198 25282
rect 35198 25230 35250 25282
rect 35250 25230 35252 25282
rect 35196 25228 35252 25230
rect 35420 24498 35476 24500
rect 35420 24446 35422 24498
rect 35422 24446 35474 24498
rect 35474 24446 35476 24498
rect 35420 24444 35476 24446
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 34860 23714 34916 23716
rect 34860 23662 34862 23714
rect 34862 23662 34914 23714
rect 34914 23662 34916 23714
rect 34860 23660 34916 23662
rect 34636 22988 34692 23044
rect 34748 22652 34804 22708
rect 35420 23548 35476 23604
rect 35644 25564 35700 25620
rect 35532 23436 35588 23492
rect 35868 26460 35924 26516
rect 35980 26402 36036 26404
rect 35980 26350 35982 26402
rect 35982 26350 36034 26402
rect 36034 26350 36036 26402
rect 35980 26348 36036 26350
rect 35868 25730 35924 25732
rect 35868 25678 35870 25730
rect 35870 25678 35922 25730
rect 35922 25678 35924 25730
rect 35868 25676 35924 25678
rect 35868 25452 35924 25508
rect 35980 24668 36036 24724
rect 35980 24332 36036 24388
rect 35980 23826 36036 23828
rect 35980 23774 35982 23826
rect 35982 23774 36034 23826
rect 36034 23774 36036 23826
rect 35980 23772 36036 23774
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35084 22540 35140 22596
rect 33964 21362 34020 21364
rect 33964 21310 33966 21362
rect 33966 21310 34018 21362
rect 34018 21310 34020 21362
rect 33964 21308 34020 21310
rect 33964 20242 34020 20244
rect 33964 20190 33966 20242
rect 33966 20190 34018 20242
rect 34018 20190 34020 20242
rect 33964 20188 34020 20190
rect 34300 20300 34356 20356
rect 34188 19516 34244 19572
rect 34300 19404 34356 19460
rect 34076 19180 34132 19236
rect 35420 22316 35476 22372
rect 36428 31836 36484 31892
rect 37996 37548 38052 37604
rect 38556 38610 38612 38612
rect 38556 38558 38558 38610
rect 38558 38558 38610 38610
rect 38610 38558 38612 38610
rect 38556 38556 38612 38558
rect 40012 38834 40068 38836
rect 40012 38782 40014 38834
rect 40014 38782 40066 38834
rect 40066 38782 40068 38834
rect 40012 38780 40068 38782
rect 39564 38722 39620 38724
rect 39564 38670 39566 38722
rect 39566 38670 39618 38722
rect 39618 38670 39620 38722
rect 39564 38668 39620 38670
rect 38332 37548 38388 37604
rect 39340 38332 39396 38388
rect 38668 36594 38724 36596
rect 38668 36542 38670 36594
rect 38670 36542 38722 36594
rect 38722 36542 38724 36594
rect 38668 36540 38724 36542
rect 38444 36204 38500 36260
rect 38668 36204 38724 36260
rect 38444 35980 38500 36036
rect 39004 35980 39060 36036
rect 39228 36316 39284 36372
rect 37100 34412 37156 34468
rect 37212 34300 37268 34356
rect 39004 34690 39060 34692
rect 39004 34638 39006 34690
rect 39006 34638 39058 34690
rect 39058 34638 39060 34690
rect 39004 34636 39060 34638
rect 37772 34300 37828 34356
rect 40460 38722 40516 38724
rect 40460 38670 40462 38722
rect 40462 38670 40514 38722
rect 40514 38670 40516 38722
rect 40460 38668 40516 38670
rect 39452 38220 39508 38276
rect 41132 36876 41188 36932
rect 40124 36482 40180 36484
rect 40124 36430 40126 36482
rect 40126 36430 40178 36482
rect 40178 36430 40180 36482
rect 40124 36428 40180 36430
rect 41132 35980 41188 36036
rect 39340 34188 39396 34244
rect 40460 34636 40516 34692
rect 38220 34018 38276 34020
rect 38220 33966 38222 34018
rect 38222 33966 38274 34018
rect 38274 33966 38276 34018
rect 38220 33964 38276 33966
rect 37436 33292 37492 33348
rect 37660 33346 37716 33348
rect 37660 33294 37662 33346
rect 37662 33294 37714 33346
rect 37714 33294 37716 33346
rect 37660 33292 37716 33294
rect 37548 32620 37604 32676
rect 36764 31276 36820 31332
rect 36428 29708 36484 29764
rect 37436 31052 37492 31108
rect 39452 33292 39508 33348
rect 41020 33292 41076 33348
rect 37996 32674 38052 32676
rect 37996 32622 37998 32674
rect 37998 32622 38050 32674
rect 38050 32622 38052 32674
rect 37996 32620 38052 32622
rect 38444 31666 38500 31668
rect 38444 31614 38446 31666
rect 38446 31614 38498 31666
rect 38498 31614 38500 31666
rect 38444 31612 38500 31614
rect 40348 31836 40404 31892
rect 38668 31612 38724 31668
rect 37884 31276 37940 31332
rect 40124 31500 40180 31556
rect 37660 30380 37716 30436
rect 36652 29820 36708 29876
rect 36540 29538 36596 29540
rect 36540 29486 36542 29538
rect 36542 29486 36594 29538
rect 36594 29486 36596 29538
rect 36540 29484 36596 29486
rect 36428 29426 36484 29428
rect 36428 29374 36430 29426
rect 36430 29374 36482 29426
rect 36482 29374 36484 29426
rect 36428 29372 36484 29374
rect 37436 29708 37492 29764
rect 38108 30434 38164 30436
rect 38108 30382 38110 30434
rect 38110 30382 38162 30434
rect 38162 30382 38164 30434
rect 38108 30380 38164 30382
rect 37884 29484 37940 29540
rect 36652 29372 36708 29428
rect 37324 29372 37380 29428
rect 36316 26850 36372 26852
rect 36316 26798 36318 26850
rect 36318 26798 36370 26850
rect 36370 26798 36372 26850
rect 36316 26796 36372 26798
rect 37772 29426 37828 29428
rect 37772 29374 37774 29426
rect 37774 29374 37826 29426
rect 37826 29374 37828 29426
rect 37772 29372 37828 29374
rect 37548 28588 37604 28644
rect 38332 29538 38388 29540
rect 38332 29486 38334 29538
rect 38334 29486 38386 29538
rect 38386 29486 38388 29538
rect 38332 29484 38388 29486
rect 38668 29538 38724 29540
rect 38668 29486 38670 29538
rect 38670 29486 38722 29538
rect 38722 29486 38724 29538
rect 38668 29484 38724 29486
rect 39116 29538 39172 29540
rect 39116 29486 39118 29538
rect 39118 29486 39170 29538
rect 39170 29486 39172 29538
rect 39116 29484 39172 29486
rect 37436 28418 37492 28420
rect 37436 28366 37438 28418
rect 37438 28366 37490 28418
rect 37490 28366 37492 28418
rect 37436 28364 37492 28366
rect 36540 27746 36596 27748
rect 36540 27694 36542 27746
rect 36542 27694 36594 27746
rect 36594 27694 36596 27746
rect 36540 27692 36596 27694
rect 36764 27468 36820 27524
rect 37548 27580 37604 27636
rect 36988 26908 37044 26964
rect 37100 27356 37156 27412
rect 36876 26460 36932 26516
rect 36764 26348 36820 26404
rect 36428 26012 36484 26068
rect 36540 25788 36596 25844
rect 37772 28140 37828 28196
rect 37772 27580 37828 27636
rect 38220 29148 38276 29204
rect 38220 28642 38276 28644
rect 38220 28590 38222 28642
rect 38222 28590 38274 28642
rect 38274 28590 38276 28642
rect 38220 28588 38276 28590
rect 38780 28700 38836 28756
rect 38444 27970 38500 27972
rect 38444 27918 38446 27970
rect 38446 27918 38498 27970
rect 38498 27918 38500 27970
rect 38444 27916 38500 27918
rect 37884 27356 37940 27412
rect 37996 27074 38052 27076
rect 37996 27022 37998 27074
rect 37998 27022 38050 27074
rect 38050 27022 38052 27074
rect 37996 27020 38052 27022
rect 37660 26908 37716 26964
rect 37100 25900 37156 25956
rect 36876 25452 36932 25508
rect 36988 25676 37044 25732
rect 36316 25228 36372 25284
rect 36764 25228 36820 25284
rect 37100 25564 37156 25620
rect 36204 24780 36260 24836
rect 36764 24834 36820 24836
rect 36764 24782 36766 24834
rect 36766 24782 36818 24834
rect 36818 24782 36820 24834
rect 36764 24780 36820 24782
rect 36316 24444 36372 24500
rect 36540 24332 36596 24388
rect 36540 23884 36596 23940
rect 36316 23826 36372 23828
rect 36316 23774 36318 23826
rect 36318 23774 36370 23826
rect 36370 23774 36372 23826
rect 36316 23772 36372 23774
rect 36540 23660 36596 23716
rect 36652 23548 36708 23604
rect 36764 24556 36820 24612
rect 36764 23212 36820 23268
rect 35868 23100 35924 23156
rect 36540 23100 36596 23156
rect 35756 23042 35812 23044
rect 35756 22990 35758 23042
rect 35758 22990 35810 23042
rect 35810 22990 35812 23042
rect 35756 22988 35812 22990
rect 35756 22540 35812 22596
rect 36092 22652 36148 22708
rect 36428 22652 36484 22708
rect 34636 20412 34692 20468
rect 34524 20300 34580 20356
rect 34972 20188 35028 20244
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35532 20860 35588 20916
rect 33964 18338 34020 18340
rect 33964 18286 33966 18338
rect 33966 18286 34018 18338
rect 34018 18286 34020 18338
rect 33964 18284 34020 18286
rect 34412 17666 34468 17668
rect 34412 17614 34414 17666
rect 34414 17614 34466 17666
rect 34466 17614 34468 17666
rect 34412 17612 34468 17614
rect 33740 17554 33796 17556
rect 33740 17502 33742 17554
rect 33742 17502 33794 17554
rect 33794 17502 33796 17554
rect 33740 17500 33796 17502
rect 33628 17442 33684 17444
rect 33628 17390 33630 17442
rect 33630 17390 33682 17442
rect 33682 17390 33684 17442
rect 33628 17388 33684 17390
rect 33628 16882 33684 16884
rect 33628 16830 33630 16882
rect 33630 16830 33682 16882
rect 33682 16830 33684 16882
rect 33628 16828 33684 16830
rect 33852 17388 33908 17444
rect 34524 17388 34580 17444
rect 34300 16492 34356 16548
rect 33740 15986 33796 15988
rect 33740 15934 33742 15986
rect 33742 15934 33794 15986
rect 33794 15934 33796 15986
rect 33740 15932 33796 15934
rect 33292 15148 33348 15204
rect 33180 14812 33236 14868
rect 33292 14306 33348 14308
rect 33292 14254 33294 14306
rect 33294 14254 33346 14306
rect 33346 14254 33348 14306
rect 33292 14252 33348 14254
rect 33180 12796 33236 12852
rect 33180 11170 33236 11172
rect 33180 11118 33182 11170
rect 33182 11118 33234 11170
rect 33234 11118 33236 11170
rect 33180 11116 33236 11118
rect 33180 10668 33236 10724
rect 33180 10050 33236 10052
rect 33180 9998 33182 10050
rect 33182 9998 33234 10050
rect 33234 9998 33236 10050
rect 33180 9996 33236 9998
rect 32844 9266 32900 9268
rect 32844 9214 32846 9266
rect 32846 9214 32898 9266
rect 32898 9214 32900 9266
rect 32844 9212 32900 9214
rect 33068 9602 33124 9604
rect 33068 9550 33070 9602
rect 33070 9550 33122 9602
rect 33122 9550 33124 9602
rect 33068 9548 33124 9550
rect 33740 15596 33796 15652
rect 33516 12066 33572 12068
rect 33516 12014 33518 12066
rect 33518 12014 33570 12066
rect 33570 12014 33572 12066
rect 33516 12012 33572 12014
rect 33628 11788 33684 11844
rect 33628 11394 33684 11396
rect 33628 11342 33630 11394
rect 33630 11342 33682 11394
rect 33682 11342 33684 11394
rect 33628 11340 33684 11342
rect 33964 12962 34020 12964
rect 33964 12910 33966 12962
rect 33966 12910 34018 12962
rect 34018 12910 34020 12962
rect 33964 12908 34020 12910
rect 33852 12850 33908 12852
rect 33852 12798 33854 12850
rect 33854 12798 33906 12850
rect 33906 12798 33908 12850
rect 33852 12796 33908 12798
rect 33964 11900 34020 11956
rect 34188 11900 34244 11956
rect 33740 10498 33796 10500
rect 33740 10446 33742 10498
rect 33742 10446 33794 10498
rect 33794 10446 33796 10498
rect 33740 10444 33796 10446
rect 33740 9996 33796 10052
rect 34524 15932 34580 15988
rect 34188 10556 34244 10612
rect 33964 10050 34020 10052
rect 33964 9998 33966 10050
rect 33966 9998 34018 10050
rect 34018 9998 34020 10050
rect 33964 9996 34020 9998
rect 33852 9212 33908 9268
rect 33292 8428 33348 8484
rect 33068 8146 33124 8148
rect 33068 8094 33070 8146
rect 33070 8094 33122 8146
rect 33122 8094 33124 8146
rect 33068 8092 33124 8094
rect 33180 8034 33236 8036
rect 33180 7982 33182 8034
rect 33182 7982 33234 8034
rect 33234 7982 33236 8034
rect 33180 7980 33236 7982
rect 32844 6690 32900 6692
rect 32844 6638 32846 6690
rect 32846 6638 32898 6690
rect 32898 6638 32900 6690
rect 32844 6636 32900 6638
rect 33068 6412 33124 6468
rect 33292 6636 33348 6692
rect 32956 4508 33012 4564
rect 33180 4620 33236 4676
rect 32732 2828 32788 2884
rect 28476 1596 28532 1652
rect 33628 8988 33684 9044
rect 34076 9660 34132 9716
rect 34412 10108 34468 10164
rect 34300 9100 34356 9156
rect 34412 9884 34468 9940
rect 34188 9042 34244 9044
rect 34188 8990 34190 9042
rect 34190 8990 34242 9042
rect 34242 8990 34244 9042
rect 34188 8988 34244 8990
rect 34412 8876 34468 8932
rect 33628 8428 33684 8484
rect 34188 8092 34244 8148
rect 34972 19404 35028 19460
rect 35420 20188 35476 20244
rect 35532 20076 35588 20132
rect 35980 21810 36036 21812
rect 35980 21758 35982 21810
rect 35982 21758 36034 21810
rect 36034 21758 36036 21810
rect 35980 21756 36036 21758
rect 36428 21308 36484 21364
rect 35868 20300 35924 20356
rect 35196 19852 35252 19908
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34860 19234 34916 19236
rect 34860 19182 34862 19234
rect 34862 19182 34914 19234
rect 34914 19182 34916 19234
rect 34860 19180 34916 19182
rect 34748 19122 34804 19124
rect 34748 19070 34750 19122
rect 34750 19070 34802 19122
rect 34802 19070 34804 19122
rect 34748 19068 34804 19070
rect 34860 18508 34916 18564
rect 34748 17836 34804 17892
rect 34748 17106 34804 17108
rect 34748 17054 34750 17106
rect 34750 17054 34802 17106
rect 34802 17054 34804 17106
rect 34748 17052 34804 17054
rect 35532 19010 35588 19012
rect 35532 18958 35534 19010
rect 35534 18958 35586 19010
rect 35586 18958 35588 19010
rect 35532 18956 35588 18958
rect 36204 20690 36260 20692
rect 36204 20638 36206 20690
rect 36206 20638 36258 20690
rect 36258 20638 36260 20690
rect 36204 20636 36260 20638
rect 36092 19852 36148 19908
rect 36204 20188 36260 20244
rect 36316 19404 36372 19460
rect 35308 18562 35364 18564
rect 35308 18510 35310 18562
rect 35310 18510 35362 18562
rect 35362 18510 35364 18562
rect 35308 18508 35364 18510
rect 35084 18396 35140 18452
rect 35756 18450 35812 18452
rect 35756 18398 35758 18450
rect 35758 18398 35810 18450
rect 35810 18398 35812 18450
rect 35756 18396 35812 18398
rect 36092 18562 36148 18564
rect 36092 18510 36094 18562
rect 36094 18510 36146 18562
rect 36146 18510 36148 18562
rect 36092 18508 36148 18510
rect 36316 18396 36372 18452
rect 35980 18284 36036 18340
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35980 17836 36036 17892
rect 34972 17052 35028 17108
rect 35084 17276 35140 17332
rect 34972 16882 35028 16884
rect 34972 16830 34974 16882
rect 34974 16830 35026 16882
rect 35026 16830 35028 16882
rect 34972 16828 35028 16830
rect 34860 16604 34916 16660
rect 35308 17052 35364 17108
rect 35532 16828 35588 16884
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35196 15874 35252 15876
rect 35196 15822 35198 15874
rect 35198 15822 35250 15874
rect 35250 15822 35252 15874
rect 35196 15820 35252 15822
rect 34860 13804 34916 13860
rect 34748 12402 34804 12404
rect 34748 12350 34750 12402
rect 34750 12350 34802 12402
rect 34802 12350 34804 12402
rect 34748 12348 34804 12350
rect 34860 11228 34916 11284
rect 34860 9938 34916 9940
rect 34860 9886 34862 9938
rect 34862 9886 34914 9938
rect 34914 9886 34916 9938
rect 34860 9884 34916 9886
rect 34748 9772 34804 9828
rect 35196 15036 35252 15092
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35308 14476 35364 14532
rect 35644 16716 35700 16772
rect 36092 17388 36148 17444
rect 35980 17276 36036 17332
rect 35980 16828 36036 16884
rect 36316 17276 36372 17332
rect 36316 16882 36372 16884
rect 36316 16830 36318 16882
rect 36318 16830 36370 16882
rect 36370 16830 36372 16882
rect 36316 16828 36372 16830
rect 36652 20972 36708 21028
rect 36540 19068 36596 19124
rect 36652 20412 36708 20468
rect 36540 18450 36596 18452
rect 36540 18398 36542 18450
rect 36542 18398 36594 18450
rect 36594 18398 36596 18450
rect 36540 18396 36596 18398
rect 37100 21698 37156 21700
rect 37100 21646 37102 21698
rect 37102 21646 37154 21698
rect 37154 21646 37156 21698
rect 37100 21644 37156 21646
rect 38444 27244 38500 27300
rect 38220 27132 38276 27188
rect 38444 27020 38500 27076
rect 38108 26908 38164 26964
rect 37772 26012 37828 26068
rect 37996 26402 38052 26404
rect 37996 26350 37998 26402
rect 37998 26350 38050 26402
rect 38050 26350 38052 26402
rect 37996 26348 38052 26350
rect 37660 25506 37716 25508
rect 37660 25454 37662 25506
rect 37662 25454 37714 25506
rect 37714 25454 37716 25506
rect 37660 25452 37716 25454
rect 37884 25394 37940 25396
rect 37884 25342 37886 25394
rect 37886 25342 37938 25394
rect 37938 25342 37940 25394
rect 37884 25340 37940 25342
rect 37324 24834 37380 24836
rect 37324 24782 37326 24834
rect 37326 24782 37378 24834
rect 37378 24782 37380 24834
rect 37324 24780 37380 24782
rect 37772 25004 37828 25060
rect 37436 23772 37492 23828
rect 37436 23548 37492 23604
rect 37548 22652 37604 22708
rect 38220 26236 38276 26292
rect 38108 25730 38164 25732
rect 38108 25678 38110 25730
rect 38110 25678 38162 25730
rect 38162 25678 38164 25730
rect 38108 25676 38164 25678
rect 38444 26012 38500 26068
rect 38332 25788 38388 25844
rect 38332 25340 38388 25396
rect 38332 25116 38388 25172
rect 38668 26962 38724 26964
rect 38668 26910 38670 26962
rect 38670 26910 38722 26962
rect 38722 26910 38724 26962
rect 38668 26908 38724 26910
rect 38668 24834 38724 24836
rect 38668 24782 38670 24834
rect 38670 24782 38722 24834
rect 38722 24782 38724 24834
rect 38668 24780 38724 24782
rect 38892 27244 38948 27300
rect 38892 26796 38948 26852
rect 38892 25900 38948 25956
rect 39228 26796 39284 26852
rect 39340 26290 39396 26292
rect 39340 26238 39342 26290
rect 39342 26238 39394 26290
rect 39394 26238 39396 26290
rect 39340 26236 39396 26238
rect 39116 26012 39172 26068
rect 39004 25788 39060 25844
rect 39228 25788 39284 25844
rect 39116 25506 39172 25508
rect 39116 25454 39118 25506
rect 39118 25454 39170 25506
rect 39170 25454 39172 25506
rect 39116 25452 39172 25454
rect 37772 22652 37828 22708
rect 37996 22482 38052 22484
rect 37996 22430 37998 22482
rect 37998 22430 38050 22482
rect 38050 22430 38052 22482
rect 37996 22428 38052 22430
rect 36988 20636 37044 20692
rect 37324 20242 37380 20244
rect 37324 20190 37326 20242
rect 37326 20190 37378 20242
rect 37378 20190 37380 20242
rect 37324 20188 37380 20190
rect 37212 20076 37268 20132
rect 37100 19740 37156 19796
rect 37996 22146 38052 22148
rect 37996 22094 37998 22146
rect 37998 22094 38050 22146
rect 38050 22094 38052 22146
rect 37996 22092 38052 22094
rect 38668 23436 38724 23492
rect 39340 25506 39396 25508
rect 39340 25454 39342 25506
rect 39342 25454 39394 25506
rect 39394 25454 39396 25506
rect 39340 25452 39396 25454
rect 39340 25228 39396 25284
rect 40012 27858 40068 27860
rect 40012 27806 40014 27858
rect 40014 27806 40066 27858
rect 40066 27806 40068 27858
rect 40012 27804 40068 27806
rect 39676 27186 39732 27188
rect 39676 27134 39678 27186
rect 39678 27134 39730 27186
rect 39730 27134 39732 27186
rect 39676 27132 39732 27134
rect 40572 31388 40628 31444
rect 40460 30828 40516 30884
rect 40908 30604 40964 30660
rect 41916 51996 41972 52052
rect 41580 51100 41636 51156
rect 41804 49922 41860 49924
rect 41804 49870 41806 49922
rect 41806 49870 41858 49922
rect 41858 49870 41860 49922
rect 41804 49868 41860 49870
rect 41692 48076 41748 48132
rect 41804 47740 41860 47796
rect 41916 47068 41972 47124
rect 41804 44322 41860 44324
rect 41804 44270 41806 44322
rect 41806 44270 41858 44322
rect 41858 44270 41860 44322
rect 41804 44268 41860 44270
rect 41804 43538 41860 43540
rect 41804 43486 41806 43538
rect 41806 43486 41858 43538
rect 41858 43486 41860 43538
rect 41804 43484 41860 43486
rect 41468 41970 41524 41972
rect 41468 41918 41470 41970
rect 41470 41918 41522 41970
rect 41522 41918 41524 41970
rect 41468 41916 41524 41918
rect 41692 40460 41748 40516
rect 41356 39676 41412 39732
rect 41804 40236 41860 40292
rect 41692 39564 41748 39620
rect 43036 53228 43092 53284
rect 42476 53058 42532 53060
rect 42476 53006 42478 53058
rect 42478 53006 42530 53058
rect 42530 53006 42532 53058
rect 42476 53004 42532 53006
rect 42364 52834 42420 52836
rect 42364 52782 42366 52834
rect 42366 52782 42418 52834
rect 42418 52782 42420 52834
rect 42364 52780 42420 52782
rect 42252 52220 42308 52276
rect 42476 52668 42532 52724
rect 43372 55020 43428 55076
rect 43932 55580 43988 55636
rect 43708 54626 43764 54628
rect 43708 54574 43710 54626
rect 43710 54574 43762 54626
rect 43762 54574 43764 54626
rect 43708 54572 43764 54574
rect 43596 54460 43652 54516
rect 43596 54290 43652 54292
rect 43596 54238 43598 54290
rect 43598 54238 43650 54290
rect 43650 54238 43652 54290
rect 43596 54236 43652 54238
rect 43596 53228 43652 53284
rect 47516 56028 47572 56084
rect 44604 55410 44660 55412
rect 44604 55358 44606 55410
rect 44606 55358 44658 55410
rect 44658 55358 44660 55410
rect 44604 55356 44660 55358
rect 45836 55410 45892 55412
rect 45836 55358 45838 55410
rect 45838 55358 45890 55410
rect 45890 55358 45892 55410
rect 45836 55356 45892 55358
rect 44492 55298 44548 55300
rect 44492 55246 44494 55298
rect 44494 55246 44546 55298
rect 44546 55246 44548 55298
rect 44492 55244 44548 55246
rect 44716 55074 44772 55076
rect 44716 55022 44718 55074
rect 44718 55022 44770 55074
rect 44770 55022 44772 55074
rect 44716 55020 44772 55022
rect 44156 54626 44212 54628
rect 44156 54574 44158 54626
rect 44158 54574 44210 54626
rect 44210 54574 44212 54626
rect 44156 54572 44212 54574
rect 44044 54236 44100 54292
rect 44044 53506 44100 53508
rect 44044 53454 44046 53506
rect 44046 53454 44098 53506
rect 44098 53454 44100 53506
rect 44044 53452 44100 53454
rect 44492 53452 44548 53508
rect 42364 51996 42420 52052
rect 42252 49868 42308 49924
rect 42140 48748 42196 48804
rect 43260 51884 43316 51940
rect 43932 52108 43988 52164
rect 43596 51324 43652 51380
rect 42476 49922 42532 49924
rect 42476 49870 42478 49922
rect 42478 49870 42530 49922
rect 42530 49870 42532 49922
rect 42476 49868 42532 49870
rect 42364 46396 42420 46452
rect 42812 49644 42868 49700
rect 42364 44604 42420 44660
rect 42364 43708 42420 43764
rect 42364 43538 42420 43540
rect 42364 43486 42366 43538
rect 42366 43486 42418 43538
rect 42418 43486 42420 43538
rect 42364 43484 42420 43486
rect 42140 40572 42196 40628
rect 42028 39788 42084 39844
rect 42700 48914 42756 48916
rect 42700 48862 42702 48914
rect 42702 48862 42754 48914
rect 42754 48862 42756 48914
rect 42700 48860 42756 48862
rect 43484 49698 43540 49700
rect 43484 49646 43486 49698
rect 43486 49646 43538 49698
rect 43538 49646 43540 49698
rect 43484 49644 43540 49646
rect 43484 48914 43540 48916
rect 43484 48862 43486 48914
rect 43486 48862 43538 48914
rect 43538 48862 43540 48914
rect 43484 48860 43540 48862
rect 43036 48300 43092 48356
rect 43372 48748 43428 48804
rect 43708 48802 43764 48804
rect 43708 48750 43710 48802
rect 43710 48750 43762 48802
rect 43762 48750 43764 48802
rect 43708 48748 43764 48750
rect 43932 48300 43988 48356
rect 43708 48130 43764 48132
rect 43708 48078 43710 48130
rect 43710 48078 43762 48130
rect 43762 48078 43764 48130
rect 43708 48076 43764 48078
rect 43372 47346 43428 47348
rect 43372 47294 43374 47346
rect 43374 47294 43426 47346
rect 43426 47294 43428 47346
rect 43372 47292 43428 47294
rect 44380 51996 44436 52052
rect 44380 51548 44436 51604
rect 44716 52386 44772 52388
rect 44716 52334 44718 52386
rect 44718 52334 44770 52386
rect 44770 52334 44772 52386
rect 44716 52332 44772 52334
rect 44604 51938 44660 51940
rect 44604 51886 44606 51938
rect 44606 51886 44658 51938
rect 44658 51886 44660 51938
rect 44604 51884 44660 51886
rect 46620 55186 46676 55188
rect 46620 55134 46622 55186
rect 46622 55134 46674 55186
rect 46674 55134 46676 55186
rect 46620 55132 46676 55134
rect 45836 54738 45892 54740
rect 45836 54686 45838 54738
rect 45838 54686 45890 54738
rect 45890 54686 45892 54738
rect 45836 54684 45892 54686
rect 45724 54012 45780 54068
rect 45388 52162 45444 52164
rect 45388 52110 45390 52162
rect 45390 52110 45442 52162
rect 45442 52110 45444 52162
rect 45388 52108 45444 52110
rect 44828 51378 44884 51380
rect 44828 51326 44830 51378
rect 44830 51326 44882 51378
rect 44882 51326 44884 51378
rect 44828 51324 44884 51326
rect 45052 51212 45108 51268
rect 46060 52332 46116 52388
rect 46060 51996 46116 52052
rect 45724 51266 45780 51268
rect 45724 51214 45726 51266
rect 45726 51214 45778 51266
rect 45778 51214 45780 51266
rect 45724 51212 45780 51214
rect 45836 51938 45892 51940
rect 45836 51886 45838 51938
rect 45838 51886 45890 51938
rect 45890 51886 45892 51938
rect 45836 51884 45892 51886
rect 45164 48860 45220 48916
rect 44716 48748 44772 48804
rect 45500 48748 45556 48804
rect 45612 48914 45668 48916
rect 45612 48862 45614 48914
rect 45614 48862 45666 48914
rect 45666 48862 45668 48914
rect 45612 48860 45668 48862
rect 44268 48354 44324 48356
rect 44268 48302 44270 48354
rect 44270 48302 44322 48354
rect 44322 48302 44324 48354
rect 44268 48300 44324 48302
rect 44492 48354 44548 48356
rect 44492 48302 44494 48354
rect 44494 48302 44546 48354
rect 44546 48302 44548 48354
rect 44492 48300 44548 48302
rect 44156 47180 44212 47236
rect 45388 48354 45444 48356
rect 45388 48302 45390 48354
rect 45390 48302 45442 48354
rect 45442 48302 45444 48354
rect 45388 48300 45444 48302
rect 45276 48130 45332 48132
rect 45276 48078 45278 48130
rect 45278 48078 45330 48130
rect 45330 48078 45332 48130
rect 45276 48076 45332 48078
rect 44604 47404 44660 47460
rect 44492 47068 44548 47124
rect 46060 47458 46116 47460
rect 46060 47406 46062 47458
rect 46062 47406 46114 47458
rect 46114 47406 46116 47458
rect 46060 47404 46116 47406
rect 44940 47180 44996 47236
rect 44380 45778 44436 45780
rect 44380 45726 44382 45778
rect 44382 45726 44434 45778
rect 44434 45726 44436 45778
rect 44380 45724 44436 45726
rect 42700 44492 42756 44548
rect 43484 44434 43540 44436
rect 43484 44382 43486 44434
rect 43486 44382 43538 44434
rect 43538 44382 43540 44434
rect 43484 44380 43540 44382
rect 43932 44268 43988 44324
rect 43148 44156 43204 44212
rect 44156 44380 44212 44436
rect 44268 44322 44324 44324
rect 44268 44270 44270 44322
rect 44270 44270 44322 44322
rect 44322 44270 44324 44322
rect 44268 44268 44324 44270
rect 44044 44156 44100 44212
rect 43372 43708 43428 43764
rect 42812 43596 42868 43652
rect 42700 43372 42756 43428
rect 43708 43650 43764 43652
rect 43708 43598 43710 43650
rect 43710 43598 43762 43650
rect 43762 43598 43764 43650
rect 43708 43596 43764 43598
rect 43260 43484 43316 43540
rect 43148 43314 43204 43316
rect 43148 43262 43150 43314
rect 43150 43262 43202 43314
rect 43202 43262 43204 43314
rect 43148 43260 43204 43262
rect 44156 43538 44212 43540
rect 44156 43486 44158 43538
rect 44158 43486 44210 43538
rect 44210 43486 44212 43538
rect 44156 43484 44212 43486
rect 44716 44322 44772 44324
rect 44716 44270 44718 44322
rect 44718 44270 44770 44322
rect 44770 44270 44772 44322
rect 44716 44268 44772 44270
rect 44380 43484 44436 43540
rect 44828 43538 44884 43540
rect 44828 43486 44830 43538
rect 44830 43486 44882 43538
rect 44882 43486 44884 43538
rect 44828 43484 44884 43486
rect 44156 43260 44212 43316
rect 44268 42754 44324 42756
rect 44268 42702 44270 42754
rect 44270 42702 44322 42754
rect 44322 42702 44324 42754
rect 44268 42700 44324 42702
rect 43708 42028 43764 42084
rect 43932 42028 43988 42084
rect 42924 41186 42980 41188
rect 42924 41134 42926 41186
rect 42926 41134 42978 41186
rect 42978 41134 42980 41186
rect 42924 41132 42980 41134
rect 43820 41186 43876 41188
rect 43820 41134 43822 41186
rect 43822 41134 43874 41186
rect 43874 41134 43876 41186
rect 43820 41132 43876 41134
rect 43260 40962 43316 40964
rect 43260 40910 43262 40962
rect 43262 40910 43314 40962
rect 43314 40910 43316 40962
rect 43260 40908 43316 40910
rect 43820 40908 43876 40964
rect 43708 40514 43764 40516
rect 43708 40462 43710 40514
rect 43710 40462 43762 40514
rect 43762 40462 43764 40514
rect 43708 40460 43764 40462
rect 42812 40348 42868 40404
rect 42364 38332 42420 38388
rect 43596 40402 43652 40404
rect 43596 40350 43598 40402
rect 43598 40350 43650 40402
rect 43650 40350 43652 40402
rect 43596 40348 43652 40350
rect 41916 38162 41972 38164
rect 41916 38110 41918 38162
rect 41918 38110 41970 38162
rect 41970 38110 41972 38162
rect 41916 38108 41972 38110
rect 41692 37996 41748 38052
rect 41356 36482 41412 36484
rect 41356 36430 41358 36482
rect 41358 36430 41410 36482
rect 41410 36430 41412 36482
rect 41356 36428 41412 36430
rect 41468 36258 41524 36260
rect 41468 36206 41470 36258
rect 41470 36206 41522 36258
rect 41522 36206 41524 36258
rect 41468 36204 41524 36206
rect 41804 36876 41860 36932
rect 42364 38050 42420 38052
rect 42364 37998 42366 38050
rect 42366 37998 42418 38050
rect 42418 37998 42420 38050
rect 42364 37996 42420 37998
rect 42588 38108 42644 38164
rect 42140 36316 42196 36372
rect 41804 36204 41860 36260
rect 41468 33346 41524 33348
rect 41468 33294 41470 33346
rect 41470 33294 41522 33346
rect 41522 33294 41524 33346
rect 41468 33292 41524 33294
rect 41132 33180 41188 33236
rect 41132 32284 41188 32340
rect 41468 31388 41524 31444
rect 43036 36988 43092 37044
rect 42476 36876 42532 36932
rect 42364 36316 42420 36372
rect 43148 36594 43204 36596
rect 43148 36542 43150 36594
rect 43150 36542 43202 36594
rect 43202 36542 43204 36594
rect 43148 36540 43204 36542
rect 42364 33964 42420 34020
rect 42252 31276 42308 31332
rect 43596 34524 43652 34580
rect 43932 40626 43988 40628
rect 43932 40574 43934 40626
rect 43934 40574 43986 40626
rect 43986 40574 43988 40626
rect 43932 40572 43988 40574
rect 45724 47234 45780 47236
rect 45724 47182 45726 47234
rect 45726 47182 45778 47234
rect 45778 47182 45780 47234
rect 45724 47180 45780 47182
rect 45500 45724 45556 45780
rect 45052 44268 45108 44324
rect 45500 44322 45556 44324
rect 45500 44270 45502 44322
rect 45502 44270 45554 44322
rect 45554 44270 45556 44322
rect 45500 44268 45556 44270
rect 45948 43538 46004 43540
rect 45948 43486 45950 43538
rect 45950 43486 46002 43538
rect 46002 43486 46004 43538
rect 45948 43484 46004 43486
rect 45164 40908 45220 40964
rect 44492 40514 44548 40516
rect 44492 40462 44494 40514
rect 44494 40462 44546 40514
rect 44546 40462 44548 40514
rect 44492 40460 44548 40462
rect 44380 40402 44436 40404
rect 44380 40350 44382 40402
rect 44382 40350 44434 40402
rect 44434 40350 44436 40402
rect 44380 40348 44436 40350
rect 46172 42700 46228 42756
rect 45724 41186 45780 41188
rect 45724 41134 45726 41186
rect 45726 41134 45778 41186
rect 45778 41134 45780 41186
rect 45724 41132 45780 41134
rect 45500 40572 45556 40628
rect 45388 40402 45444 40404
rect 45388 40350 45390 40402
rect 45390 40350 45442 40402
rect 45442 40350 45444 40402
rect 45388 40348 45444 40350
rect 45612 40460 45668 40516
rect 45612 36540 45668 36596
rect 43708 33516 43764 33572
rect 46284 33628 46340 33684
rect 43036 33404 43092 33460
rect 44492 33458 44548 33460
rect 44492 33406 44494 33458
rect 44494 33406 44546 33458
rect 44546 33406 44548 33458
rect 44492 33404 44548 33406
rect 46172 32450 46228 32452
rect 46172 32398 46174 32450
rect 46174 32398 46226 32450
rect 46226 32398 46228 32450
rect 46172 32396 46228 32398
rect 43596 31554 43652 31556
rect 43596 31502 43598 31554
rect 43598 31502 43650 31554
rect 43650 31502 43652 31554
rect 43596 31500 43652 31502
rect 46060 31164 46116 31220
rect 42252 30828 42308 30884
rect 41692 30098 41748 30100
rect 41692 30046 41694 30098
rect 41694 30046 41746 30098
rect 41746 30046 41748 30098
rect 41692 30044 41748 30046
rect 41356 29596 41412 29652
rect 40684 29484 40740 29540
rect 40348 28754 40404 28756
rect 40348 28702 40350 28754
rect 40350 28702 40402 28754
rect 40402 28702 40404 28754
rect 40348 28700 40404 28702
rect 40908 28812 40964 28868
rect 40796 28642 40852 28644
rect 40796 28590 40798 28642
rect 40798 28590 40850 28642
rect 40850 28590 40852 28642
rect 40796 28588 40852 28590
rect 40572 27020 40628 27076
rect 40124 26850 40180 26852
rect 40124 26798 40126 26850
rect 40126 26798 40178 26850
rect 40178 26798 40180 26850
rect 40124 26796 40180 26798
rect 39788 26402 39844 26404
rect 39788 26350 39790 26402
rect 39790 26350 39842 26402
rect 39842 26350 39844 26402
rect 39788 26348 39844 26350
rect 40124 25900 40180 25956
rect 40348 25676 40404 25732
rect 41356 28588 41412 28644
rect 42028 29708 42084 29764
rect 41916 29650 41972 29652
rect 41916 29598 41918 29650
rect 41918 29598 41970 29650
rect 41970 29598 41972 29650
rect 41916 29596 41972 29598
rect 41580 29538 41636 29540
rect 41580 29486 41582 29538
rect 41582 29486 41634 29538
rect 41634 29486 41636 29538
rect 41580 29484 41636 29486
rect 41468 28700 41524 28756
rect 41580 28812 41636 28868
rect 41132 27804 41188 27860
rect 41132 27020 41188 27076
rect 39564 25228 39620 25284
rect 40124 25228 40180 25284
rect 38780 22876 38836 22932
rect 38556 22316 38612 22372
rect 38108 21532 38164 21588
rect 37772 20188 37828 20244
rect 38444 20636 38500 20692
rect 38444 20412 38500 20468
rect 37884 19964 37940 20020
rect 37884 19740 37940 19796
rect 36876 18732 36932 18788
rect 36988 17948 37044 18004
rect 37100 18508 37156 18564
rect 36988 17500 37044 17556
rect 36764 17106 36820 17108
rect 36764 17054 36766 17106
rect 36766 17054 36818 17106
rect 36818 17054 36820 17106
rect 36764 17052 36820 17054
rect 35868 16658 35924 16660
rect 35868 16606 35870 16658
rect 35870 16606 35922 16658
rect 35922 16606 35924 16658
rect 35868 16604 35924 16606
rect 35980 15484 36036 15540
rect 36428 16322 36484 16324
rect 36428 16270 36430 16322
rect 36430 16270 36482 16322
rect 36482 16270 36484 16322
rect 36428 16268 36484 16270
rect 36764 16828 36820 16884
rect 36652 16156 36708 16212
rect 36652 15986 36708 15988
rect 36652 15934 36654 15986
rect 36654 15934 36706 15986
rect 36706 15934 36708 15986
rect 36652 15932 36708 15934
rect 36764 15820 36820 15876
rect 36988 17276 37044 17332
rect 36876 15596 36932 15652
rect 36988 16492 37044 16548
rect 36652 15148 36708 15204
rect 35756 14364 35812 14420
rect 35196 13970 35252 13972
rect 35196 13918 35198 13970
rect 35198 13918 35250 13970
rect 35250 13918 35252 13970
rect 35196 13916 35252 13918
rect 35868 14140 35924 14196
rect 36316 14252 36372 14308
rect 35756 13746 35812 13748
rect 35756 13694 35758 13746
rect 35758 13694 35810 13746
rect 35810 13694 35812 13746
rect 35756 13692 35812 13694
rect 35420 13580 35476 13636
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 36204 13580 36260 13636
rect 36540 13746 36596 13748
rect 36540 13694 36542 13746
rect 36542 13694 36594 13746
rect 36594 13694 36596 13746
rect 36540 13692 36596 13694
rect 35084 12348 35140 12404
rect 35532 12348 35588 12404
rect 35868 12348 35924 12404
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35084 11228 35140 11284
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35084 9996 35140 10052
rect 35532 9938 35588 9940
rect 35532 9886 35534 9938
rect 35534 9886 35586 9938
rect 35586 9886 35588 9938
rect 35532 9884 35588 9886
rect 36428 12236 36484 12292
rect 36204 12124 36260 12180
rect 36092 11954 36148 11956
rect 36092 11902 36094 11954
rect 36094 11902 36146 11954
rect 36146 11902 36148 11954
rect 36092 11900 36148 11902
rect 35980 11282 36036 11284
rect 35980 11230 35982 11282
rect 35982 11230 36034 11282
rect 36034 11230 36036 11282
rect 35980 11228 36036 11230
rect 36876 15036 36932 15092
rect 36988 14252 37044 14308
rect 37996 19010 38052 19012
rect 37996 18958 37998 19010
rect 37998 18958 38050 19010
rect 38050 18958 38052 19010
rect 37996 18956 38052 18958
rect 37884 18508 37940 18564
rect 37548 18396 37604 18452
rect 38332 19234 38388 19236
rect 38332 19182 38334 19234
rect 38334 19182 38386 19234
rect 38386 19182 38388 19234
rect 38332 19180 38388 19182
rect 38220 18508 38276 18564
rect 38108 18396 38164 18452
rect 37436 18338 37492 18340
rect 37436 18286 37438 18338
rect 37438 18286 37490 18338
rect 37490 18286 37492 18338
rect 37436 18284 37492 18286
rect 37996 18284 38052 18340
rect 37212 18172 37268 18228
rect 37436 17948 37492 18004
rect 37660 17554 37716 17556
rect 37660 17502 37662 17554
rect 37662 17502 37714 17554
rect 37714 17502 37716 17554
rect 37660 17500 37716 17502
rect 37548 17052 37604 17108
rect 37660 17276 37716 17332
rect 37436 16994 37492 16996
rect 37436 16942 37438 16994
rect 37438 16942 37490 16994
rect 37490 16942 37492 16994
rect 37436 16940 37492 16942
rect 37212 16604 37268 16660
rect 37436 16604 37492 16660
rect 37100 15484 37156 15540
rect 37100 15148 37156 15204
rect 37212 15708 37268 15764
rect 37772 17164 37828 17220
rect 37996 17052 38052 17108
rect 38108 17164 38164 17220
rect 38220 16994 38276 16996
rect 38220 16942 38222 16994
rect 38222 16942 38274 16994
rect 38274 16942 38276 16994
rect 38220 16940 38276 16942
rect 37772 16044 37828 16100
rect 37884 15932 37940 15988
rect 36876 13132 36932 13188
rect 36652 12572 36708 12628
rect 36764 12348 36820 12404
rect 36540 11116 36596 11172
rect 36316 10892 36372 10948
rect 35756 9938 35812 9940
rect 35756 9886 35758 9938
rect 35758 9886 35810 9938
rect 35810 9886 35812 9938
rect 35756 9884 35812 9886
rect 38108 15484 38164 15540
rect 38220 15596 38276 15652
rect 38220 15260 38276 15316
rect 38668 22146 38724 22148
rect 38668 22094 38670 22146
rect 38670 22094 38722 22146
rect 38722 22094 38724 22146
rect 38668 22092 38724 22094
rect 38892 22316 38948 22372
rect 39228 22258 39284 22260
rect 39228 22206 39230 22258
rect 39230 22206 39282 22258
rect 39282 22206 39284 22258
rect 39228 22204 39284 22206
rect 40348 25116 40404 25172
rect 40572 26124 40628 26180
rect 41580 27970 41636 27972
rect 41580 27918 41582 27970
rect 41582 27918 41634 27970
rect 41634 27918 41636 27970
rect 41580 27916 41636 27918
rect 41916 27858 41972 27860
rect 41916 27806 41918 27858
rect 41918 27806 41970 27858
rect 41970 27806 41972 27858
rect 41916 27804 41972 27806
rect 41916 27356 41972 27412
rect 41580 27074 41636 27076
rect 41580 27022 41582 27074
rect 41582 27022 41634 27074
rect 41634 27022 41636 27074
rect 41580 27020 41636 27022
rect 41356 26124 41412 26180
rect 41132 25788 41188 25844
rect 40684 25452 40740 25508
rect 40908 25340 40964 25396
rect 40572 24780 40628 24836
rect 39788 23996 39844 24052
rect 39676 23436 39732 23492
rect 40236 23548 40292 23604
rect 41132 25394 41188 25396
rect 41132 25342 41134 25394
rect 41134 25342 41186 25394
rect 41186 25342 41188 25394
rect 41132 25340 41188 25342
rect 41468 24610 41524 24612
rect 41468 24558 41470 24610
rect 41470 24558 41522 24610
rect 41522 24558 41524 24610
rect 41468 24556 41524 24558
rect 41804 25900 41860 25956
rect 42028 26684 42084 26740
rect 42140 26178 42196 26180
rect 42140 26126 42142 26178
rect 42142 26126 42194 26178
rect 42194 26126 42196 26178
rect 42140 26124 42196 26126
rect 43820 30716 43876 30772
rect 42364 30156 42420 30212
rect 42364 29650 42420 29652
rect 42364 29598 42366 29650
rect 42366 29598 42418 29650
rect 42418 29598 42420 29650
rect 42364 29596 42420 29598
rect 42476 30098 42532 30100
rect 42476 30046 42478 30098
rect 42478 30046 42530 30098
rect 42530 30046 42532 30098
rect 42476 30044 42532 30046
rect 43932 30210 43988 30212
rect 43932 30158 43934 30210
rect 43934 30158 43986 30210
rect 43986 30158 43988 30210
rect 43932 30156 43988 30158
rect 43820 30044 43876 30100
rect 43708 29708 43764 29764
rect 43260 29650 43316 29652
rect 43260 29598 43262 29650
rect 43262 29598 43314 29650
rect 43314 29598 43316 29650
rect 43260 29596 43316 29598
rect 42700 28812 42756 28868
rect 42588 28364 42644 28420
rect 42700 27692 42756 27748
rect 44492 30940 44548 30996
rect 44156 30098 44212 30100
rect 44156 30046 44158 30098
rect 44158 30046 44210 30098
rect 44210 30046 44212 30098
rect 44156 30044 44212 30046
rect 44044 29708 44100 29764
rect 44380 29650 44436 29652
rect 44380 29598 44382 29650
rect 44382 29598 44434 29650
rect 44434 29598 44436 29650
rect 44380 29596 44436 29598
rect 45724 30994 45780 30996
rect 45724 30942 45726 30994
rect 45726 30942 45778 30994
rect 45778 30942 45780 30994
rect 45724 30940 45780 30942
rect 45388 30828 45444 30884
rect 45388 30044 45444 30100
rect 44716 29708 44772 29764
rect 44828 29538 44884 29540
rect 44828 29486 44830 29538
rect 44830 29486 44882 29538
rect 44882 29486 44884 29538
rect 44828 29484 44884 29486
rect 43484 28530 43540 28532
rect 43484 28478 43486 28530
rect 43486 28478 43538 28530
rect 43538 28478 43540 28530
rect 43484 28476 43540 28478
rect 42812 27580 42868 27636
rect 42924 28364 42980 28420
rect 42588 27356 42644 27412
rect 42364 26962 42420 26964
rect 42364 26910 42366 26962
rect 42366 26910 42418 26962
rect 42418 26910 42420 26962
rect 42364 26908 42420 26910
rect 42588 26850 42644 26852
rect 42588 26798 42590 26850
rect 42590 26798 42642 26850
rect 42642 26798 42644 26850
rect 42588 26796 42644 26798
rect 42252 25282 42308 25284
rect 42252 25230 42254 25282
rect 42254 25230 42306 25282
rect 42306 25230 42308 25282
rect 42252 25228 42308 25230
rect 42364 26684 42420 26740
rect 42588 24780 42644 24836
rect 43036 27916 43092 27972
rect 43372 27916 43428 27972
rect 43148 27804 43204 27860
rect 42924 26908 42980 26964
rect 43260 26908 43316 26964
rect 43148 26348 43204 26404
rect 43148 25618 43204 25620
rect 43148 25566 43150 25618
rect 43150 25566 43202 25618
rect 43202 25566 43204 25618
rect 43148 25564 43204 25566
rect 43260 25452 43316 25508
rect 41020 23660 41076 23716
rect 40460 23324 40516 23380
rect 40012 22482 40068 22484
rect 40012 22430 40014 22482
rect 40014 22430 40066 22482
rect 40066 22430 40068 22482
rect 40012 22428 40068 22430
rect 38780 21756 38836 21812
rect 39340 22092 39396 22148
rect 38668 21644 38724 21700
rect 39452 21810 39508 21812
rect 39452 21758 39454 21810
rect 39454 21758 39506 21810
rect 39506 21758 39508 21810
rect 39452 21756 39508 21758
rect 38780 21084 38836 21140
rect 39452 21532 39508 21588
rect 39564 21420 39620 21476
rect 38668 20802 38724 20804
rect 38668 20750 38670 20802
rect 38670 20750 38722 20802
rect 38722 20750 38724 20802
rect 38668 20748 38724 20750
rect 39340 20748 39396 20804
rect 39004 20130 39060 20132
rect 39004 20078 39006 20130
rect 39006 20078 39058 20130
rect 39058 20078 39060 20130
rect 39004 20076 39060 20078
rect 39452 20300 39508 20356
rect 39564 20076 39620 20132
rect 38780 19516 38836 19572
rect 38892 19180 38948 19236
rect 37548 14252 37604 14308
rect 38108 13692 38164 13748
rect 37996 12908 38052 12964
rect 38556 18508 38612 18564
rect 39340 19404 39396 19460
rect 39116 19122 39172 19124
rect 39116 19070 39118 19122
rect 39118 19070 39170 19122
rect 39170 19070 39172 19122
rect 39116 19068 39172 19070
rect 39228 19292 39284 19348
rect 39004 19010 39060 19012
rect 39004 18958 39006 19010
rect 39006 18958 39058 19010
rect 39058 18958 39060 19010
rect 39004 18956 39060 18958
rect 40348 23154 40404 23156
rect 40348 23102 40350 23154
rect 40350 23102 40402 23154
rect 40402 23102 40404 23154
rect 40348 23100 40404 23102
rect 40236 22258 40292 22260
rect 40236 22206 40238 22258
rect 40238 22206 40290 22258
rect 40290 22206 40292 22258
rect 40236 22204 40292 22206
rect 39900 22092 39956 22148
rect 39900 20188 39956 20244
rect 39900 19740 39956 19796
rect 40012 19292 40068 19348
rect 40124 22092 40180 22148
rect 39676 19180 39732 19236
rect 40012 19122 40068 19124
rect 40012 19070 40014 19122
rect 40014 19070 40066 19122
rect 40066 19070 40068 19122
rect 40012 19068 40068 19070
rect 40572 22428 40628 22484
rect 40796 22988 40852 23044
rect 40460 21980 40516 22036
rect 40684 22316 40740 22372
rect 40236 21810 40292 21812
rect 40236 21758 40238 21810
rect 40238 21758 40290 21810
rect 40290 21758 40292 21810
rect 40236 21756 40292 21758
rect 40460 21586 40516 21588
rect 40460 21534 40462 21586
rect 40462 21534 40514 21586
rect 40514 21534 40516 21586
rect 40460 21532 40516 21534
rect 40908 22258 40964 22260
rect 40908 22206 40910 22258
rect 40910 22206 40962 22258
rect 40962 22206 40964 22258
rect 40908 22204 40964 22206
rect 40908 21308 40964 21364
rect 40348 20524 40404 20580
rect 40348 20130 40404 20132
rect 40348 20078 40350 20130
rect 40350 20078 40402 20130
rect 40402 20078 40404 20130
rect 40348 20076 40404 20078
rect 40908 20300 40964 20356
rect 39564 18844 39620 18900
rect 40684 19516 40740 19572
rect 39004 18508 39060 18564
rect 38892 18284 38948 18340
rect 38668 17442 38724 17444
rect 38668 17390 38670 17442
rect 38670 17390 38722 17442
rect 38722 17390 38724 17442
rect 38668 17388 38724 17390
rect 39228 18284 39284 18340
rect 39116 18172 39172 18228
rect 39004 17890 39060 17892
rect 39004 17838 39006 17890
rect 39006 17838 39058 17890
rect 39058 17838 39060 17890
rect 39004 17836 39060 17838
rect 38780 16940 38836 16996
rect 38668 16098 38724 16100
rect 38668 16046 38670 16098
rect 38670 16046 38722 16098
rect 38722 16046 38724 16098
rect 38668 16044 38724 16046
rect 39228 17666 39284 17668
rect 39228 17614 39230 17666
rect 39230 17614 39282 17666
rect 39282 17614 39284 17666
rect 39228 17612 39284 17614
rect 39900 18284 39956 18340
rect 40012 18396 40068 18452
rect 39900 17890 39956 17892
rect 39900 17838 39902 17890
rect 39902 17838 39954 17890
rect 39954 17838 39956 17890
rect 39900 17836 39956 17838
rect 40236 18060 40292 18116
rect 40348 18396 40404 18452
rect 40796 19404 40852 19460
rect 40796 18620 40852 18676
rect 40460 17500 40516 17556
rect 39900 17164 39956 17220
rect 39676 16940 39732 16996
rect 39452 16882 39508 16884
rect 39452 16830 39454 16882
rect 39454 16830 39506 16882
rect 39506 16830 39508 16882
rect 39452 16828 39508 16830
rect 39340 16044 39396 16100
rect 39116 15596 39172 15652
rect 39564 15372 39620 15428
rect 38444 14364 38500 14420
rect 38444 12908 38500 12964
rect 37100 12290 37156 12292
rect 37100 12238 37102 12290
rect 37102 12238 37154 12290
rect 37154 12238 37156 12290
rect 37100 12236 37156 12238
rect 37212 12178 37268 12180
rect 37212 12126 37214 12178
rect 37214 12126 37266 12178
rect 37266 12126 37268 12178
rect 37212 12124 37268 12126
rect 37324 11900 37380 11956
rect 37100 10892 37156 10948
rect 37884 12124 37940 12180
rect 37548 11788 37604 11844
rect 39228 14530 39284 14532
rect 39228 14478 39230 14530
rect 39230 14478 39282 14530
rect 39282 14478 39284 14530
rect 39228 14476 39284 14478
rect 38780 14140 38836 14196
rect 38892 14252 38948 14308
rect 38668 13916 38724 13972
rect 39004 13916 39060 13972
rect 39564 14306 39620 14308
rect 39564 14254 39566 14306
rect 39566 14254 39618 14306
rect 39618 14254 39620 14306
rect 39564 14252 39620 14254
rect 40684 17164 40740 17220
rect 40684 16994 40740 16996
rect 40684 16942 40686 16994
rect 40686 16942 40738 16994
rect 40738 16942 40740 16994
rect 40684 16940 40740 16942
rect 40236 15708 40292 15764
rect 40348 15596 40404 15652
rect 40124 14924 40180 14980
rect 40684 15036 40740 15092
rect 41468 23436 41524 23492
rect 41132 22988 41188 23044
rect 41356 23324 41412 23380
rect 41356 22316 41412 22372
rect 41132 22204 41188 22260
rect 41244 21980 41300 22036
rect 41468 21980 41524 22036
rect 41356 21084 41412 21140
rect 41244 20972 41300 21028
rect 41132 19740 41188 19796
rect 41132 17948 41188 18004
rect 41244 17836 41300 17892
rect 41244 17388 41300 17444
rect 41804 23660 41860 23716
rect 42028 23714 42084 23716
rect 42028 23662 42030 23714
rect 42030 23662 42082 23714
rect 42082 23662 42084 23714
rect 42028 23660 42084 23662
rect 42364 23938 42420 23940
rect 42364 23886 42366 23938
rect 42366 23886 42418 23938
rect 42418 23886 42420 23938
rect 42364 23884 42420 23886
rect 42140 23212 42196 23268
rect 42252 22764 42308 22820
rect 41916 21756 41972 21812
rect 42028 22652 42084 22708
rect 41468 19740 41524 19796
rect 41580 19010 41636 19012
rect 41580 18958 41582 19010
rect 41582 18958 41634 19010
rect 41634 18958 41636 19010
rect 41580 18956 41636 18958
rect 41916 21308 41972 21364
rect 42028 20972 42084 21028
rect 41580 17052 41636 17108
rect 41468 16882 41524 16884
rect 41468 16830 41470 16882
rect 41470 16830 41522 16882
rect 41522 16830 41524 16882
rect 41468 16828 41524 16830
rect 40012 14140 40068 14196
rect 40796 14530 40852 14532
rect 40796 14478 40798 14530
rect 40798 14478 40850 14530
rect 40850 14478 40852 14530
rect 40796 14476 40852 14478
rect 40684 14418 40740 14420
rect 40684 14366 40686 14418
rect 40686 14366 40738 14418
rect 40738 14366 40740 14418
rect 40684 14364 40740 14366
rect 39676 13858 39732 13860
rect 39676 13806 39678 13858
rect 39678 13806 39730 13858
rect 39730 13806 39732 13858
rect 39676 13804 39732 13806
rect 39452 13356 39508 13412
rect 39676 13468 39732 13524
rect 39116 12796 39172 12852
rect 39228 13244 39284 13300
rect 39116 12572 39172 12628
rect 38780 12178 38836 12180
rect 38780 12126 38782 12178
rect 38782 12126 38834 12178
rect 38834 12126 38836 12178
rect 38780 12124 38836 12126
rect 38556 11788 38612 11844
rect 38892 11676 38948 11732
rect 39452 13074 39508 13076
rect 39452 13022 39454 13074
rect 39454 13022 39506 13074
rect 39506 13022 39508 13074
rect 39452 13020 39508 13022
rect 39340 12908 39396 12964
rect 40236 13916 40292 13972
rect 39900 13746 39956 13748
rect 39900 13694 39902 13746
rect 39902 13694 39954 13746
rect 39954 13694 39956 13746
rect 39900 13692 39956 13694
rect 39788 13020 39844 13076
rect 35868 9660 35924 9716
rect 35980 9996 36036 10052
rect 35420 9436 35476 9492
rect 35868 9436 35924 9492
rect 34636 9212 34692 9268
rect 35196 9212 35252 9268
rect 34636 8370 34692 8372
rect 34636 8318 34638 8370
rect 34638 8318 34690 8370
rect 34690 8318 34692 8370
rect 34636 8316 34692 8318
rect 35532 9154 35588 9156
rect 35532 9102 35534 9154
rect 35534 9102 35586 9154
rect 35586 9102 35588 9154
rect 35532 9100 35588 9102
rect 36540 9772 36596 9828
rect 36092 9714 36148 9716
rect 36092 9662 36094 9714
rect 36094 9662 36146 9714
rect 36146 9662 36148 9714
rect 36092 9660 36148 9662
rect 36764 9826 36820 9828
rect 36764 9774 36766 9826
rect 36766 9774 36818 9826
rect 36818 9774 36820 9826
rect 36764 9772 36820 9774
rect 35868 9100 35924 9156
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35532 8316 35588 8372
rect 36316 9042 36372 9044
rect 36316 8990 36318 9042
rect 36318 8990 36370 9042
rect 36370 8990 36372 9042
rect 36316 8988 36372 8990
rect 36092 8428 36148 8484
rect 35084 7980 35140 8036
rect 35196 8092 35252 8148
rect 34636 7868 34692 7924
rect 34524 7420 34580 7476
rect 35084 7250 35140 7252
rect 35084 7198 35086 7250
rect 35086 7198 35138 7250
rect 35138 7198 35140 7250
rect 35084 7196 35140 7198
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35308 6748 35364 6804
rect 33740 6636 33796 6692
rect 34636 6690 34692 6692
rect 34636 6638 34638 6690
rect 34638 6638 34690 6690
rect 34690 6638 34692 6690
rect 34636 6636 34692 6638
rect 35084 6466 35140 6468
rect 35084 6414 35086 6466
rect 35086 6414 35138 6466
rect 35138 6414 35140 6466
rect 35084 6412 35140 6414
rect 33740 6076 33796 6132
rect 33628 6018 33684 6020
rect 33628 5966 33630 6018
rect 33630 5966 33682 6018
rect 33682 5966 33684 6018
rect 33628 5964 33684 5966
rect 33964 5906 34020 5908
rect 33964 5854 33966 5906
rect 33966 5854 34018 5906
rect 34018 5854 34020 5906
rect 33964 5852 34020 5854
rect 35532 6412 35588 6468
rect 35196 5852 35252 5908
rect 35756 5906 35812 5908
rect 35756 5854 35758 5906
rect 35758 5854 35810 5906
rect 35810 5854 35812 5906
rect 35756 5852 35812 5854
rect 36764 8930 36820 8932
rect 36764 8878 36766 8930
rect 36766 8878 36818 8930
rect 36818 8878 36820 8930
rect 36764 8876 36820 8878
rect 36428 8370 36484 8372
rect 36428 8318 36430 8370
rect 36430 8318 36482 8370
rect 36482 8318 36484 8370
rect 36428 8316 36484 8318
rect 36540 8204 36596 8260
rect 36540 7586 36596 7588
rect 36540 7534 36542 7586
rect 36542 7534 36594 7586
rect 36594 7534 36596 7586
rect 36540 7532 36596 7534
rect 36204 6748 36260 6804
rect 36540 6748 36596 6804
rect 36316 6636 36372 6692
rect 35980 6412 36036 6468
rect 34188 5794 34244 5796
rect 34188 5742 34190 5794
rect 34190 5742 34242 5794
rect 34242 5742 34244 5794
rect 34188 5740 34244 5742
rect 33740 5292 33796 5348
rect 35308 5794 35364 5796
rect 35308 5742 35310 5794
rect 35310 5742 35362 5794
rect 35362 5742 35364 5794
rect 35308 5740 35364 5742
rect 35980 5794 36036 5796
rect 35980 5742 35982 5794
rect 35982 5742 36034 5794
rect 36034 5742 36036 5794
rect 35980 5740 36036 5742
rect 36652 5794 36708 5796
rect 36652 5742 36654 5794
rect 36654 5742 36706 5794
rect 36706 5742 36708 5794
rect 36652 5740 36708 5742
rect 34636 5516 34692 5572
rect 34524 5180 34580 5236
rect 33516 4956 33572 5012
rect 33516 4620 33572 4676
rect 33852 4396 33908 4452
rect 33292 1484 33348 1540
rect 33628 3612 33684 3668
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 36540 5234 36596 5236
rect 36540 5182 36542 5234
rect 36542 5182 36594 5234
rect 36594 5182 36596 5234
rect 36540 5180 36596 5182
rect 34972 4338 35028 4340
rect 34972 4286 34974 4338
rect 34974 4286 35026 4338
rect 35026 4286 35028 4338
rect 34972 4284 35028 4286
rect 35644 4284 35700 4340
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 34524 3666 34580 3668
rect 34524 3614 34526 3666
rect 34526 3614 34578 3666
rect 34578 3614 34580 3666
rect 34524 3612 34580 3614
rect 36988 8316 37044 8372
rect 37212 8316 37268 8372
rect 37548 8258 37604 8260
rect 37548 8206 37550 8258
rect 37550 8206 37602 8258
rect 37602 8206 37604 8258
rect 37548 8204 37604 8206
rect 36988 7756 37044 7812
rect 38668 10722 38724 10724
rect 38668 10670 38670 10722
rect 38670 10670 38722 10722
rect 38722 10670 38724 10722
rect 38668 10668 38724 10670
rect 38668 10220 38724 10276
rect 38556 9826 38612 9828
rect 38556 9774 38558 9826
rect 38558 9774 38610 9826
rect 38610 9774 38612 9826
rect 38556 9772 38612 9774
rect 40348 13858 40404 13860
rect 40348 13806 40350 13858
rect 40350 13806 40402 13858
rect 40402 13806 40404 13858
rect 40348 13804 40404 13806
rect 40684 13468 40740 13524
rect 40348 13356 40404 13412
rect 40348 12738 40404 12740
rect 40348 12686 40350 12738
rect 40350 12686 40402 12738
rect 40402 12686 40404 12738
rect 40348 12684 40404 12686
rect 40572 13020 40628 13076
rect 40572 12290 40628 12292
rect 40572 12238 40574 12290
rect 40574 12238 40626 12290
rect 40626 12238 40628 12290
rect 40572 12236 40628 12238
rect 40684 11900 40740 11956
rect 41020 13692 41076 13748
rect 41468 15036 41524 15092
rect 41580 14924 41636 14980
rect 41804 18396 41860 18452
rect 42028 19346 42084 19348
rect 42028 19294 42030 19346
rect 42030 19294 42082 19346
rect 42082 19294 42084 19346
rect 42028 19292 42084 19294
rect 42140 18732 42196 18788
rect 42476 22988 42532 23044
rect 42924 23660 42980 23716
rect 42588 22540 42644 22596
rect 42700 23100 42756 23156
rect 42588 22370 42644 22372
rect 42588 22318 42590 22370
rect 42590 22318 42642 22370
rect 42642 22318 42644 22370
rect 42588 22316 42644 22318
rect 42812 22764 42868 22820
rect 42364 21644 42420 21700
rect 42476 21420 42532 21476
rect 42364 20802 42420 20804
rect 42364 20750 42366 20802
rect 42366 20750 42418 20802
rect 42418 20750 42420 20802
rect 42364 20748 42420 20750
rect 43036 22988 43092 23044
rect 43372 25340 43428 25396
rect 43148 22316 43204 22372
rect 43036 22146 43092 22148
rect 43036 22094 43038 22146
rect 43038 22094 43090 22146
rect 43090 22094 43092 22146
rect 43036 22092 43092 22094
rect 43596 27580 43652 27636
rect 43596 27356 43652 27412
rect 43820 28418 43876 28420
rect 43820 28366 43822 28418
rect 43822 28366 43874 28418
rect 43874 28366 43876 28418
rect 43820 28364 43876 28366
rect 43820 27692 43876 27748
rect 43820 27132 43876 27188
rect 44156 26796 44212 26852
rect 43820 26236 43876 26292
rect 43708 25564 43764 25620
rect 44492 27916 44548 27972
rect 44716 27916 44772 27972
rect 44492 27468 44548 27524
rect 44492 26962 44548 26964
rect 44492 26910 44494 26962
rect 44494 26910 44546 26962
rect 44546 26910 44548 26962
rect 44492 26908 44548 26910
rect 46060 30940 46116 30996
rect 46172 30380 46228 30436
rect 45948 29596 46004 29652
rect 45836 29260 45892 29316
rect 46060 29260 46116 29316
rect 45948 28924 46004 28980
rect 46620 33180 46676 33236
rect 47180 55186 47236 55188
rect 47180 55134 47182 55186
rect 47182 55134 47234 55186
rect 47234 55134 47236 55186
rect 47180 55132 47236 55134
rect 55804 57148 55860 57204
rect 52780 56082 52836 56084
rect 52780 56030 52782 56082
rect 52782 56030 52834 56082
rect 52834 56030 52836 56082
rect 52780 56028 52836 56030
rect 51772 55916 51828 55972
rect 53452 55970 53508 55972
rect 53452 55918 53454 55970
rect 53454 55918 53506 55970
rect 53506 55918 53508 55970
rect 53452 55916 53508 55918
rect 56028 55410 56084 55412
rect 56028 55358 56030 55410
rect 56030 55358 56082 55410
rect 56082 55358 56084 55410
rect 56028 55356 56084 55358
rect 57148 55356 57204 55412
rect 47068 54908 47124 54964
rect 46844 40402 46900 40404
rect 46844 40350 46846 40402
rect 46846 40350 46898 40402
rect 46898 40350 46900 40402
rect 46844 40348 46900 40350
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 49532 53788 49588 53844
rect 48748 52108 48804 52164
rect 47404 48914 47460 48916
rect 47404 48862 47406 48914
rect 47406 48862 47458 48914
rect 47458 48862 47460 48914
rect 47404 48860 47460 48862
rect 47852 40460 47908 40516
rect 47852 35868 47908 35924
rect 47068 34860 47124 34916
rect 53900 53788 53956 53844
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 52892 52780 52948 52836
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 49532 34524 49588 34580
rect 52780 35756 52836 35812
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 52332 33628 52388 33684
rect 46732 32844 46788 32900
rect 47516 33180 47572 33236
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 51660 32674 51716 32676
rect 51660 32622 51662 32674
rect 51662 32622 51714 32674
rect 51714 32622 51716 32674
rect 51660 32620 51716 32622
rect 47516 32562 47572 32564
rect 47516 32510 47518 32562
rect 47518 32510 47570 32562
rect 47570 32510 47572 32562
rect 47516 32508 47572 32510
rect 48076 32396 48132 32452
rect 51100 32450 51156 32452
rect 51100 32398 51102 32450
rect 51102 32398 51154 32450
rect 51154 32398 51156 32450
rect 51100 32396 51156 32398
rect 51548 31778 51604 31780
rect 51548 31726 51550 31778
rect 51550 31726 51602 31778
rect 51602 31726 51604 31778
rect 51548 31724 51604 31726
rect 46284 29986 46340 29988
rect 46284 29934 46286 29986
rect 46286 29934 46338 29986
rect 46338 29934 46340 29986
rect 46284 29932 46340 29934
rect 46508 30994 46564 30996
rect 46508 30942 46510 30994
rect 46510 30942 46562 30994
rect 46562 30942 46564 30994
rect 46508 30940 46564 30942
rect 46844 30882 46900 30884
rect 46844 30830 46846 30882
rect 46846 30830 46898 30882
rect 46898 30830 46900 30882
rect 46844 30828 46900 30830
rect 47516 31554 47572 31556
rect 47516 31502 47518 31554
rect 47518 31502 47570 31554
rect 47570 31502 47572 31554
rect 47516 31500 47572 31502
rect 47852 31500 47908 31556
rect 48076 30940 48132 30996
rect 47180 30828 47236 30884
rect 46620 30156 46676 30212
rect 46172 28588 46228 28644
rect 46508 29596 46564 29652
rect 45276 26908 45332 26964
rect 44268 26066 44324 26068
rect 44268 26014 44270 26066
rect 44270 26014 44322 26066
rect 44322 26014 44324 26066
rect 44268 26012 44324 26014
rect 44156 25506 44212 25508
rect 44156 25454 44158 25506
rect 44158 25454 44210 25506
rect 44210 25454 44212 25506
rect 44156 25452 44212 25454
rect 44044 25116 44100 25172
rect 43708 23938 43764 23940
rect 43708 23886 43710 23938
rect 43710 23886 43762 23938
rect 43762 23886 43764 23938
rect 43708 23884 43764 23886
rect 43932 24556 43988 24612
rect 44044 24108 44100 24164
rect 44156 24220 44212 24276
rect 43596 23100 43652 23156
rect 43708 23548 43764 23604
rect 43932 23548 43988 23604
rect 43708 22652 43764 22708
rect 43820 23324 43876 23380
rect 43596 22540 43652 22596
rect 43148 21420 43204 21476
rect 43596 22204 43652 22260
rect 43036 21308 43092 21364
rect 42476 20300 42532 20356
rect 42252 18620 42308 18676
rect 42364 19516 42420 19572
rect 42140 18508 42196 18564
rect 41916 18172 41972 18228
rect 41916 17052 41972 17108
rect 42252 18338 42308 18340
rect 42252 18286 42254 18338
rect 42254 18286 42306 18338
rect 42306 18286 42308 18338
rect 42252 18284 42308 18286
rect 42476 18172 42532 18228
rect 43036 20412 43092 20468
rect 42812 19292 42868 19348
rect 44380 24722 44436 24724
rect 44380 24670 44382 24722
rect 44382 24670 44434 24722
rect 44434 24670 44436 24722
rect 44380 24668 44436 24670
rect 44492 23772 44548 23828
rect 44828 26460 44884 26516
rect 44604 24556 44660 24612
rect 44268 23436 44324 23492
rect 44380 23548 44436 23604
rect 44156 22876 44212 22932
rect 44156 22316 44212 22372
rect 43932 22092 43988 22148
rect 43484 20748 43540 20804
rect 43820 20802 43876 20804
rect 43820 20750 43822 20802
rect 43822 20750 43874 20802
rect 43874 20750 43876 20802
rect 43820 20748 43876 20750
rect 43708 20690 43764 20692
rect 43708 20638 43710 20690
rect 43710 20638 43762 20690
rect 43762 20638 43764 20690
rect 43708 20636 43764 20638
rect 43708 20300 43764 20356
rect 44044 21756 44100 21812
rect 44156 21980 44212 22036
rect 44044 20690 44100 20692
rect 44044 20638 44046 20690
rect 44046 20638 44098 20690
rect 44098 20638 44100 20690
rect 44044 20636 44100 20638
rect 44156 20578 44212 20580
rect 44156 20526 44158 20578
rect 44158 20526 44210 20578
rect 44210 20526 44212 20578
rect 44156 20524 44212 20526
rect 44604 23324 44660 23380
rect 44716 25452 44772 25508
rect 44492 22540 44548 22596
rect 44492 21980 44548 22036
rect 44156 20300 44212 20356
rect 43820 19906 43876 19908
rect 43820 19854 43822 19906
rect 43822 19854 43874 19906
rect 43874 19854 43876 19906
rect 43820 19852 43876 19854
rect 44380 21756 44436 21812
rect 44492 21532 44548 21588
rect 44492 20860 44548 20916
rect 44380 20300 44436 20356
rect 44268 19852 44324 19908
rect 43260 19180 43316 19236
rect 44380 19234 44436 19236
rect 44380 19182 44382 19234
rect 44382 19182 44434 19234
rect 44434 19182 44436 19234
rect 44380 19180 44436 19182
rect 43596 19068 43652 19124
rect 42812 18732 42868 18788
rect 42700 18284 42756 18340
rect 42252 17612 42308 17668
rect 41692 14700 41748 14756
rect 41692 14530 41748 14532
rect 41692 14478 41694 14530
rect 41694 14478 41746 14530
rect 41746 14478 41748 14530
rect 41692 14476 41748 14478
rect 41916 16044 41972 16100
rect 42140 16156 42196 16212
rect 42812 17612 42868 17668
rect 42588 17164 42644 17220
rect 42588 16940 42644 16996
rect 43596 18732 43652 18788
rect 44156 18844 44212 18900
rect 42924 17276 42980 17332
rect 43148 18620 43204 18676
rect 42700 16828 42756 16884
rect 43932 18674 43988 18676
rect 43932 18622 43934 18674
rect 43934 18622 43986 18674
rect 43986 18622 43988 18674
rect 43932 18620 43988 18622
rect 44044 18562 44100 18564
rect 44044 18510 44046 18562
rect 44046 18510 44098 18562
rect 44098 18510 44100 18562
rect 44044 18508 44100 18510
rect 43820 18450 43876 18452
rect 43820 18398 43822 18450
rect 43822 18398 43874 18450
rect 43874 18398 43876 18450
rect 43820 18396 43876 18398
rect 44716 21980 44772 22036
rect 44716 20972 44772 21028
rect 44828 19516 44884 19572
rect 45276 24220 45332 24276
rect 45052 23042 45108 23044
rect 45052 22990 45054 23042
rect 45054 22990 45106 23042
rect 45106 22990 45108 23042
rect 45052 22988 45108 22990
rect 45052 22204 45108 22260
rect 45052 21586 45108 21588
rect 45052 21534 45054 21586
rect 45054 21534 45106 21586
rect 45106 21534 45108 21586
rect 45052 21532 45108 21534
rect 45164 21420 45220 21476
rect 44940 19180 44996 19236
rect 45052 19516 45108 19572
rect 44380 18562 44436 18564
rect 44380 18510 44382 18562
rect 44382 18510 44434 18562
rect 44434 18510 44436 18562
rect 44380 18508 44436 18510
rect 44268 18396 44324 18452
rect 44492 18396 44548 18452
rect 43708 18172 43764 18228
rect 43372 17164 43428 17220
rect 42028 15596 42084 15652
rect 41916 14924 41972 14980
rect 41916 14700 41972 14756
rect 41356 14306 41412 14308
rect 41356 14254 41358 14306
rect 41358 14254 41410 14306
rect 41410 14254 41412 14306
rect 41356 14252 41412 14254
rect 41468 14140 41524 14196
rect 41356 13916 41412 13972
rect 41244 13468 41300 13524
rect 41468 13580 41524 13636
rect 41580 13356 41636 13412
rect 40796 11228 40852 11284
rect 41468 11228 41524 11284
rect 39452 10610 39508 10612
rect 39452 10558 39454 10610
rect 39454 10558 39506 10610
rect 39506 10558 39508 10610
rect 39452 10556 39508 10558
rect 40236 11004 40292 11060
rect 41916 13858 41972 13860
rect 41916 13806 41918 13858
rect 41918 13806 41970 13858
rect 41970 13806 41972 13858
rect 41916 13804 41972 13806
rect 41692 11004 41748 11060
rect 41804 13746 41860 13748
rect 41804 13694 41806 13746
rect 41806 13694 41858 13746
rect 41858 13694 41860 13746
rect 41804 13692 41860 13694
rect 42476 15820 42532 15876
rect 42364 15708 42420 15764
rect 42476 15372 42532 15428
rect 42476 15148 42532 15204
rect 42476 15036 42532 15092
rect 42924 16268 42980 16324
rect 42812 15874 42868 15876
rect 42812 15822 42814 15874
rect 42814 15822 42866 15874
rect 42866 15822 42868 15874
rect 42812 15820 42868 15822
rect 42812 15426 42868 15428
rect 42812 15374 42814 15426
rect 42814 15374 42866 15426
rect 42866 15374 42868 15426
rect 42812 15372 42868 15374
rect 42700 15148 42756 15204
rect 43260 16322 43316 16324
rect 43260 16270 43262 16322
rect 43262 16270 43314 16322
rect 43314 16270 43316 16322
rect 43260 16268 43316 16270
rect 43260 15596 43316 15652
rect 44156 18060 44212 18116
rect 44380 17890 44436 17892
rect 44380 17838 44382 17890
rect 44382 17838 44434 17890
rect 44434 17838 44436 17890
rect 44380 17836 44436 17838
rect 43932 17276 43988 17332
rect 44380 17500 44436 17556
rect 43708 16828 43764 16884
rect 43596 16156 43652 16212
rect 43484 16098 43540 16100
rect 43484 16046 43486 16098
rect 43486 16046 43538 16098
rect 43538 16046 43540 16098
rect 43484 16044 43540 16046
rect 43708 15596 43764 15652
rect 43596 15372 43652 15428
rect 43260 14700 43316 14756
rect 42028 13020 42084 13076
rect 42476 13692 42532 13748
rect 42140 12908 42196 12964
rect 42252 13580 42308 13636
rect 41916 12684 41972 12740
rect 42364 12124 42420 12180
rect 41916 11116 41972 11172
rect 42028 11004 42084 11060
rect 42028 10780 42084 10836
rect 40236 10610 40292 10612
rect 40236 10558 40238 10610
rect 40238 10558 40290 10610
rect 40290 10558 40292 10610
rect 40236 10556 40292 10558
rect 39116 9772 39172 9828
rect 38668 9548 38724 9604
rect 38220 9042 38276 9044
rect 38220 8990 38222 9042
rect 38222 8990 38274 9042
rect 38274 8990 38276 9042
rect 38220 8988 38276 8990
rect 37772 8876 37828 8932
rect 37772 8428 37828 8484
rect 37884 8034 37940 8036
rect 37884 7982 37886 8034
rect 37886 7982 37938 8034
rect 37938 7982 37940 8034
rect 37884 7980 37940 7982
rect 38332 7980 38388 8036
rect 38444 8092 38500 8148
rect 37660 7532 37716 7588
rect 36876 4284 36932 4340
rect 36876 3612 36932 3668
rect 37100 6524 37156 6580
rect 37100 5740 37156 5796
rect 37212 5180 37268 5236
rect 37324 5852 37380 5908
rect 37884 7308 37940 7364
rect 38332 6748 38388 6804
rect 37772 5122 37828 5124
rect 37772 5070 37774 5122
rect 37774 5070 37826 5122
rect 37826 5070 37828 5122
rect 37772 5068 37828 5070
rect 37436 4562 37492 4564
rect 37436 4510 37438 4562
rect 37438 4510 37490 4562
rect 37490 4510 37492 4562
rect 37436 4508 37492 4510
rect 37548 4396 37604 4452
rect 37996 6636 38052 6692
rect 40012 9826 40068 9828
rect 40012 9774 40014 9826
rect 40014 9774 40066 9826
rect 40066 9774 40068 9826
rect 40012 9772 40068 9774
rect 39340 9602 39396 9604
rect 39340 9550 39342 9602
rect 39342 9550 39394 9602
rect 39394 9550 39396 9602
rect 39340 9548 39396 9550
rect 39900 9436 39956 9492
rect 40348 9660 40404 9716
rect 38668 8876 38724 8932
rect 39004 8258 39060 8260
rect 39004 8206 39006 8258
rect 39006 8206 39058 8258
rect 39058 8206 39060 8258
rect 39004 8204 39060 8206
rect 38780 8146 38836 8148
rect 38780 8094 38782 8146
rect 38782 8094 38834 8146
rect 38834 8094 38836 8146
rect 38780 8092 38836 8094
rect 40348 9266 40404 9268
rect 40348 9214 40350 9266
rect 40350 9214 40402 9266
rect 40402 9214 40404 9266
rect 40348 9212 40404 9214
rect 39340 9154 39396 9156
rect 39340 9102 39342 9154
rect 39342 9102 39394 9154
rect 39394 9102 39396 9154
rect 39340 9100 39396 9102
rect 39452 9042 39508 9044
rect 39452 8990 39454 9042
rect 39454 8990 39506 9042
rect 39506 8990 39508 9042
rect 39452 8988 39508 8990
rect 39228 8370 39284 8372
rect 39228 8318 39230 8370
rect 39230 8318 39282 8370
rect 39282 8318 39284 8370
rect 39228 8316 39284 8318
rect 39676 8316 39732 8372
rect 41468 9826 41524 9828
rect 41468 9774 41470 9826
rect 41470 9774 41522 9826
rect 41522 9774 41524 9826
rect 41468 9772 41524 9774
rect 40908 9266 40964 9268
rect 40908 9214 40910 9266
rect 40910 9214 40962 9266
rect 40962 9214 40964 9266
rect 40908 9212 40964 9214
rect 40796 8316 40852 8372
rect 39452 8204 39508 8260
rect 41132 8258 41188 8260
rect 41132 8206 41134 8258
rect 41134 8206 41186 8258
rect 41186 8206 41188 8258
rect 41132 8204 41188 8206
rect 41692 9772 41748 9828
rect 39900 8092 39956 8148
rect 41580 7756 41636 7812
rect 41468 7644 41524 7700
rect 39900 6972 39956 7028
rect 38556 6636 38612 6692
rect 38780 6690 38836 6692
rect 38780 6638 38782 6690
rect 38782 6638 38834 6690
rect 38834 6638 38836 6690
rect 38780 6636 38836 6638
rect 38220 5180 38276 5236
rect 38444 4956 38500 5012
rect 37996 4284 38052 4340
rect 38780 4562 38836 4564
rect 38780 4510 38782 4562
rect 38782 4510 38834 4562
rect 38834 4510 38836 4562
rect 38780 4508 38836 4510
rect 40908 6018 40964 6020
rect 40908 5966 40910 6018
rect 40910 5966 40962 6018
rect 40962 5966 40964 6018
rect 40908 5964 40964 5966
rect 40124 4508 40180 4564
rect 41132 4508 41188 4564
rect 39340 4450 39396 4452
rect 39340 4398 39342 4450
rect 39342 4398 39394 4450
rect 39394 4398 39396 4450
rect 39340 4396 39396 4398
rect 39452 4284 39508 4340
rect 40012 4338 40068 4340
rect 40012 4286 40014 4338
rect 40014 4286 40066 4338
rect 40066 4286 40068 4338
rect 40012 4284 40068 4286
rect 40012 3554 40068 3556
rect 40012 3502 40014 3554
rect 40014 3502 40066 3554
rect 40066 3502 40068 3554
rect 40012 3500 40068 3502
rect 40908 3554 40964 3556
rect 40908 3502 40910 3554
rect 40910 3502 40962 3554
rect 40962 3502 40964 3554
rect 40908 3500 40964 3502
rect 42364 10780 42420 10836
rect 43148 14530 43204 14532
rect 43148 14478 43150 14530
rect 43150 14478 43202 14530
rect 43202 14478 43204 14530
rect 43148 14476 43204 14478
rect 42924 13916 42980 13972
rect 43260 13916 43316 13972
rect 42812 13804 42868 13860
rect 42700 13580 42756 13636
rect 42924 13692 42980 13748
rect 42924 13468 42980 13524
rect 42924 13020 42980 13076
rect 42700 12460 42756 12516
rect 42700 12066 42756 12068
rect 42700 12014 42702 12066
rect 42702 12014 42754 12066
rect 42754 12014 42756 12066
rect 42700 12012 42756 12014
rect 42924 11228 42980 11284
rect 43484 13692 43540 13748
rect 43484 13244 43540 13300
rect 43148 11618 43204 11620
rect 43148 11566 43150 11618
rect 43150 11566 43202 11618
rect 43202 11566 43204 11618
rect 43148 11564 43204 11566
rect 43260 11506 43316 11508
rect 43260 11454 43262 11506
rect 43262 11454 43314 11506
rect 43314 11454 43316 11506
rect 43260 11452 43316 11454
rect 43820 14924 43876 14980
rect 43708 13746 43764 13748
rect 43708 13694 43710 13746
rect 43710 13694 43762 13746
rect 43762 13694 43764 13746
rect 43708 13692 43764 13694
rect 44156 16268 44212 16324
rect 44828 18508 44884 18564
rect 44716 18284 44772 18340
rect 44828 17500 44884 17556
rect 44716 16994 44772 16996
rect 44716 16942 44718 16994
rect 44718 16942 44770 16994
rect 44770 16942 44772 16994
rect 44716 16940 44772 16942
rect 44156 15986 44212 15988
rect 44156 15934 44158 15986
rect 44158 15934 44210 15986
rect 44210 15934 44212 15986
rect 44156 15932 44212 15934
rect 44268 15596 44324 15652
rect 44268 15148 44324 15204
rect 44604 15426 44660 15428
rect 44604 15374 44606 15426
rect 44606 15374 44658 15426
rect 44658 15374 44660 15426
rect 44604 15372 44660 15374
rect 44044 14924 44100 14980
rect 43932 13970 43988 13972
rect 43932 13918 43934 13970
rect 43934 13918 43986 13970
rect 43986 13918 43988 13970
rect 43932 13916 43988 13918
rect 43932 13580 43988 13636
rect 44268 14418 44324 14420
rect 44268 14366 44270 14418
rect 44270 14366 44322 14418
rect 44322 14366 44324 14418
rect 44268 14364 44324 14366
rect 44268 13804 44324 13860
rect 44492 14140 44548 14196
rect 44604 14924 44660 14980
rect 44156 13244 44212 13300
rect 44156 12796 44212 12852
rect 44380 12796 44436 12852
rect 43596 11228 43652 11284
rect 43148 9996 43204 10052
rect 41916 9938 41972 9940
rect 41916 9886 41918 9938
rect 41918 9886 41970 9938
rect 41970 9886 41972 9938
rect 41916 9884 41972 9886
rect 42812 9826 42868 9828
rect 42812 9774 42814 9826
rect 42814 9774 42866 9826
rect 42866 9774 42868 9826
rect 42812 9772 42868 9774
rect 42476 9714 42532 9716
rect 42476 9662 42478 9714
rect 42478 9662 42530 9714
rect 42530 9662 42532 9714
rect 42476 9660 42532 9662
rect 42140 9212 42196 9268
rect 42476 9324 42532 9380
rect 42028 8428 42084 8484
rect 42364 8428 42420 8484
rect 41916 8204 41972 8260
rect 42924 9324 42980 9380
rect 42924 8764 42980 8820
rect 42924 8482 42980 8484
rect 42924 8430 42926 8482
rect 42926 8430 42978 8482
rect 42978 8430 42980 8482
rect 42924 8428 42980 8430
rect 42588 8316 42644 8372
rect 42476 7698 42532 7700
rect 42476 7646 42478 7698
rect 42478 7646 42530 7698
rect 42530 7646 42532 7698
rect 42476 7644 42532 7646
rect 42700 8258 42756 8260
rect 42700 8206 42702 8258
rect 42702 8206 42754 8258
rect 42754 8206 42756 8258
rect 42700 8204 42756 8206
rect 42700 7756 42756 7812
rect 43148 8876 43204 8932
rect 43260 8764 43316 8820
rect 43372 7644 43428 7700
rect 44492 12236 44548 12292
rect 45612 27916 45668 27972
rect 45612 27468 45668 27524
rect 46620 29426 46676 29428
rect 46620 29374 46622 29426
rect 46622 29374 46674 29426
rect 46674 29374 46676 29426
rect 46620 29372 46676 29374
rect 46620 28812 46676 28868
rect 47628 29986 47684 29988
rect 47628 29934 47630 29986
rect 47630 29934 47682 29986
rect 47682 29934 47684 29986
rect 47628 29932 47684 29934
rect 47404 29650 47460 29652
rect 47404 29598 47406 29650
rect 47406 29598 47458 29650
rect 47458 29598 47460 29650
rect 47404 29596 47460 29598
rect 47292 29484 47348 29540
rect 47180 29260 47236 29316
rect 47740 28812 47796 28868
rect 47964 29372 48020 29428
rect 45836 26850 45892 26852
rect 45836 26798 45838 26850
rect 45838 26798 45890 26850
rect 45890 26798 45892 26850
rect 45836 26796 45892 26798
rect 45836 26124 45892 26180
rect 45500 25452 45556 25508
rect 45500 25228 45556 25284
rect 45388 24108 45444 24164
rect 45388 23714 45444 23716
rect 45388 23662 45390 23714
rect 45390 23662 45442 23714
rect 45442 23662 45444 23714
rect 45388 23660 45444 23662
rect 45724 24444 45780 24500
rect 45612 23660 45668 23716
rect 45724 23772 45780 23828
rect 45500 23212 45556 23268
rect 45500 23042 45556 23044
rect 45500 22990 45502 23042
rect 45502 22990 45554 23042
rect 45554 22990 45556 23042
rect 45500 22988 45556 22990
rect 45612 22876 45668 22932
rect 45388 22258 45444 22260
rect 45388 22206 45390 22258
rect 45390 22206 45442 22258
rect 45442 22206 45444 22258
rect 45388 22204 45444 22206
rect 45500 21756 45556 21812
rect 45388 21698 45444 21700
rect 45388 21646 45390 21698
rect 45390 21646 45442 21698
rect 45442 21646 45444 21698
rect 45388 21644 45444 21646
rect 45388 21084 45444 21140
rect 45500 20242 45556 20244
rect 45500 20190 45502 20242
rect 45502 20190 45554 20242
rect 45554 20190 45556 20242
rect 45500 20188 45556 20190
rect 45276 19516 45332 19572
rect 45164 19292 45220 19348
rect 45276 19180 45332 19236
rect 45500 20018 45556 20020
rect 45500 19966 45502 20018
rect 45502 19966 45554 20018
rect 45554 19966 45556 20018
rect 45500 19964 45556 19966
rect 45612 19852 45668 19908
rect 45164 17500 45220 17556
rect 45388 17052 45444 17108
rect 45612 18732 45668 18788
rect 45948 24780 46004 24836
rect 46956 27804 47012 27860
rect 47068 28028 47124 28084
rect 46844 27692 46900 27748
rect 46956 27634 47012 27636
rect 46956 27582 46958 27634
rect 46958 27582 47010 27634
rect 47010 27582 47012 27634
rect 46956 27580 47012 27582
rect 46396 26908 46452 26964
rect 46172 26012 46228 26068
rect 45948 24610 46004 24612
rect 45948 24558 45950 24610
rect 45950 24558 46002 24610
rect 46002 24558 46004 24610
rect 45948 24556 46004 24558
rect 45836 23436 45892 23492
rect 45948 23772 46004 23828
rect 45836 23212 45892 23268
rect 46284 23436 46340 23492
rect 46620 27468 46676 27524
rect 46508 26684 46564 26740
rect 47628 27858 47684 27860
rect 47628 27806 47630 27858
rect 47630 27806 47682 27858
rect 47682 27806 47684 27858
rect 47628 27804 47684 27806
rect 47180 27692 47236 27748
rect 47628 27580 47684 27636
rect 47516 27468 47572 27524
rect 47068 26290 47124 26292
rect 47068 26238 47070 26290
rect 47070 26238 47122 26290
rect 47122 26238 47124 26290
rect 47068 26236 47124 26238
rect 46844 26012 46900 26068
rect 46732 25282 46788 25284
rect 46732 25230 46734 25282
rect 46734 25230 46786 25282
rect 46786 25230 46788 25282
rect 46732 25228 46788 25230
rect 47404 25340 47460 25396
rect 47740 26962 47796 26964
rect 47740 26910 47742 26962
rect 47742 26910 47794 26962
rect 47794 26910 47796 26962
rect 47740 26908 47796 26910
rect 47628 25394 47684 25396
rect 47628 25342 47630 25394
rect 47630 25342 47682 25394
rect 47682 25342 47684 25394
rect 47628 25340 47684 25342
rect 47740 25506 47796 25508
rect 47740 25454 47742 25506
rect 47742 25454 47794 25506
rect 47794 25454 47796 25506
rect 47740 25452 47796 25454
rect 46956 25228 47012 25284
rect 47964 27970 48020 27972
rect 47964 27918 47966 27970
rect 47966 27918 48018 27970
rect 48018 27918 48020 27970
rect 47964 27916 48020 27918
rect 48636 31500 48692 31556
rect 49084 31554 49140 31556
rect 49084 31502 49086 31554
rect 49086 31502 49138 31554
rect 49138 31502 49140 31554
rect 49084 31500 49140 31502
rect 50204 31554 50260 31556
rect 50204 31502 50206 31554
rect 50206 31502 50258 31554
rect 50258 31502 50260 31554
rect 50204 31500 50260 31502
rect 49532 31106 49588 31108
rect 49532 31054 49534 31106
rect 49534 31054 49586 31106
rect 49586 31054 49588 31106
rect 49532 31052 49588 31054
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50652 31218 50708 31220
rect 50652 31166 50654 31218
rect 50654 31166 50706 31218
rect 50706 31166 50708 31218
rect 50652 31164 50708 31166
rect 50428 30994 50484 30996
rect 50428 30942 50430 30994
rect 50430 30942 50482 30994
rect 50482 30942 50484 30994
rect 50428 30940 50484 30942
rect 48188 29314 48244 29316
rect 48188 29262 48190 29314
rect 48190 29262 48242 29314
rect 48242 29262 48244 29314
rect 48188 29260 48244 29262
rect 48188 28476 48244 28532
rect 48524 29932 48580 29988
rect 48524 28812 48580 28868
rect 48412 28754 48468 28756
rect 48412 28702 48414 28754
rect 48414 28702 48466 28754
rect 48466 28702 48468 28754
rect 48412 28700 48468 28702
rect 49756 30156 49812 30212
rect 49308 30098 49364 30100
rect 49308 30046 49310 30098
rect 49310 30046 49362 30098
rect 49362 30046 49364 30098
rect 49308 30044 49364 30046
rect 49644 30098 49700 30100
rect 49644 30046 49646 30098
rect 49646 30046 49698 30098
rect 49698 30046 49700 30098
rect 49644 30044 49700 30046
rect 48748 29596 48804 29652
rect 49644 29650 49700 29652
rect 49644 29598 49646 29650
rect 49646 29598 49698 29650
rect 49698 29598 49700 29650
rect 49644 29596 49700 29598
rect 50652 30492 50708 30548
rect 50204 30098 50260 30100
rect 50204 30046 50206 30098
rect 50206 30046 50258 30098
rect 50258 30046 50260 30098
rect 50204 30044 50260 30046
rect 50876 29932 50932 29988
rect 50988 30156 51044 30212
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50428 29596 50484 29652
rect 50204 29484 50260 29540
rect 48636 28028 48692 28084
rect 48300 27804 48356 27860
rect 48524 27804 48580 27860
rect 48188 27186 48244 27188
rect 48188 27134 48190 27186
rect 48190 27134 48242 27186
rect 48242 27134 48244 27186
rect 48188 27132 48244 27134
rect 47964 27020 48020 27076
rect 48076 26796 48132 26852
rect 48636 27746 48692 27748
rect 48636 27694 48638 27746
rect 48638 27694 48690 27746
rect 48690 27694 48692 27746
rect 48636 27692 48692 27694
rect 48860 27916 48916 27972
rect 48972 29260 49028 29316
rect 48300 26012 48356 26068
rect 48188 25282 48244 25284
rect 48188 25230 48190 25282
rect 48190 25230 48242 25282
rect 48242 25230 48244 25282
rect 48188 25228 48244 25230
rect 48076 25116 48132 25172
rect 46956 24834 47012 24836
rect 46956 24782 46958 24834
rect 46958 24782 47010 24834
rect 47010 24782 47012 24834
rect 46956 24780 47012 24782
rect 47180 24834 47236 24836
rect 47180 24782 47182 24834
rect 47182 24782 47234 24834
rect 47234 24782 47236 24834
rect 47180 24780 47236 24782
rect 47292 24668 47348 24724
rect 46620 23996 46676 24052
rect 46620 23714 46676 23716
rect 46620 23662 46622 23714
rect 46622 23662 46674 23714
rect 46674 23662 46676 23714
rect 46620 23660 46676 23662
rect 46396 23212 46452 23268
rect 46508 23436 46564 23492
rect 46172 22988 46228 23044
rect 46060 22316 46116 22372
rect 46396 22876 46452 22932
rect 45948 22146 46004 22148
rect 45948 22094 45950 22146
rect 45950 22094 46002 22146
rect 46002 22094 46004 22146
rect 45948 22092 46004 22094
rect 45948 21698 46004 21700
rect 45948 21646 45950 21698
rect 45950 21646 46002 21698
rect 46002 21646 46004 21698
rect 45948 21644 46004 21646
rect 45948 19122 46004 19124
rect 45948 19070 45950 19122
rect 45950 19070 46002 19122
rect 46002 19070 46004 19122
rect 45948 19068 46004 19070
rect 46956 23938 47012 23940
rect 46956 23886 46958 23938
rect 46958 23886 47010 23938
rect 47010 23886 47012 23938
rect 46956 23884 47012 23886
rect 46844 23436 46900 23492
rect 46844 22764 46900 22820
rect 46732 22316 46788 22372
rect 47180 23826 47236 23828
rect 47180 23774 47182 23826
rect 47182 23774 47234 23826
rect 47234 23774 47236 23826
rect 47180 23772 47236 23774
rect 47292 23660 47348 23716
rect 47180 23212 47236 23268
rect 46956 22204 47012 22260
rect 46172 21644 46228 21700
rect 47852 24780 47908 24836
rect 47628 24610 47684 24612
rect 47628 24558 47630 24610
rect 47630 24558 47682 24610
rect 47682 24558 47684 24610
rect 47628 24556 47684 24558
rect 47516 24220 47572 24276
rect 47740 24444 47796 24500
rect 47740 23378 47796 23380
rect 47740 23326 47742 23378
rect 47742 23326 47794 23378
rect 47794 23326 47796 23378
rect 47740 23324 47796 23326
rect 47180 22764 47236 22820
rect 46732 21756 46788 21812
rect 46284 20802 46340 20804
rect 46284 20750 46286 20802
rect 46286 20750 46338 20802
rect 46338 20750 46340 20802
rect 46284 20748 46340 20750
rect 46844 21084 46900 21140
rect 46396 19964 46452 20020
rect 46172 19852 46228 19908
rect 46284 19628 46340 19684
rect 46732 20802 46788 20804
rect 46732 20750 46734 20802
rect 46734 20750 46786 20802
rect 46786 20750 46788 20802
rect 46732 20748 46788 20750
rect 46620 19964 46676 20020
rect 46732 20300 46788 20356
rect 46396 19292 46452 19348
rect 46172 19180 46228 19236
rect 45836 18396 45892 18452
rect 45724 18172 45780 18228
rect 45836 17106 45892 17108
rect 45836 17054 45838 17106
rect 45838 17054 45890 17106
rect 45890 17054 45892 17106
rect 45836 17052 45892 17054
rect 45500 16716 45556 16772
rect 45052 15596 45108 15652
rect 45276 15932 45332 15988
rect 44828 14476 44884 14532
rect 44716 12572 44772 12628
rect 44492 11788 44548 11844
rect 44156 11618 44212 11620
rect 44156 11566 44158 11618
rect 44158 11566 44210 11618
rect 44210 11566 44212 11618
rect 44156 11564 44212 11566
rect 44268 11676 44324 11732
rect 44044 11340 44100 11396
rect 43932 11228 43988 11284
rect 44380 11618 44436 11620
rect 44380 11566 44382 11618
rect 44382 11566 44434 11618
rect 44434 11566 44436 11618
rect 44380 11564 44436 11566
rect 44268 11004 44324 11060
rect 45164 14140 45220 14196
rect 45724 16828 45780 16884
rect 45836 16044 45892 16100
rect 45724 15036 45780 15092
rect 45500 14418 45556 14420
rect 45500 14366 45502 14418
rect 45502 14366 45554 14418
rect 45554 14366 45556 14418
rect 45500 14364 45556 14366
rect 45724 14364 45780 14420
rect 46060 17724 46116 17780
rect 46172 17612 46228 17668
rect 46060 16828 46116 16884
rect 46172 16492 46228 16548
rect 46620 18396 46676 18452
rect 46732 18284 46788 18340
rect 46620 17612 46676 17668
rect 46956 16492 47012 16548
rect 46396 15820 46452 15876
rect 46172 15314 46228 15316
rect 46172 15262 46174 15314
rect 46174 15262 46226 15314
rect 46226 15262 46228 15314
rect 46172 15260 46228 15262
rect 45388 14252 45444 14308
rect 45500 14140 45556 14196
rect 47068 19628 47124 19684
rect 47516 22652 47572 22708
rect 47516 22428 47572 22484
rect 47404 22092 47460 22148
rect 48748 26908 48804 26964
rect 48860 26684 48916 26740
rect 48748 25676 48804 25732
rect 48636 25564 48692 25620
rect 47964 23996 48020 24052
rect 48412 25228 48468 25284
rect 48636 25116 48692 25172
rect 48524 24108 48580 24164
rect 48748 24108 48804 24164
rect 49308 28476 49364 28532
rect 49308 27356 49364 27412
rect 49084 27074 49140 27076
rect 49084 27022 49086 27074
rect 49086 27022 49138 27074
rect 49138 27022 49140 27074
rect 49084 27020 49140 27022
rect 49756 29148 49812 29204
rect 49756 28700 49812 28756
rect 49644 28140 49700 28196
rect 50316 29372 50372 29428
rect 50428 29148 50484 29204
rect 50428 28754 50484 28756
rect 50428 28702 50430 28754
rect 50430 28702 50482 28754
rect 50482 28702 50484 28754
rect 50428 28700 50484 28702
rect 50652 28476 50708 28532
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50876 28028 50932 28084
rect 49532 27692 49588 27748
rect 50876 27244 50932 27300
rect 49196 26962 49252 26964
rect 49196 26910 49198 26962
rect 49198 26910 49250 26962
rect 49250 26910 49252 26962
rect 49196 26908 49252 26910
rect 49196 26684 49252 26740
rect 49532 26460 49588 26516
rect 49420 26012 49476 26068
rect 49308 25452 49364 25508
rect 49868 26178 49924 26180
rect 49868 26126 49870 26178
rect 49870 26126 49922 26178
rect 49922 26126 49924 26178
rect 49868 26124 49924 26126
rect 49532 25452 49588 25508
rect 49084 23996 49140 24052
rect 48300 23436 48356 23492
rect 48188 23042 48244 23044
rect 48188 22990 48190 23042
rect 48190 22990 48242 23042
rect 48242 22990 48244 23042
rect 48188 22988 48244 22990
rect 48188 22258 48244 22260
rect 48188 22206 48190 22258
rect 48190 22206 48242 22258
rect 48242 22206 48244 22258
rect 48188 22204 48244 22206
rect 48300 22092 48356 22148
rect 48076 21756 48132 21812
rect 48972 23436 49028 23492
rect 49196 23324 49252 23380
rect 49420 25228 49476 25284
rect 49084 22988 49140 23044
rect 48860 22876 48916 22932
rect 49196 22876 49252 22932
rect 49196 22540 49252 22596
rect 47964 21308 48020 21364
rect 48300 21196 48356 21252
rect 47516 20076 47572 20132
rect 47292 19404 47348 19460
rect 47180 16322 47236 16324
rect 47180 16270 47182 16322
rect 47182 16270 47234 16322
rect 47234 16270 47236 16322
rect 47180 16268 47236 16270
rect 47404 17666 47460 17668
rect 47404 17614 47406 17666
rect 47406 17614 47458 17666
rect 47458 17614 47460 17666
rect 47404 17612 47460 17614
rect 47628 19068 47684 19124
rect 47516 17276 47572 17332
rect 47404 16716 47460 16772
rect 47516 16604 47572 16660
rect 46956 15820 47012 15876
rect 46956 15596 47012 15652
rect 47404 15596 47460 15652
rect 47180 15314 47236 15316
rect 47180 15262 47182 15314
rect 47182 15262 47234 15314
rect 47234 15262 47236 15314
rect 47180 15260 47236 15262
rect 46172 14252 46228 14308
rect 45724 13468 45780 13524
rect 45948 13074 46004 13076
rect 45948 13022 45950 13074
rect 45950 13022 46002 13074
rect 46002 13022 46004 13074
rect 45948 13020 46004 13022
rect 45164 12460 45220 12516
rect 45276 12572 45332 12628
rect 45836 12796 45892 12852
rect 45164 11788 45220 11844
rect 44940 11564 44996 11620
rect 45052 11676 45108 11732
rect 45276 11228 45332 11284
rect 44492 10220 44548 10276
rect 43820 9212 43876 9268
rect 43820 8876 43876 8932
rect 44716 10050 44772 10052
rect 44716 9998 44718 10050
rect 44718 9998 44770 10050
rect 44770 9998 44772 10050
rect 44716 9996 44772 9998
rect 43484 8204 43540 8260
rect 44044 8258 44100 8260
rect 44044 8206 44046 8258
rect 44046 8206 44098 8258
rect 44098 8206 44100 8258
rect 44044 8204 44100 8206
rect 44380 7868 44436 7924
rect 43820 7756 43876 7812
rect 44380 7698 44436 7700
rect 44380 7646 44382 7698
rect 44382 7646 44434 7698
rect 44434 7646 44436 7698
rect 44380 7644 44436 7646
rect 43596 6690 43652 6692
rect 43596 6638 43598 6690
rect 43598 6638 43650 6690
rect 43650 6638 43652 6690
rect 43596 6636 43652 6638
rect 45164 9884 45220 9940
rect 44492 6636 44548 6692
rect 44604 6972 44660 7028
rect 42588 6300 42644 6356
rect 42812 6018 42868 6020
rect 42812 5966 42814 6018
rect 42814 5966 42866 6018
rect 42866 5966 42868 6018
rect 42812 5964 42868 5966
rect 43036 5740 43092 5796
rect 43484 5740 43540 5796
rect 41916 5122 41972 5124
rect 41916 5070 41918 5122
rect 41918 5070 41970 5122
rect 41970 5070 41972 5122
rect 41916 5068 41972 5070
rect 42588 5068 42644 5124
rect 44044 6300 44100 6356
rect 43820 6018 43876 6020
rect 43820 5966 43822 6018
rect 43822 5966 43874 6018
rect 43874 5966 43876 6018
rect 43820 5964 43876 5966
rect 44380 6188 44436 6244
rect 45388 11116 45444 11172
rect 45724 11676 45780 11732
rect 45836 11788 45892 11844
rect 45948 12012 46004 12068
rect 45724 11004 45780 11060
rect 45724 10668 45780 10724
rect 45724 9100 45780 9156
rect 46172 13580 46228 13636
rect 46732 14306 46788 14308
rect 46732 14254 46734 14306
rect 46734 14254 46786 14306
rect 46786 14254 46788 14306
rect 46732 14252 46788 14254
rect 46172 12290 46228 12292
rect 46172 12238 46174 12290
rect 46174 12238 46226 12290
rect 46226 12238 46228 12290
rect 46172 12236 46228 12238
rect 46284 11788 46340 11844
rect 46060 10834 46116 10836
rect 46060 10782 46062 10834
rect 46062 10782 46114 10834
rect 46114 10782 46116 10834
rect 46060 10780 46116 10782
rect 45836 9996 45892 10052
rect 45500 7756 45556 7812
rect 45388 6412 45444 6468
rect 45276 6300 45332 6356
rect 44380 6018 44436 6020
rect 44380 5966 44382 6018
rect 44382 5966 44434 6018
rect 44434 5966 44436 6018
rect 44380 5964 44436 5966
rect 45388 6130 45444 6132
rect 45388 6078 45390 6130
rect 45390 6078 45442 6130
rect 45442 6078 45444 6130
rect 45388 6076 45444 6078
rect 45948 10668 46004 10724
rect 46508 14028 46564 14084
rect 46732 13858 46788 13860
rect 46732 13806 46734 13858
rect 46734 13806 46786 13858
rect 46786 13806 46788 13858
rect 46732 13804 46788 13806
rect 46508 13746 46564 13748
rect 46508 13694 46510 13746
rect 46510 13694 46562 13746
rect 46562 13694 46564 13746
rect 46508 13692 46564 13694
rect 46732 13468 46788 13524
rect 46508 12962 46564 12964
rect 46508 12910 46510 12962
rect 46510 12910 46562 12962
rect 46562 12910 46564 12962
rect 46508 12908 46564 12910
rect 47068 14418 47124 14420
rect 47068 14366 47070 14418
rect 47070 14366 47122 14418
rect 47122 14366 47124 14418
rect 47068 14364 47124 14366
rect 47180 14252 47236 14308
rect 46956 13804 47012 13860
rect 47068 14140 47124 14196
rect 46508 12012 46564 12068
rect 47516 15372 47572 15428
rect 47404 15148 47460 15204
rect 48188 20018 48244 20020
rect 48188 19966 48190 20018
rect 48190 19966 48242 20018
rect 48242 19966 48244 20018
rect 48188 19964 48244 19966
rect 48412 19740 48468 19796
rect 48076 19516 48132 19572
rect 50428 26962 50484 26964
rect 50428 26910 50430 26962
rect 50430 26910 50482 26962
rect 50482 26910 50484 26962
rect 50428 26908 50484 26910
rect 51996 32396 52052 32452
rect 52668 32674 52724 32676
rect 52668 32622 52670 32674
rect 52670 32622 52722 32674
rect 52722 32622 52724 32674
rect 52668 32620 52724 32622
rect 52444 31778 52500 31780
rect 52444 31726 52446 31778
rect 52446 31726 52498 31778
rect 52498 31726 52500 31778
rect 52444 31724 52500 31726
rect 52108 30828 52164 30884
rect 52332 30770 52388 30772
rect 52332 30718 52334 30770
rect 52334 30718 52386 30770
rect 52386 30718 52388 30770
rect 52332 30716 52388 30718
rect 51324 30156 51380 30212
rect 51436 30268 51492 30324
rect 51212 29820 51268 29876
rect 51100 29484 51156 29540
rect 51212 29596 51268 29652
rect 51324 29036 51380 29092
rect 51212 28812 51268 28868
rect 51548 29260 51604 29316
rect 51772 29820 51828 29876
rect 51772 29260 51828 29316
rect 51884 29484 51940 29540
rect 52108 29148 52164 29204
rect 51884 28588 51940 28644
rect 51660 28530 51716 28532
rect 51660 28478 51662 28530
rect 51662 28478 51714 28530
rect 51714 28478 51716 28530
rect 51660 28476 51716 28478
rect 51212 28028 51268 28084
rect 51212 27020 51268 27076
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50204 26124 50260 26180
rect 50988 26178 51044 26180
rect 50988 26126 50990 26178
rect 50990 26126 51042 26178
rect 51042 26126 51044 26178
rect 50988 26124 51044 26126
rect 50092 25282 50148 25284
rect 50092 25230 50094 25282
rect 50094 25230 50146 25282
rect 50146 25230 50148 25282
rect 50092 25228 50148 25230
rect 49980 24834 50036 24836
rect 49980 24782 49982 24834
rect 49982 24782 50034 24834
rect 50034 24782 50036 24834
rect 49980 24780 50036 24782
rect 49644 24498 49700 24500
rect 49644 24446 49646 24498
rect 49646 24446 49698 24498
rect 49698 24446 49700 24498
rect 49644 24444 49700 24446
rect 49756 24108 49812 24164
rect 49868 23996 49924 24052
rect 49532 23436 49588 23492
rect 49532 22540 49588 22596
rect 49420 22316 49476 22372
rect 49532 22146 49588 22148
rect 49532 22094 49534 22146
rect 49534 22094 49586 22146
rect 49586 22094 49588 22146
rect 49532 22092 49588 22094
rect 49756 22876 49812 22932
rect 50316 24668 50372 24724
rect 49868 22988 49924 23044
rect 49868 22428 49924 22484
rect 50204 24444 50260 24500
rect 50092 22988 50148 23044
rect 49980 22146 50036 22148
rect 49980 22094 49982 22146
rect 49982 22094 50034 22146
rect 50034 22094 50036 22146
rect 49980 22092 50036 22094
rect 49756 21980 49812 22036
rect 48972 21756 49028 21812
rect 49420 21756 49476 21812
rect 49756 21756 49812 21812
rect 48748 21586 48804 21588
rect 48748 21534 48750 21586
rect 48750 21534 48802 21586
rect 48802 21534 48804 21586
rect 48748 21532 48804 21534
rect 49532 21586 49588 21588
rect 49532 21534 49534 21586
rect 49534 21534 49586 21586
rect 49586 21534 49588 21586
rect 49532 21532 49588 21534
rect 48636 20972 48692 21028
rect 49532 21026 49588 21028
rect 49532 20974 49534 21026
rect 49534 20974 49586 21026
rect 49586 20974 49588 21026
rect 49532 20972 49588 20974
rect 49196 20748 49252 20804
rect 48636 20188 48692 20244
rect 48636 20018 48692 20020
rect 48636 19966 48638 20018
rect 48638 19966 48690 20018
rect 48690 19966 48692 20018
rect 48636 19964 48692 19966
rect 48524 19516 48580 19572
rect 48188 18732 48244 18788
rect 48412 18674 48468 18676
rect 48412 18622 48414 18674
rect 48414 18622 48466 18674
rect 48466 18622 48468 18674
rect 48412 18620 48468 18622
rect 48300 18562 48356 18564
rect 48300 18510 48302 18562
rect 48302 18510 48354 18562
rect 48354 18510 48356 18562
rect 48300 18508 48356 18510
rect 48300 18172 48356 18228
rect 48300 17276 48356 17332
rect 47852 16940 47908 16996
rect 47852 15820 47908 15876
rect 47964 16716 48020 16772
rect 49084 20578 49140 20580
rect 49084 20526 49086 20578
rect 49086 20526 49138 20578
rect 49138 20526 49140 20578
rect 49084 20524 49140 20526
rect 48860 20412 48916 20468
rect 48860 19740 48916 19796
rect 48972 19852 49028 19908
rect 49420 20802 49476 20804
rect 49420 20750 49422 20802
rect 49422 20750 49474 20802
rect 49474 20750 49476 20802
rect 49420 20748 49476 20750
rect 49756 20972 49812 21028
rect 49644 20412 49700 20468
rect 49420 19346 49476 19348
rect 49420 19294 49422 19346
rect 49422 19294 49474 19346
rect 49474 19294 49476 19346
rect 49420 19292 49476 19294
rect 49196 18956 49252 19012
rect 48860 18284 48916 18340
rect 48972 18396 49028 18452
rect 48748 17164 48804 17220
rect 48860 17836 48916 17892
rect 48300 16716 48356 16772
rect 48748 16770 48804 16772
rect 48748 16718 48750 16770
rect 48750 16718 48802 16770
rect 48802 16718 48804 16770
rect 48748 16716 48804 16718
rect 48188 16604 48244 16660
rect 48412 16268 48468 16324
rect 48300 16044 48356 16100
rect 47740 15036 47796 15092
rect 48076 15596 48132 15652
rect 47404 13916 47460 13972
rect 47740 14364 47796 14420
rect 47740 13916 47796 13972
rect 47404 13580 47460 13636
rect 47516 12460 47572 12516
rect 47068 12236 47124 12292
rect 46844 11676 46900 11732
rect 47516 12012 47572 12068
rect 46620 10892 46676 10948
rect 46508 9938 46564 9940
rect 46508 9886 46510 9938
rect 46510 9886 46562 9938
rect 46562 9886 46564 9938
rect 46508 9884 46564 9886
rect 47180 11340 47236 11396
rect 45724 7586 45780 7588
rect 45724 7534 45726 7586
rect 45726 7534 45778 7586
rect 45778 7534 45780 7586
rect 45724 7532 45780 7534
rect 45612 7084 45668 7140
rect 46396 7868 46452 7924
rect 46172 7308 46228 7364
rect 46060 6578 46116 6580
rect 46060 6526 46062 6578
rect 46062 6526 46114 6578
rect 46114 6526 46116 6578
rect 46060 6524 46116 6526
rect 45948 6188 46004 6244
rect 46732 8988 46788 9044
rect 46844 11116 46900 11172
rect 46844 8428 46900 8484
rect 47404 9548 47460 9604
rect 47964 14700 48020 14756
rect 47964 14140 48020 14196
rect 48524 15986 48580 15988
rect 48524 15934 48526 15986
rect 48526 15934 48578 15986
rect 48578 15934 48580 15986
rect 48524 15932 48580 15934
rect 48412 15426 48468 15428
rect 48412 15374 48414 15426
rect 48414 15374 48466 15426
rect 48466 15374 48468 15426
rect 48412 15372 48468 15374
rect 48188 14252 48244 14308
rect 48412 13746 48468 13748
rect 48412 13694 48414 13746
rect 48414 13694 48466 13746
rect 48466 13694 48468 13746
rect 48412 13692 48468 13694
rect 47852 11340 47908 11396
rect 48188 13580 48244 13636
rect 48076 12908 48132 12964
rect 48300 13468 48356 13524
rect 48188 12066 48244 12068
rect 48188 12014 48190 12066
rect 48190 12014 48242 12066
rect 48242 12014 48244 12066
rect 48188 12012 48244 12014
rect 48300 11506 48356 11508
rect 48300 11454 48302 11506
rect 48302 11454 48354 11506
rect 48354 11454 48356 11506
rect 48300 11452 48356 11454
rect 47852 9996 47908 10052
rect 47292 9266 47348 9268
rect 47292 9214 47294 9266
rect 47294 9214 47346 9266
rect 47346 9214 47348 9266
rect 47292 9212 47348 9214
rect 48748 15596 48804 15652
rect 48972 17164 49028 17220
rect 49420 17052 49476 17108
rect 49084 15596 49140 15652
rect 48860 14700 48916 14756
rect 48972 14924 49028 14980
rect 48972 14588 49028 14644
rect 48972 14140 49028 14196
rect 48748 11452 48804 11508
rect 48860 13804 48916 13860
rect 48748 11282 48804 11284
rect 48748 11230 48750 11282
rect 48750 11230 48802 11282
rect 48802 11230 48804 11282
rect 48748 11228 48804 11230
rect 48636 10108 48692 10164
rect 48188 9602 48244 9604
rect 48188 9550 48190 9602
rect 48190 9550 48242 9602
rect 48242 9550 48244 9602
rect 48188 9548 48244 9550
rect 47516 8876 47572 8932
rect 47068 8316 47124 8372
rect 47292 8428 47348 8484
rect 46844 8204 46900 8260
rect 46732 8146 46788 8148
rect 46732 8094 46734 8146
rect 46734 8094 46786 8146
rect 46786 8094 46788 8146
rect 46732 8092 46788 8094
rect 46620 7756 46676 7812
rect 46956 7868 47012 7924
rect 46844 7532 46900 7588
rect 47180 8034 47236 8036
rect 47180 7982 47182 8034
rect 47182 7982 47234 8034
rect 47234 7982 47236 8034
rect 47180 7980 47236 7982
rect 47068 7532 47124 7588
rect 46732 7308 46788 7364
rect 46620 6690 46676 6692
rect 46620 6638 46622 6690
rect 46622 6638 46674 6690
rect 46674 6638 46676 6690
rect 46620 6636 46676 6638
rect 47516 7698 47572 7700
rect 47516 7646 47518 7698
rect 47518 7646 47570 7698
rect 47570 7646 47572 7698
rect 47516 7644 47572 7646
rect 47516 6972 47572 7028
rect 47404 6524 47460 6580
rect 47404 5740 47460 5796
rect 46732 5234 46788 5236
rect 46732 5182 46734 5234
rect 46734 5182 46786 5234
rect 46786 5182 46788 5234
rect 46732 5180 46788 5182
rect 46844 5404 46900 5460
rect 43596 4956 43652 5012
rect 47740 8258 47796 8260
rect 47740 8206 47742 8258
rect 47742 8206 47794 8258
rect 47794 8206 47796 8258
rect 47740 8204 47796 8206
rect 47964 8876 48020 8932
rect 48076 8204 48132 8260
rect 47852 8092 47908 8148
rect 47852 7532 47908 7588
rect 47628 6636 47684 6692
rect 47964 7196 48020 7252
rect 48188 7698 48244 7700
rect 48188 7646 48190 7698
rect 48190 7646 48242 7698
rect 48242 7646 48244 7698
rect 48188 7644 48244 7646
rect 48076 6972 48132 7028
rect 48188 6690 48244 6692
rect 48188 6638 48190 6690
rect 48190 6638 48242 6690
rect 48242 6638 48244 6690
rect 48188 6636 48244 6638
rect 47628 5404 47684 5460
rect 48076 6188 48132 6244
rect 48188 6076 48244 6132
rect 48412 8316 48468 8372
rect 48524 9660 48580 9716
rect 48636 8428 48692 8484
rect 48524 6748 48580 6804
rect 48412 6524 48468 6580
rect 47964 5292 48020 5348
rect 48300 5404 48356 5460
rect 47852 5234 47908 5236
rect 47852 5182 47854 5234
rect 47854 5182 47906 5234
rect 47906 5182 47908 5234
rect 47852 5180 47908 5182
rect 49868 19740 49924 19796
rect 49868 19346 49924 19348
rect 49868 19294 49870 19346
rect 49870 19294 49922 19346
rect 49922 19294 49924 19346
rect 49868 19292 49924 19294
rect 50092 21586 50148 21588
rect 50092 21534 50094 21586
rect 50094 21534 50146 21586
rect 50146 21534 50148 21586
rect 50092 21532 50148 21534
rect 50092 20524 50148 20580
rect 49980 19068 50036 19124
rect 49980 18620 50036 18676
rect 49644 18450 49700 18452
rect 49644 18398 49646 18450
rect 49646 18398 49698 18450
rect 49698 18398 49700 18450
rect 49644 18396 49700 18398
rect 49644 17948 49700 18004
rect 49644 17666 49700 17668
rect 49644 17614 49646 17666
rect 49646 17614 49698 17666
rect 49698 17614 49700 17666
rect 49644 17612 49700 17614
rect 49756 17554 49812 17556
rect 49756 17502 49758 17554
rect 49758 17502 49810 17554
rect 49810 17502 49812 17554
rect 49756 17500 49812 17502
rect 49980 18172 50036 18228
rect 50876 25394 50932 25396
rect 50876 25342 50878 25394
rect 50878 25342 50930 25394
rect 50930 25342 50932 25394
rect 50876 25340 50932 25342
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 51772 28082 51828 28084
rect 51772 28030 51774 28082
rect 51774 28030 51826 28082
rect 51826 28030 51828 28082
rect 51772 28028 51828 28030
rect 51324 26348 51380 26404
rect 51996 29036 52052 29092
rect 51884 27132 51940 27188
rect 51324 25788 51380 25844
rect 51548 25788 51604 25844
rect 51548 25452 51604 25508
rect 51772 26348 51828 26404
rect 51772 26066 51828 26068
rect 51772 26014 51774 26066
rect 51774 26014 51826 26066
rect 51826 26014 51828 26066
rect 51772 26012 51828 26014
rect 51772 25340 51828 25396
rect 50764 24050 50820 24052
rect 50764 23998 50766 24050
rect 50766 23998 50818 24050
rect 50818 23998 50820 24050
rect 50764 23996 50820 23998
rect 50428 23714 50484 23716
rect 50428 23662 50430 23714
rect 50430 23662 50482 23714
rect 50482 23662 50484 23714
rect 50428 23660 50484 23662
rect 50988 23938 51044 23940
rect 50988 23886 50990 23938
rect 50990 23886 51042 23938
rect 51042 23886 51044 23938
rect 50988 23884 51044 23886
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50428 23324 50484 23380
rect 50652 23324 50708 23380
rect 50540 23042 50596 23044
rect 50540 22990 50542 23042
rect 50542 22990 50594 23042
rect 50594 22990 50596 23042
rect 50540 22988 50596 22990
rect 50988 23154 51044 23156
rect 50988 23102 50990 23154
rect 50990 23102 51042 23154
rect 51042 23102 51044 23154
rect 50988 23100 51044 23102
rect 50316 21084 50372 21140
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50988 21868 51044 21924
rect 50652 21756 50708 21812
rect 50540 21084 50596 21140
rect 50988 21586 51044 21588
rect 50988 21534 50990 21586
rect 50990 21534 51042 21586
rect 51042 21534 51044 21586
rect 50988 21532 51044 21534
rect 50316 20690 50372 20692
rect 50316 20638 50318 20690
rect 50318 20638 50370 20690
rect 50370 20638 50372 20690
rect 50316 20636 50372 20638
rect 50876 20578 50932 20580
rect 50876 20526 50878 20578
rect 50878 20526 50930 20578
rect 50930 20526 50932 20578
rect 50876 20524 50932 20526
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50988 20412 51044 20468
rect 50764 20356 50820 20358
rect 50764 20130 50820 20132
rect 50764 20078 50766 20130
rect 50766 20078 50818 20130
rect 50818 20078 50820 20130
rect 50764 20076 50820 20078
rect 51660 24892 51716 24948
rect 52108 28642 52164 28644
rect 52108 28590 52110 28642
rect 52110 28590 52162 28642
rect 52162 28590 52164 28642
rect 52108 28588 52164 28590
rect 52220 28476 52276 28532
rect 52332 27746 52388 27748
rect 52332 27694 52334 27746
rect 52334 27694 52386 27746
rect 52386 27694 52388 27746
rect 52332 27692 52388 27694
rect 51996 24892 52052 24948
rect 52332 26012 52388 26068
rect 52332 25618 52388 25620
rect 52332 25566 52334 25618
rect 52334 25566 52386 25618
rect 52386 25566 52388 25618
rect 52332 25564 52388 25566
rect 52108 25340 52164 25396
rect 52332 25228 52388 25284
rect 51772 24498 51828 24500
rect 51772 24446 51774 24498
rect 51774 24446 51826 24498
rect 51826 24446 51828 24498
rect 51772 24444 51828 24446
rect 51660 23996 51716 24052
rect 51772 23772 51828 23828
rect 51660 23154 51716 23156
rect 51660 23102 51662 23154
rect 51662 23102 51714 23154
rect 51714 23102 51716 23154
rect 51660 23100 51716 23102
rect 51548 22988 51604 23044
rect 51436 21644 51492 21700
rect 51436 21474 51492 21476
rect 51436 21422 51438 21474
rect 51438 21422 51490 21474
rect 51490 21422 51492 21474
rect 51436 21420 51492 21422
rect 51324 20076 51380 20132
rect 50540 19628 50596 19684
rect 50540 19404 50596 19460
rect 50876 19404 50932 19460
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50764 18450 50820 18452
rect 50764 18398 50766 18450
rect 50766 18398 50818 18450
rect 50818 18398 50820 18450
rect 50764 18396 50820 18398
rect 51884 23660 51940 23716
rect 51884 23378 51940 23380
rect 51884 23326 51886 23378
rect 51886 23326 51938 23378
rect 51938 23326 51940 23378
rect 51884 23324 51940 23326
rect 52108 24668 52164 24724
rect 52556 29372 52612 29428
rect 52892 34636 52948 34692
rect 53900 32508 53956 32564
rect 54908 52162 54964 52164
rect 54908 52110 54910 52162
rect 54910 52110 54962 52162
rect 54962 52110 54964 52162
rect 54908 52108 54964 52110
rect 56028 51772 56084 51828
rect 58156 48860 58212 48916
rect 55356 46396 55412 46452
rect 56140 45724 56196 45780
rect 56700 45836 56756 45892
rect 57372 45890 57428 45892
rect 57372 45838 57374 45890
rect 57374 45838 57426 45890
rect 57426 45838 57428 45890
rect 57372 45836 57428 45838
rect 57148 45778 57204 45780
rect 57148 45726 57150 45778
rect 57150 45726 57202 45778
rect 57202 45726 57204 45778
rect 57148 45724 57204 45726
rect 55356 40348 55412 40404
rect 56140 39452 56196 39508
rect 54348 35922 54404 35924
rect 54348 35870 54350 35922
rect 54350 35870 54402 35922
rect 54402 35870 54404 35922
rect 54348 35868 54404 35870
rect 54908 35868 54964 35924
rect 56028 34972 56084 35028
rect 56588 32732 56644 32788
rect 56700 39564 56756 39620
rect 57372 39618 57428 39620
rect 57372 39566 57374 39618
rect 57374 39566 57426 39618
rect 57426 39566 57428 39618
rect 57372 39564 57428 39566
rect 57148 39506 57204 39508
rect 57148 39454 57150 39506
rect 57150 39454 57202 39506
rect 57202 39454 57204 39506
rect 57148 39452 57204 39454
rect 54236 32060 54292 32116
rect 53900 31948 53956 32004
rect 54684 31948 54740 32004
rect 55020 31948 55076 32004
rect 55356 31948 55412 32004
rect 52780 29372 52836 29428
rect 52892 30828 52948 30884
rect 52668 29260 52724 29316
rect 52668 27074 52724 27076
rect 52668 27022 52670 27074
rect 52670 27022 52722 27074
rect 52722 27022 52724 27074
rect 52668 27020 52724 27022
rect 53340 30828 53396 30884
rect 53788 30882 53844 30884
rect 53788 30830 53790 30882
rect 53790 30830 53842 30882
rect 53842 30830 53844 30882
rect 53788 30828 53844 30830
rect 53116 30268 53172 30324
rect 53788 30268 53844 30324
rect 53452 29596 53508 29652
rect 53564 29426 53620 29428
rect 53564 29374 53566 29426
rect 53566 29374 53618 29426
rect 53618 29374 53620 29426
rect 53564 29372 53620 29374
rect 53004 29314 53060 29316
rect 53004 29262 53006 29314
rect 53006 29262 53058 29314
rect 53058 29262 53060 29314
rect 53004 29260 53060 29262
rect 53452 28530 53508 28532
rect 53452 28478 53454 28530
rect 53454 28478 53506 28530
rect 53506 28478 53508 28530
rect 53452 28476 53508 28478
rect 53004 27580 53060 27636
rect 53676 27916 53732 27972
rect 54236 30268 54292 30324
rect 55244 30828 55300 30884
rect 55692 30882 55748 30884
rect 55692 30830 55694 30882
rect 55694 30830 55746 30882
rect 55746 30830 55748 30882
rect 55692 30828 55748 30830
rect 54460 30268 54516 30324
rect 54572 30380 54628 30436
rect 55356 30268 55412 30324
rect 54908 29986 54964 29988
rect 54908 29934 54910 29986
rect 54910 29934 54962 29986
rect 54962 29934 54964 29986
rect 54908 29932 54964 29934
rect 54572 29820 54628 29876
rect 54348 29538 54404 29540
rect 54348 29486 54350 29538
rect 54350 29486 54402 29538
rect 54402 29486 54404 29538
rect 54348 29484 54404 29486
rect 54908 29426 54964 29428
rect 54908 29374 54910 29426
rect 54910 29374 54962 29426
rect 54962 29374 54964 29426
rect 54908 29372 54964 29374
rect 54012 28364 54068 28420
rect 53900 28082 53956 28084
rect 53900 28030 53902 28082
rect 53902 28030 53954 28082
rect 53954 28030 53956 28082
rect 53900 28028 53956 28030
rect 53228 27020 53284 27076
rect 53900 27580 53956 27636
rect 52556 26348 52612 26404
rect 52668 26290 52724 26292
rect 52668 26238 52670 26290
rect 52670 26238 52722 26290
rect 52722 26238 52724 26290
rect 52668 26236 52724 26238
rect 52892 25788 52948 25844
rect 52668 25676 52724 25732
rect 52668 25228 52724 25284
rect 52556 25116 52612 25172
rect 52220 23324 52276 23380
rect 52108 23212 52164 23268
rect 51884 22988 51940 23044
rect 51884 22764 51940 22820
rect 51996 22652 52052 22708
rect 51772 21980 51828 22036
rect 51660 21644 51716 21700
rect 51884 21586 51940 21588
rect 51884 21534 51886 21586
rect 51886 21534 51938 21586
rect 51938 21534 51940 21586
rect 51884 21532 51940 21534
rect 51884 21084 51940 21140
rect 52108 21980 52164 22036
rect 51772 20412 51828 20468
rect 51548 19964 51604 20020
rect 52108 20524 52164 20580
rect 51324 19906 51380 19908
rect 51324 19854 51326 19906
rect 51326 19854 51378 19906
rect 51378 19854 51380 19906
rect 51324 19852 51380 19854
rect 51772 19628 51828 19684
rect 51324 19404 51380 19460
rect 50988 19234 51044 19236
rect 50988 19182 50990 19234
rect 50990 19182 51042 19234
rect 51042 19182 51044 19234
rect 50988 19180 51044 19182
rect 50988 18732 51044 18788
rect 50988 18508 51044 18564
rect 50988 18060 51044 18116
rect 50876 17724 50932 17780
rect 50316 17442 50372 17444
rect 50316 17390 50318 17442
rect 50318 17390 50370 17442
rect 50370 17390 50372 17442
rect 50316 17388 50372 17390
rect 49532 16156 49588 16212
rect 49308 14418 49364 14420
rect 49308 14366 49310 14418
rect 49310 14366 49362 14418
rect 49362 14366 49364 14418
rect 49308 14364 49364 14366
rect 49420 13746 49476 13748
rect 49420 13694 49422 13746
rect 49422 13694 49474 13746
rect 49474 13694 49476 13746
rect 49420 13692 49476 13694
rect 49980 16716 50036 16772
rect 49868 16098 49924 16100
rect 49868 16046 49870 16098
rect 49870 16046 49922 16098
rect 49922 16046 49924 16098
rect 49868 16044 49924 16046
rect 49756 15986 49812 15988
rect 49756 15934 49758 15986
rect 49758 15934 49810 15986
rect 49810 15934 49812 15986
rect 49756 15932 49812 15934
rect 50092 16268 50148 16324
rect 50204 15932 50260 15988
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50764 16770 50820 16772
rect 50764 16718 50766 16770
rect 50766 16718 50818 16770
rect 50818 16718 50820 16770
rect 50764 16716 50820 16718
rect 50540 16322 50596 16324
rect 50540 16270 50542 16322
rect 50542 16270 50594 16322
rect 50594 16270 50596 16322
rect 50540 16268 50596 16270
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 51996 19404 52052 19460
rect 51324 18450 51380 18452
rect 51324 18398 51326 18450
rect 51326 18398 51378 18450
rect 51378 18398 51380 18450
rect 51324 18396 51380 18398
rect 52780 25004 52836 25060
rect 52780 24220 52836 24276
rect 53564 26572 53620 26628
rect 52556 23660 52612 23716
rect 52668 23938 52724 23940
rect 52668 23886 52670 23938
rect 52670 23886 52722 23938
rect 52722 23886 52724 23938
rect 52668 23884 52724 23886
rect 52668 23548 52724 23604
rect 52556 22594 52612 22596
rect 52556 22542 52558 22594
rect 52558 22542 52610 22594
rect 52610 22542 52612 22594
rect 52556 22540 52612 22542
rect 52556 22316 52612 22372
rect 52668 21868 52724 21924
rect 52668 21420 52724 21476
rect 51548 19122 51604 19124
rect 51548 19070 51550 19122
rect 51550 19070 51602 19122
rect 51602 19070 51604 19122
rect 51548 19068 51604 19070
rect 51996 18844 52052 18900
rect 51660 18620 51716 18676
rect 51884 18396 51940 18452
rect 51324 17948 51380 18004
rect 51212 17666 51268 17668
rect 51212 17614 51214 17666
rect 51214 17614 51266 17666
rect 51266 17614 51268 17666
rect 51212 17612 51268 17614
rect 51100 15986 51156 15988
rect 51100 15934 51102 15986
rect 51102 15934 51154 15986
rect 51154 15934 51156 15986
rect 51100 15932 51156 15934
rect 50316 14924 50372 14980
rect 50204 14642 50260 14644
rect 50204 14590 50206 14642
rect 50206 14590 50258 14642
rect 50258 14590 50260 14642
rect 50204 14588 50260 14590
rect 50540 14530 50596 14532
rect 50540 14478 50542 14530
rect 50542 14478 50594 14530
rect 50594 14478 50596 14530
rect 50540 14476 50596 14478
rect 50316 13916 50372 13972
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 49980 13858 50036 13860
rect 49980 13806 49982 13858
rect 49982 13806 50034 13858
rect 50034 13806 50036 13858
rect 49980 13804 50036 13806
rect 49644 12908 49700 12964
rect 49196 11506 49252 11508
rect 49196 11454 49198 11506
rect 49198 11454 49250 11506
rect 49250 11454 49252 11506
rect 49196 11452 49252 11454
rect 49084 10892 49140 10948
rect 49084 10556 49140 10612
rect 49532 12460 49588 12516
rect 49644 11170 49700 11172
rect 49644 11118 49646 11170
rect 49646 11118 49698 11170
rect 49698 11118 49700 11170
rect 49644 11116 49700 11118
rect 49532 10834 49588 10836
rect 49532 10782 49534 10834
rect 49534 10782 49586 10834
rect 49586 10782 49588 10834
rect 49532 10780 49588 10782
rect 49756 10444 49812 10500
rect 49868 12908 49924 12964
rect 49868 12236 49924 12292
rect 49532 8370 49588 8372
rect 49532 8318 49534 8370
rect 49534 8318 49586 8370
rect 49586 8318 49588 8370
rect 49532 8316 49588 8318
rect 49420 8092 49476 8148
rect 48860 7308 48916 7364
rect 49084 7980 49140 8036
rect 48636 6524 48692 6580
rect 48524 6076 48580 6132
rect 48524 4450 48580 4452
rect 48524 4398 48526 4450
rect 48526 4398 48578 4450
rect 48578 4398 48580 4450
rect 48524 4396 48580 4398
rect 47964 4172 48020 4228
rect 48300 4172 48356 4228
rect 44268 3554 44324 3556
rect 44268 3502 44270 3554
rect 44270 3502 44322 3554
rect 44322 3502 44324 3554
rect 44268 3500 44324 3502
rect 45164 3554 45220 3556
rect 45164 3502 45166 3554
rect 45166 3502 45218 3554
rect 45218 3502 45220 3554
rect 45164 3500 45220 3502
rect 41804 3276 41860 3332
rect 44940 3330 44996 3332
rect 44940 3278 44942 3330
rect 44942 3278 44994 3330
rect 44994 3278 44996 3330
rect 44940 3276 44996 3278
rect 50428 13468 50484 13524
rect 50316 13244 50372 13300
rect 50092 12236 50148 12292
rect 49980 10668 50036 10724
rect 50204 11340 50260 11396
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50764 12348 50820 12404
rect 50764 12012 50820 12068
rect 51548 15874 51604 15876
rect 51548 15822 51550 15874
rect 51550 15822 51602 15874
rect 51602 15822 51604 15874
rect 51548 15820 51604 15822
rect 51212 14476 51268 14532
rect 51324 15708 51380 15764
rect 51100 13916 51156 13972
rect 50988 13468 51044 13524
rect 51100 13132 51156 13188
rect 50988 12290 51044 12292
rect 50988 12238 50990 12290
rect 50990 12238 51042 12290
rect 51042 12238 51044 12290
rect 50988 12236 51044 12238
rect 51436 15148 51492 15204
rect 51436 14588 51492 14644
rect 51436 14140 51492 14196
rect 51548 14476 51604 14532
rect 51100 11788 51156 11844
rect 51100 11506 51156 11508
rect 51100 11454 51102 11506
rect 51102 11454 51154 11506
rect 51154 11454 51156 11506
rect 51100 11452 51156 11454
rect 50316 11282 50372 11284
rect 50316 11230 50318 11282
rect 50318 11230 50370 11282
rect 50370 11230 50372 11282
rect 50316 11228 50372 11230
rect 49980 10444 50036 10500
rect 50652 11394 50708 11396
rect 50652 11342 50654 11394
rect 50654 11342 50706 11394
rect 50706 11342 50708 11394
rect 50652 11340 50708 11342
rect 50764 11116 50820 11172
rect 50876 11228 50932 11284
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50316 9938 50372 9940
rect 50316 9886 50318 9938
rect 50318 9886 50370 9938
rect 50370 9886 50372 9938
rect 50316 9884 50372 9886
rect 50092 9660 50148 9716
rect 50428 9660 50484 9716
rect 50316 9548 50372 9604
rect 49196 6802 49252 6804
rect 49196 6750 49198 6802
rect 49198 6750 49250 6802
rect 49250 6750 49252 6802
rect 49196 6748 49252 6750
rect 49308 6690 49364 6692
rect 49308 6638 49310 6690
rect 49310 6638 49362 6690
rect 49362 6638 49364 6690
rect 49308 6636 49364 6638
rect 49420 5852 49476 5908
rect 49980 7980 50036 8036
rect 50092 7644 50148 7700
rect 49644 7250 49700 7252
rect 49644 7198 49646 7250
rect 49646 7198 49698 7250
rect 49698 7198 49700 7250
rect 49644 7196 49700 7198
rect 49532 6748 49588 6804
rect 50204 7362 50260 7364
rect 50204 7310 50206 7362
rect 50206 7310 50258 7362
rect 50258 7310 50260 7362
rect 50204 7308 50260 7310
rect 50316 7196 50372 7252
rect 49868 6636 49924 6692
rect 49756 6130 49812 6132
rect 49756 6078 49758 6130
rect 49758 6078 49810 6130
rect 49810 6078 49812 6130
rect 49756 6076 49812 6078
rect 49980 6412 50036 6468
rect 49644 4956 49700 5012
rect 49644 3612 49700 3668
rect 50316 5794 50372 5796
rect 50316 5742 50318 5794
rect 50318 5742 50370 5794
rect 50370 5742 50372 5794
rect 50316 5740 50372 5742
rect 50540 9548 50596 9604
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 50764 9100 50820 9156
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50652 7698 50708 7700
rect 50652 7646 50654 7698
rect 50654 7646 50706 7698
rect 50706 7646 50708 7698
rect 50652 7644 50708 7646
rect 50652 6690 50708 6692
rect 50652 6638 50654 6690
rect 50654 6638 50706 6690
rect 50706 6638 50708 6690
rect 50652 6636 50708 6638
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 51436 12572 51492 12628
rect 51884 17388 51940 17444
rect 52108 18060 52164 18116
rect 51772 17276 51828 17332
rect 51996 17164 52052 17220
rect 51772 15314 51828 15316
rect 51772 15262 51774 15314
rect 51774 15262 51826 15314
rect 51826 15262 51828 15314
rect 51772 15260 51828 15262
rect 51772 13468 51828 13524
rect 51996 16268 52052 16324
rect 52444 18060 52500 18116
rect 52332 17052 52388 17108
rect 53004 23884 53060 23940
rect 53004 23660 53060 23716
rect 53228 24610 53284 24612
rect 53228 24558 53230 24610
rect 53230 24558 53282 24610
rect 53282 24558 53284 24610
rect 53228 24556 53284 24558
rect 53788 27020 53844 27076
rect 53452 26348 53508 26404
rect 53452 26124 53508 26180
rect 53676 26012 53732 26068
rect 53900 26460 53956 26516
rect 54012 26348 54068 26404
rect 53452 23938 53508 23940
rect 53452 23886 53454 23938
rect 53454 23886 53506 23938
rect 53506 23886 53508 23938
rect 53452 23884 53508 23886
rect 53564 23548 53620 23604
rect 53116 22764 53172 22820
rect 53004 22316 53060 22372
rect 54684 28588 54740 28644
rect 55020 28588 55076 28644
rect 54572 27916 54628 27972
rect 54236 27746 54292 27748
rect 54236 27694 54238 27746
rect 54238 27694 54290 27746
rect 54290 27694 54292 27746
rect 54236 27692 54292 27694
rect 54236 27468 54292 27524
rect 54348 27074 54404 27076
rect 54348 27022 54350 27074
rect 54350 27022 54402 27074
rect 54402 27022 54404 27074
rect 54348 27020 54404 27022
rect 54684 27356 54740 27412
rect 54908 26402 54964 26404
rect 54908 26350 54910 26402
rect 54910 26350 54962 26402
rect 54962 26350 54964 26402
rect 54908 26348 54964 26350
rect 54236 25394 54292 25396
rect 54236 25342 54238 25394
rect 54238 25342 54290 25394
rect 54290 25342 54292 25394
rect 54236 25340 54292 25342
rect 54124 24780 54180 24836
rect 54012 23826 54068 23828
rect 54012 23774 54014 23826
rect 54014 23774 54066 23826
rect 54066 23774 54068 23826
rect 54012 23772 54068 23774
rect 53900 23714 53956 23716
rect 53900 23662 53902 23714
rect 53902 23662 53954 23714
rect 53954 23662 53956 23714
rect 53900 23660 53956 23662
rect 54012 23548 54068 23604
rect 53788 23266 53844 23268
rect 53788 23214 53790 23266
rect 53790 23214 53842 23266
rect 53842 23214 53844 23266
rect 53788 23212 53844 23214
rect 53228 21644 53284 21700
rect 53228 21474 53284 21476
rect 53228 21422 53230 21474
rect 53230 21422 53282 21474
rect 53282 21422 53284 21474
rect 53228 21420 53284 21422
rect 52780 20188 52836 20244
rect 52892 19964 52948 20020
rect 52892 19516 52948 19572
rect 53452 22764 53508 22820
rect 53900 23324 53956 23380
rect 53900 22652 53956 22708
rect 54012 22540 54068 22596
rect 53676 22204 53732 22260
rect 53452 21980 53508 22036
rect 53788 21980 53844 22036
rect 53004 20524 53060 20580
rect 54236 21868 54292 21924
rect 54236 21644 54292 21700
rect 54124 21586 54180 21588
rect 54124 21534 54126 21586
rect 54126 21534 54178 21586
rect 54178 21534 54180 21586
rect 54124 21532 54180 21534
rect 54012 20860 54068 20916
rect 53452 20524 53508 20580
rect 52668 18508 52724 18564
rect 52780 18450 52836 18452
rect 52780 18398 52782 18450
rect 52782 18398 52834 18450
rect 52834 18398 52836 18450
rect 52780 18396 52836 18398
rect 52780 18060 52836 18116
rect 52556 17948 52612 18004
rect 53340 20242 53396 20244
rect 53340 20190 53342 20242
rect 53342 20190 53394 20242
rect 53394 20190 53396 20242
rect 53340 20188 53396 20190
rect 52220 16492 52276 16548
rect 52220 16268 52276 16324
rect 52668 17052 52724 17108
rect 52108 15092 52164 15148
rect 53004 17106 53060 17108
rect 53004 17054 53006 17106
rect 53006 17054 53058 17106
rect 53058 17054 53060 17106
rect 53004 17052 53060 17054
rect 53788 20018 53844 20020
rect 53788 19966 53790 20018
rect 53790 19966 53842 20018
rect 53842 19966 53844 20018
rect 53788 19964 53844 19966
rect 53340 19516 53396 19572
rect 54124 20802 54180 20804
rect 54124 20750 54126 20802
rect 54126 20750 54178 20802
rect 54178 20750 54180 20802
rect 54124 20748 54180 20750
rect 54124 20412 54180 20468
rect 54012 19010 54068 19012
rect 54012 18958 54014 19010
rect 54014 18958 54066 19010
rect 54066 18958 54068 19010
rect 54012 18956 54068 18958
rect 53900 18844 53956 18900
rect 53676 18450 53732 18452
rect 53676 18398 53678 18450
rect 53678 18398 53730 18450
rect 53730 18398 53732 18450
rect 53676 18396 53732 18398
rect 53900 18450 53956 18452
rect 53900 18398 53902 18450
rect 53902 18398 53954 18450
rect 53954 18398 53956 18450
rect 53900 18396 53956 18398
rect 53340 18284 53396 18340
rect 53452 17666 53508 17668
rect 53452 17614 53454 17666
rect 53454 17614 53506 17666
rect 53506 17614 53508 17666
rect 53452 17612 53508 17614
rect 53340 17388 53396 17444
rect 53228 17276 53284 17332
rect 53788 17052 53844 17108
rect 53452 16994 53508 16996
rect 53452 16942 53454 16994
rect 53454 16942 53506 16994
rect 53506 16942 53508 16994
rect 53452 16940 53508 16942
rect 53228 16268 53284 16324
rect 53340 15874 53396 15876
rect 53340 15822 53342 15874
rect 53342 15822 53394 15874
rect 53394 15822 53396 15874
rect 53340 15820 53396 15822
rect 52668 15426 52724 15428
rect 52668 15374 52670 15426
rect 52670 15374 52722 15426
rect 52722 15374 52724 15426
rect 52668 15372 52724 15374
rect 52556 15314 52612 15316
rect 52556 15262 52558 15314
rect 52558 15262 52610 15314
rect 52610 15262 52612 15314
rect 52556 15260 52612 15262
rect 52780 15148 52836 15204
rect 52108 14924 52164 14980
rect 52332 14924 52388 14980
rect 52220 13746 52276 13748
rect 52220 13694 52222 13746
rect 52222 13694 52274 13746
rect 52274 13694 52276 13746
rect 52220 13692 52276 13694
rect 52332 14700 52388 14756
rect 52220 13356 52276 13412
rect 51660 12572 51716 12628
rect 51772 13020 51828 13076
rect 51996 12796 52052 12852
rect 51884 12684 51940 12740
rect 51324 12124 51380 12180
rect 51660 12236 51716 12292
rect 51772 12124 51828 12180
rect 51212 11228 51268 11284
rect 51436 12012 51492 12068
rect 51100 10722 51156 10724
rect 51100 10670 51102 10722
rect 51102 10670 51154 10722
rect 51154 10670 51156 10722
rect 51100 10668 51156 10670
rect 51100 10108 51156 10164
rect 50988 8146 51044 8148
rect 50988 8094 50990 8146
rect 50990 8094 51042 8146
rect 51042 8094 51044 8146
rect 50988 8092 51044 8094
rect 51212 9884 51268 9940
rect 51660 11788 51716 11844
rect 51660 11564 51716 11620
rect 51548 11340 51604 11396
rect 51884 11564 51940 11620
rect 51996 12236 52052 12292
rect 51660 10108 51716 10164
rect 51324 9714 51380 9716
rect 51324 9662 51326 9714
rect 51326 9662 51378 9714
rect 51378 9662 51380 9714
rect 51324 9660 51380 9662
rect 51324 9100 51380 9156
rect 51884 9548 51940 9604
rect 51884 8988 51940 9044
rect 52220 11564 52276 11620
rect 52108 9884 52164 9940
rect 52108 9714 52164 9716
rect 52108 9662 52110 9714
rect 52110 9662 52162 9714
rect 52162 9662 52164 9714
rect 52108 9660 52164 9662
rect 51212 7980 51268 8036
rect 51100 6972 51156 7028
rect 50988 6524 51044 6580
rect 51660 8146 51716 8148
rect 51660 8094 51662 8146
rect 51662 8094 51714 8146
rect 51714 8094 51716 8146
rect 51660 8092 51716 8094
rect 51772 8034 51828 8036
rect 51772 7982 51774 8034
rect 51774 7982 51826 8034
rect 51826 7982 51828 8034
rect 51772 7980 51828 7982
rect 51324 6914 51380 6916
rect 51324 6862 51326 6914
rect 51326 6862 51378 6914
rect 51378 6862 51380 6914
rect 51324 6860 51380 6862
rect 51996 8316 52052 8372
rect 51996 7196 52052 7252
rect 52108 6524 52164 6580
rect 51996 6466 52052 6468
rect 51996 6414 51998 6466
rect 51998 6414 52050 6466
rect 52050 6414 52052 6466
rect 51996 6412 52052 6414
rect 52556 14306 52612 14308
rect 52556 14254 52558 14306
rect 52558 14254 52610 14306
rect 52610 14254 52612 14306
rect 52556 14252 52612 14254
rect 52444 14140 52500 14196
rect 52444 13970 52500 13972
rect 52444 13918 52446 13970
rect 52446 13918 52498 13970
rect 52498 13918 52500 13970
rect 52444 13916 52500 13918
rect 52556 13468 52612 13524
rect 52668 13074 52724 13076
rect 52668 13022 52670 13074
rect 52670 13022 52722 13074
rect 52722 13022 52724 13074
rect 52668 13020 52724 13022
rect 52556 12684 52612 12740
rect 52332 9884 52388 9940
rect 52444 11676 52500 11732
rect 52668 12066 52724 12068
rect 52668 12014 52670 12066
rect 52670 12014 52722 12066
rect 52722 12014 52724 12066
rect 52668 12012 52724 12014
rect 52556 11170 52612 11172
rect 52556 11118 52558 11170
rect 52558 11118 52610 11170
rect 52610 11118 52612 11170
rect 52556 11116 52612 11118
rect 52556 9938 52612 9940
rect 52556 9886 52558 9938
rect 52558 9886 52610 9938
rect 52610 9886 52612 9938
rect 52556 9884 52612 9886
rect 53228 15314 53284 15316
rect 53228 15262 53230 15314
rect 53230 15262 53282 15314
rect 53282 15262 53284 15314
rect 53228 15260 53284 15262
rect 53340 15148 53396 15204
rect 52892 14364 52948 14420
rect 53004 12684 53060 12740
rect 53116 14924 53172 14980
rect 54124 17948 54180 18004
rect 54460 25116 54516 25172
rect 54796 24834 54852 24836
rect 54796 24782 54798 24834
rect 54798 24782 54850 24834
rect 54850 24782 54852 24834
rect 54796 24780 54852 24782
rect 54908 24556 54964 24612
rect 55468 29986 55524 29988
rect 55468 29934 55470 29986
rect 55470 29934 55522 29986
rect 55522 29934 55524 29986
rect 55468 29932 55524 29934
rect 55580 29484 55636 29540
rect 55468 27970 55524 27972
rect 55468 27918 55470 27970
rect 55470 27918 55522 27970
rect 55522 27918 55524 27970
rect 55468 27916 55524 27918
rect 55244 25564 55300 25620
rect 55356 26572 55412 26628
rect 55132 25506 55188 25508
rect 55132 25454 55134 25506
rect 55134 25454 55186 25506
rect 55186 25454 55188 25506
rect 55132 25452 55188 25454
rect 55356 25116 55412 25172
rect 55132 24108 55188 24164
rect 55020 23378 55076 23380
rect 55020 23326 55022 23378
rect 55022 23326 55074 23378
rect 55074 23326 55076 23378
rect 55020 23324 55076 23326
rect 55244 23324 55300 23380
rect 55468 24444 55524 24500
rect 55804 27580 55860 27636
rect 55692 25452 55748 25508
rect 56700 31836 56756 31892
rect 56364 31500 56420 31556
rect 56700 30604 56756 30660
rect 56028 28924 56084 28980
rect 56140 28700 56196 28756
rect 56364 29820 56420 29876
rect 56364 29260 56420 29316
rect 56588 29484 56644 29540
rect 57372 32450 57428 32452
rect 57372 32398 57374 32450
rect 57374 32398 57426 32450
rect 57426 32398 57428 32450
rect 57372 32396 57428 32398
rect 57148 31500 57204 31556
rect 57036 30604 57092 30660
rect 56924 29820 56980 29876
rect 56700 28588 56756 28644
rect 56476 28476 56532 28532
rect 56588 28364 56644 28420
rect 56364 27804 56420 27860
rect 56252 27298 56308 27300
rect 56252 27246 56254 27298
rect 56254 27246 56306 27298
rect 56306 27246 56308 27298
rect 56252 27244 56308 27246
rect 56028 25676 56084 25732
rect 56252 26290 56308 26292
rect 56252 26238 56254 26290
rect 56254 26238 56306 26290
rect 56306 26238 56308 26290
rect 56252 26236 56308 26238
rect 55916 25116 55972 25172
rect 56028 25004 56084 25060
rect 56140 25228 56196 25284
rect 55580 23324 55636 23380
rect 55132 23042 55188 23044
rect 55132 22990 55134 23042
rect 55134 22990 55186 23042
rect 55186 22990 55188 23042
rect 55132 22988 55188 22990
rect 55244 22540 55300 22596
rect 56812 26796 56868 26852
rect 56812 26236 56868 26292
rect 56476 25506 56532 25508
rect 56476 25454 56478 25506
rect 56478 25454 56530 25506
rect 56530 25454 56532 25506
rect 56476 25452 56532 25454
rect 56140 24610 56196 24612
rect 56140 24558 56142 24610
rect 56142 24558 56194 24610
rect 56194 24558 56196 24610
rect 56140 24556 56196 24558
rect 55804 24498 55860 24500
rect 55804 24446 55806 24498
rect 55806 24446 55858 24498
rect 55858 24446 55860 24498
rect 55804 24444 55860 24446
rect 55692 22764 55748 22820
rect 54348 20860 54404 20916
rect 54684 22428 54740 22484
rect 54796 22258 54852 22260
rect 54796 22206 54798 22258
rect 54798 22206 54850 22258
rect 54850 22206 54852 22258
rect 54796 22204 54852 22206
rect 55132 22146 55188 22148
rect 55132 22094 55134 22146
rect 55134 22094 55186 22146
rect 55186 22094 55188 22146
rect 55132 22092 55188 22094
rect 55580 22146 55636 22148
rect 55580 22094 55582 22146
rect 55582 22094 55634 22146
rect 55634 22094 55636 22146
rect 55580 22092 55636 22094
rect 55132 21868 55188 21924
rect 54348 20188 54404 20244
rect 54572 20636 54628 20692
rect 54460 19964 54516 20020
rect 54348 19122 54404 19124
rect 54348 19070 54350 19122
rect 54350 19070 54402 19122
rect 54402 19070 54404 19122
rect 54348 19068 54404 19070
rect 54348 18732 54404 18788
rect 54460 18620 54516 18676
rect 54460 18450 54516 18452
rect 54460 18398 54462 18450
rect 54462 18398 54514 18450
rect 54514 18398 54516 18450
rect 54460 18396 54516 18398
rect 54236 17612 54292 17668
rect 54236 17442 54292 17444
rect 54236 17390 54238 17442
rect 54238 17390 54290 17442
rect 54290 17390 54292 17442
rect 54236 17388 54292 17390
rect 54684 20412 54740 20468
rect 55020 21698 55076 21700
rect 55020 21646 55022 21698
rect 55022 21646 55074 21698
rect 55074 21646 55076 21698
rect 55020 21644 55076 21646
rect 54796 20018 54852 20020
rect 54796 19966 54798 20018
rect 54798 19966 54850 20018
rect 54850 19966 54852 20018
rect 54796 19964 54852 19966
rect 55916 24332 55972 24388
rect 55244 21644 55300 21700
rect 55804 22316 55860 22372
rect 54908 19068 54964 19124
rect 55020 20972 55076 21028
rect 55132 19964 55188 20020
rect 55692 21474 55748 21476
rect 55692 21422 55694 21474
rect 55694 21422 55746 21474
rect 55746 21422 55748 21474
rect 55692 21420 55748 21422
rect 55580 20578 55636 20580
rect 55580 20526 55582 20578
rect 55582 20526 55634 20578
rect 55634 20526 55636 20578
rect 55580 20524 55636 20526
rect 55580 19404 55636 19460
rect 54684 18284 54740 18340
rect 54796 18844 54852 18900
rect 54124 16044 54180 16100
rect 53676 15484 53732 15540
rect 54012 15932 54068 15988
rect 53676 15148 53732 15204
rect 53788 14812 53844 14868
rect 53228 14252 53284 14308
rect 53228 12684 53284 12740
rect 53452 13858 53508 13860
rect 53452 13806 53454 13858
rect 53454 13806 53506 13858
rect 53506 13806 53508 13858
rect 53452 13804 53508 13806
rect 53564 14252 53620 14308
rect 53564 14028 53620 14084
rect 53788 13580 53844 13636
rect 54124 15036 54180 15092
rect 54236 15260 54292 15316
rect 54124 14418 54180 14420
rect 54124 14366 54126 14418
rect 54126 14366 54178 14418
rect 54178 14366 54180 14418
rect 54124 14364 54180 14366
rect 54460 16268 54516 16324
rect 54460 15372 54516 15428
rect 54348 14252 54404 14308
rect 54236 13580 54292 13636
rect 54012 13356 54068 13412
rect 54124 13468 54180 13524
rect 53900 13244 53956 13300
rect 53452 12850 53508 12852
rect 53452 12798 53454 12850
rect 53454 12798 53506 12850
rect 53506 12798 53508 12850
rect 53452 12796 53508 12798
rect 53676 12738 53732 12740
rect 53676 12686 53678 12738
rect 53678 12686 53730 12738
rect 53730 12686 53732 12738
rect 53676 12684 53732 12686
rect 53452 12236 53508 12292
rect 52780 10892 52836 10948
rect 52892 11228 52948 11284
rect 52780 10722 52836 10724
rect 52780 10670 52782 10722
rect 52782 10670 52834 10722
rect 52834 10670 52836 10722
rect 52780 10668 52836 10670
rect 52668 9100 52724 9156
rect 53676 12236 53732 12292
rect 53004 9548 53060 9604
rect 53116 11900 53172 11956
rect 52444 8258 52500 8260
rect 52444 8206 52446 8258
rect 52446 8206 52498 8258
rect 52498 8206 52500 8258
rect 52444 8204 52500 8206
rect 53004 8204 53060 8260
rect 52780 8034 52836 8036
rect 52780 7982 52782 8034
rect 52782 7982 52834 8034
rect 52834 7982 52836 8034
rect 52780 7980 52836 7982
rect 52556 6690 52612 6692
rect 52556 6638 52558 6690
rect 52558 6638 52610 6690
rect 52610 6638 52612 6690
rect 52556 6636 52612 6638
rect 50204 4956 50260 5012
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 53004 7196 53060 7252
rect 53004 6018 53060 6020
rect 53004 5966 53006 6018
rect 53006 5966 53058 6018
rect 53058 5966 53060 6018
rect 53004 5964 53060 5966
rect 52780 4508 52836 4564
rect 50652 4396 50708 4452
rect 50428 3612 50484 3668
rect 49868 2940 49924 2996
rect 49084 2828 49140 2884
rect 51324 3666 51380 3668
rect 51324 3614 51326 3666
rect 51326 3614 51378 3666
rect 51378 3614 51380 3666
rect 51324 3612 51380 3614
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 53564 12178 53620 12180
rect 53564 12126 53566 12178
rect 53566 12126 53618 12178
rect 53618 12126 53620 12178
rect 53564 12124 53620 12126
rect 53228 11228 53284 11284
rect 53452 12012 53508 12068
rect 53340 10722 53396 10724
rect 53340 10670 53342 10722
rect 53342 10670 53394 10722
rect 53394 10670 53396 10722
rect 53340 10668 53396 10670
rect 53340 9826 53396 9828
rect 53340 9774 53342 9826
rect 53342 9774 53394 9826
rect 53394 9774 53396 9826
rect 53340 9772 53396 9774
rect 53788 11564 53844 11620
rect 53788 11394 53844 11396
rect 53788 11342 53790 11394
rect 53790 11342 53842 11394
rect 53842 11342 53844 11394
rect 53788 11340 53844 11342
rect 54236 12796 54292 12852
rect 54236 12460 54292 12516
rect 54236 12290 54292 12292
rect 54236 12238 54238 12290
rect 54238 12238 54290 12290
rect 54290 12238 54292 12290
rect 54236 12236 54292 12238
rect 53564 11116 53620 11172
rect 53900 11170 53956 11172
rect 53900 11118 53902 11170
rect 53902 11118 53954 11170
rect 53954 11118 53956 11170
rect 53900 11116 53956 11118
rect 54124 11676 54180 11732
rect 54460 14028 54516 14084
rect 54460 13580 54516 13636
rect 54460 11564 54516 11620
rect 54908 17666 54964 17668
rect 54908 17614 54910 17666
rect 54910 17614 54962 17666
rect 54962 17614 54964 17666
rect 54908 17612 54964 17614
rect 54796 16716 54852 16772
rect 54908 17276 54964 17332
rect 54796 15036 54852 15092
rect 54684 14476 54740 14532
rect 54796 14252 54852 14308
rect 54684 12796 54740 12852
rect 54796 13356 54852 13412
rect 54684 12402 54740 12404
rect 54684 12350 54686 12402
rect 54686 12350 54738 12402
rect 54738 12350 54740 12402
rect 54684 12348 54740 12350
rect 53788 9938 53844 9940
rect 53788 9886 53790 9938
rect 53790 9886 53842 9938
rect 53842 9886 53844 9938
rect 53788 9884 53844 9886
rect 53340 8204 53396 8260
rect 53452 9100 53508 9156
rect 53228 7980 53284 8036
rect 53340 7308 53396 7364
rect 53564 8930 53620 8932
rect 53564 8878 53566 8930
rect 53566 8878 53618 8930
rect 53618 8878 53620 8930
rect 53564 8876 53620 8878
rect 53788 8370 53844 8372
rect 53788 8318 53790 8370
rect 53790 8318 53842 8370
rect 53842 8318 53844 8370
rect 53788 8316 53844 8318
rect 53788 7868 53844 7924
rect 53788 7084 53844 7140
rect 53564 6860 53620 6916
rect 53452 6690 53508 6692
rect 53452 6638 53454 6690
rect 53454 6638 53506 6690
rect 53506 6638 53508 6690
rect 53452 6636 53508 6638
rect 53788 6130 53844 6132
rect 53788 6078 53790 6130
rect 53790 6078 53842 6130
rect 53842 6078 53844 6130
rect 53788 6076 53844 6078
rect 54012 10220 54068 10276
rect 54348 9714 54404 9716
rect 54348 9662 54350 9714
rect 54350 9662 54402 9714
rect 54402 9662 54404 9714
rect 54348 9660 54404 9662
rect 54684 11004 54740 11060
rect 54572 10834 54628 10836
rect 54572 10782 54574 10834
rect 54574 10782 54626 10834
rect 54626 10782 54628 10834
rect 54572 10780 54628 10782
rect 54572 10444 54628 10500
rect 55132 19068 55188 19124
rect 55356 19292 55412 19348
rect 55468 19234 55524 19236
rect 55468 19182 55470 19234
rect 55470 19182 55522 19234
rect 55522 19182 55524 19234
rect 55468 19180 55524 19182
rect 55244 18844 55300 18900
rect 55132 16882 55188 16884
rect 55132 16830 55134 16882
rect 55134 16830 55186 16882
rect 55186 16830 55188 16882
rect 55132 16828 55188 16830
rect 55020 15820 55076 15876
rect 55020 15596 55076 15652
rect 55692 18620 55748 18676
rect 55468 17052 55524 17108
rect 55356 16716 55412 16772
rect 55020 14530 55076 14532
rect 55020 14478 55022 14530
rect 55022 14478 55074 14530
rect 55074 14478 55076 14530
rect 55020 14476 55076 14478
rect 55580 16380 55636 16436
rect 55692 16604 55748 16660
rect 55692 15986 55748 15988
rect 55692 15934 55694 15986
rect 55694 15934 55746 15986
rect 55746 15934 55748 15986
rect 55692 15932 55748 15934
rect 56028 23548 56084 23604
rect 56140 23378 56196 23380
rect 56140 23326 56142 23378
rect 56142 23326 56194 23378
rect 56194 23326 56196 23378
rect 56140 23324 56196 23326
rect 56028 20972 56084 21028
rect 56476 23324 56532 23380
rect 56700 22316 56756 22372
rect 57708 31554 57764 31556
rect 57708 31502 57710 31554
rect 57710 31502 57762 31554
rect 57762 31502 57764 31554
rect 57708 31500 57764 31502
rect 57820 30882 57876 30884
rect 57820 30830 57822 30882
rect 57822 30830 57874 30882
rect 57874 30830 57876 30882
rect 57820 30828 57876 30830
rect 57372 29484 57428 29540
rect 57596 28642 57652 28644
rect 57596 28590 57598 28642
rect 57598 28590 57650 28642
rect 57650 28590 57652 28642
rect 57596 28588 57652 28590
rect 57260 28530 57316 28532
rect 57260 28478 57262 28530
rect 57262 28478 57314 28530
rect 57314 28478 57316 28530
rect 57260 28476 57316 28478
rect 57372 27970 57428 27972
rect 57372 27918 57374 27970
rect 57374 27918 57426 27970
rect 57426 27918 57428 27970
rect 57372 27916 57428 27918
rect 57372 26850 57428 26852
rect 57372 26798 57374 26850
rect 57374 26798 57426 26850
rect 57426 26798 57428 26850
rect 57372 26796 57428 26798
rect 57372 26402 57428 26404
rect 57372 26350 57374 26402
rect 57374 26350 57426 26402
rect 57426 26350 57428 26402
rect 57372 26348 57428 26350
rect 58044 28642 58100 28644
rect 58044 28590 58046 28642
rect 58046 28590 58098 28642
rect 58098 28590 58100 28642
rect 58044 28588 58100 28590
rect 57820 28364 57876 28420
rect 57820 27746 57876 27748
rect 57820 27694 57822 27746
rect 57822 27694 57874 27746
rect 57874 27694 57876 27746
rect 57820 27692 57876 27694
rect 57708 26572 57764 26628
rect 57036 24444 57092 24500
rect 56924 24108 56980 24164
rect 57820 25116 57876 25172
rect 56924 23324 56980 23380
rect 56812 22204 56868 22260
rect 56476 21644 56532 21700
rect 56364 21308 56420 21364
rect 56588 20300 56644 20356
rect 56140 19180 56196 19236
rect 56252 18562 56308 18564
rect 56252 18510 56254 18562
rect 56254 18510 56306 18562
rect 56306 18510 56308 18562
rect 56252 18508 56308 18510
rect 55916 18172 55972 18228
rect 56028 17724 56084 17780
rect 57372 24444 57428 24500
rect 57596 24162 57652 24164
rect 57596 24110 57598 24162
rect 57598 24110 57650 24162
rect 57650 24110 57652 24162
rect 57596 24108 57652 24110
rect 57820 23996 57876 24052
rect 58044 25116 58100 25172
rect 57484 23378 57540 23380
rect 57484 23326 57486 23378
rect 57486 23326 57538 23378
rect 57538 23326 57540 23378
rect 57484 23324 57540 23326
rect 58380 32396 58436 32452
rect 58268 30828 58324 30884
rect 58156 22876 58212 22932
rect 57708 21868 57764 21924
rect 57260 21084 57316 21140
rect 57260 19292 57316 19348
rect 56476 18450 56532 18452
rect 56476 18398 56478 18450
rect 56478 18398 56530 18450
rect 56530 18398 56532 18450
rect 56476 18396 56532 18398
rect 56588 18284 56644 18340
rect 56364 16828 56420 16884
rect 56476 17388 56532 17444
rect 56700 17554 56756 17556
rect 56700 17502 56702 17554
rect 56702 17502 56754 17554
rect 56754 17502 56756 17554
rect 56700 17500 56756 17502
rect 56028 16492 56084 16548
rect 55804 15314 55860 15316
rect 55804 15262 55806 15314
rect 55806 15262 55858 15314
rect 55858 15262 55860 15314
rect 55804 15260 55860 15262
rect 55132 14418 55188 14420
rect 55132 14366 55134 14418
rect 55134 14366 55186 14418
rect 55186 14366 55188 14418
rect 55132 14364 55188 14366
rect 55692 15202 55748 15204
rect 55692 15150 55694 15202
rect 55694 15150 55746 15202
rect 55746 15150 55748 15202
rect 55692 15148 55748 15150
rect 55132 14028 55188 14084
rect 55020 13468 55076 13524
rect 54908 13074 54964 13076
rect 54908 13022 54910 13074
rect 54910 13022 54962 13074
rect 54962 13022 54964 13074
rect 54908 13020 54964 13022
rect 54796 9772 54852 9828
rect 54460 9212 54516 9268
rect 54348 8428 54404 8484
rect 54572 8258 54628 8260
rect 54572 8206 54574 8258
rect 54574 8206 54626 8258
rect 54626 8206 54628 8258
rect 54572 8204 54628 8206
rect 54460 7868 54516 7924
rect 54348 7084 54404 7140
rect 54236 6690 54292 6692
rect 54236 6638 54238 6690
rect 54238 6638 54290 6690
rect 54290 6638 54292 6690
rect 54236 6636 54292 6638
rect 54012 6076 54068 6132
rect 54124 6524 54180 6580
rect 54012 5852 54068 5908
rect 53116 2492 53172 2548
rect 54908 12796 54964 12852
rect 54908 11900 54964 11956
rect 55020 11564 55076 11620
rect 55132 11506 55188 11508
rect 55132 11454 55134 11506
rect 55134 11454 55186 11506
rect 55186 11454 55188 11506
rect 55132 11452 55188 11454
rect 55356 14306 55412 14308
rect 55356 14254 55358 14306
rect 55358 14254 55410 14306
rect 55410 14254 55412 14306
rect 55356 14252 55412 14254
rect 55580 14140 55636 14196
rect 55468 14028 55524 14084
rect 56028 15820 56084 15876
rect 56700 16828 56756 16884
rect 56364 15932 56420 15988
rect 56700 16604 56756 16660
rect 56252 15820 56308 15876
rect 56812 15932 56868 15988
rect 56364 15314 56420 15316
rect 56364 15262 56366 15314
rect 56366 15262 56418 15314
rect 56418 15262 56420 15314
rect 56364 15260 56420 15262
rect 56140 14418 56196 14420
rect 56140 14366 56142 14418
rect 56142 14366 56194 14418
rect 56194 14366 56196 14418
rect 56140 14364 56196 14366
rect 55356 13858 55412 13860
rect 55356 13806 55358 13858
rect 55358 13806 55410 13858
rect 55410 13806 55412 13858
rect 55356 13804 55412 13806
rect 55580 13468 55636 13524
rect 55356 12236 55412 12292
rect 55020 10444 55076 10500
rect 55244 9938 55300 9940
rect 55244 9886 55246 9938
rect 55246 9886 55298 9938
rect 55298 9886 55300 9938
rect 55244 9884 55300 9886
rect 55020 8876 55076 8932
rect 55244 8204 55300 8260
rect 54908 7196 54964 7252
rect 54348 5234 54404 5236
rect 54348 5182 54350 5234
rect 54350 5182 54402 5234
rect 54402 5182 54404 5234
rect 54348 5180 54404 5182
rect 54908 6018 54964 6020
rect 54908 5966 54910 6018
rect 54910 5966 54962 6018
rect 54962 5966 54964 6018
rect 54908 5964 54964 5966
rect 55244 7868 55300 7924
rect 55804 13020 55860 13076
rect 55692 12066 55748 12068
rect 55692 12014 55694 12066
rect 55694 12014 55746 12066
rect 55746 12014 55748 12066
rect 55692 12012 55748 12014
rect 56028 12402 56084 12404
rect 56028 12350 56030 12402
rect 56030 12350 56082 12402
rect 56082 12350 56084 12402
rect 56028 12348 56084 12350
rect 56140 12124 56196 12180
rect 56028 10498 56084 10500
rect 56028 10446 56030 10498
rect 56030 10446 56082 10498
rect 56082 10446 56084 10498
rect 56028 10444 56084 10446
rect 55580 9996 55636 10052
rect 56028 9602 56084 9604
rect 56028 9550 56030 9602
rect 56030 9550 56082 9602
rect 56082 9550 56084 9602
rect 56028 9548 56084 9550
rect 56028 9324 56084 9380
rect 55468 8428 55524 8484
rect 55916 8204 55972 8260
rect 55468 8034 55524 8036
rect 55468 7982 55470 8034
rect 55470 7982 55522 8034
rect 55522 7982 55524 8034
rect 55468 7980 55524 7982
rect 55804 8034 55860 8036
rect 55804 7982 55806 8034
rect 55806 7982 55858 8034
rect 55858 7982 55860 8034
rect 55804 7980 55860 7982
rect 55356 6748 55412 6804
rect 55356 6578 55412 6580
rect 55356 6526 55358 6578
rect 55358 6526 55410 6578
rect 55410 6526 55412 6578
rect 55356 6524 55412 6526
rect 55804 7420 55860 7476
rect 56028 8092 56084 8148
rect 57148 18284 57204 18340
rect 57484 21196 57540 21252
rect 57820 22316 57876 22372
rect 59388 24556 59444 24612
rect 58604 22876 58660 22932
rect 57484 20242 57540 20244
rect 57484 20190 57486 20242
rect 57486 20190 57538 20242
rect 57538 20190 57540 20242
rect 57484 20188 57540 20190
rect 57484 18562 57540 18564
rect 57484 18510 57486 18562
rect 57486 18510 57538 18562
rect 57538 18510 57540 18562
rect 57484 18508 57540 18510
rect 57708 18284 57764 18340
rect 57036 17500 57092 17556
rect 56700 15426 56756 15428
rect 56700 15374 56702 15426
rect 56702 15374 56754 15426
rect 56754 15374 56756 15426
rect 56700 15372 56756 15374
rect 56364 13804 56420 13860
rect 56700 14140 56756 14196
rect 56476 13692 56532 13748
rect 56588 13634 56644 13636
rect 56588 13582 56590 13634
rect 56590 13582 56642 13634
rect 56642 13582 56644 13634
rect 56588 13580 56644 13582
rect 57932 19740 57988 19796
rect 58044 18284 58100 18340
rect 58044 18060 58100 18116
rect 58268 18732 58324 18788
rect 57148 16492 57204 16548
rect 57372 15986 57428 15988
rect 57372 15934 57374 15986
rect 57374 15934 57426 15986
rect 57426 15934 57428 15986
rect 57372 15932 57428 15934
rect 56812 12908 56868 12964
rect 57260 15596 57316 15652
rect 56812 12572 56868 12628
rect 57036 14306 57092 14308
rect 57036 14254 57038 14306
rect 57038 14254 57090 14306
rect 57090 14254 57092 14306
rect 57036 14252 57092 14254
rect 57484 15314 57540 15316
rect 57484 15262 57486 15314
rect 57486 15262 57538 15314
rect 57538 15262 57540 15314
rect 57484 15260 57540 15262
rect 57484 14140 57540 14196
rect 57372 13692 57428 13748
rect 57260 13074 57316 13076
rect 57260 13022 57262 13074
rect 57262 13022 57314 13074
rect 57314 13022 57316 13074
rect 57260 13020 57316 13022
rect 57036 12908 57092 12964
rect 57036 12012 57092 12068
rect 57148 12460 57204 12516
rect 56476 11452 56532 11508
rect 56476 10892 56532 10948
rect 57036 10780 57092 10836
rect 57372 11506 57428 11508
rect 57372 11454 57374 11506
rect 57374 11454 57426 11506
rect 57426 11454 57428 11506
rect 57372 11452 57428 11454
rect 56364 10556 56420 10612
rect 57372 9996 57428 10052
rect 57372 9660 57428 9716
rect 56476 9602 56532 9604
rect 56476 9550 56478 9602
rect 56478 9550 56530 9602
rect 56530 9550 56532 9602
rect 56476 9548 56532 9550
rect 56476 9266 56532 9268
rect 56476 9214 56478 9266
rect 56478 9214 56530 9266
rect 56530 9214 56532 9266
rect 56476 9212 56532 9214
rect 55468 5852 55524 5908
rect 57484 8370 57540 8372
rect 57484 8318 57486 8370
rect 57486 8318 57538 8370
rect 57538 8318 57540 8370
rect 57484 8316 57540 8318
rect 56812 7698 56868 7700
rect 56812 7646 56814 7698
rect 56814 7646 56866 7698
rect 56866 7646 56868 7698
rect 56812 7644 56868 7646
rect 56812 6690 56868 6692
rect 56812 6638 56814 6690
rect 56814 6638 56866 6690
rect 56866 6638 56868 6690
rect 56812 6636 56868 6638
rect 55580 5234 55636 5236
rect 55580 5182 55582 5234
rect 55582 5182 55634 5234
rect 55634 5182 55636 5234
rect 55580 5180 55636 5182
rect 57708 16828 57764 16884
rect 58044 14642 58100 14644
rect 58044 14590 58046 14642
rect 58046 14590 58098 14642
rect 58098 14590 58100 14642
rect 58044 14588 58100 14590
rect 57932 14028 57988 14084
rect 57708 13804 57764 13860
rect 58044 13804 58100 13860
rect 57708 12738 57764 12740
rect 57708 12686 57710 12738
rect 57710 12686 57762 12738
rect 57762 12686 57764 12738
rect 57708 12684 57764 12686
rect 57932 12572 57988 12628
rect 57820 12066 57876 12068
rect 57820 12014 57822 12066
rect 57822 12014 57874 12066
rect 57874 12014 57876 12066
rect 57820 12012 57876 12014
rect 57708 11788 57764 11844
rect 58044 12236 58100 12292
rect 58156 12348 58212 12404
rect 57932 11564 57988 11620
rect 57820 10834 57876 10836
rect 57820 10782 57822 10834
rect 57822 10782 57874 10834
rect 57874 10782 57876 10834
rect 57820 10780 57876 10782
rect 57708 9884 57764 9940
rect 58044 9826 58100 9828
rect 58044 9774 58046 9826
rect 58046 9774 58098 9826
rect 58098 9774 58100 9826
rect 58044 9772 58100 9774
rect 57932 8092 57988 8148
rect 58380 11452 58436 11508
rect 58492 18284 58548 18340
rect 58492 9996 58548 10052
rect 58268 9324 58324 9380
rect 57148 6972 57204 7028
rect 58044 7698 58100 7700
rect 58044 7646 58046 7698
rect 58046 7646 58098 7698
rect 58098 7646 58100 7698
rect 58044 7644 58100 7646
rect 57372 5906 57428 5908
rect 57372 5854 57374 5906
rect 57374 5854 57426 5906
rect 57426 5854 57428 5906
rect 57372 5852 57428 5854
rect 56924 4956 56980 5012
rect 54236 4844 54292 4900
rect 55916 4396 55972 4452
rect 54348 4284 54404 4340
rect 54908 4338 54964 4340
rect 54908 4286 54910 4338
rect 54910 4286 54962 4338
rect 54962 4286 54964 4338
rect 54908 4284 54964 4286
rect 54124 1596 54180 1652
rect 55244 1372 55300 1428
rect 57484 4450 57540 4452
rect 57484 4398 57486 4450
rect 57486 4398 57538 4450
rect 57538 4398 57540 4450
rect 57484 4396 57540 4398
rect 56700 4338 56756 4340
rect 56700 4286 56702 4338
rect 56702 4286 56754 4338
rect 56754 4286 56756 4338
rect 56700 4284 56756 4286
rect 57708 4338 57764 4340
rect 57708 4286 57710 4338
rect 57710 4286 57762 4338
rect 57762 4286 57764 4338
rect 57708 4284 57764 4286
rect 58828 18508 58884 18564
rect 58716 16940 58772 16996
rect 58940 16828 58996 16884
rect 59388 13132 59444 13188
rect 58940 12348 58996 12404
rect 58828 8316 58884 8372
rect 58716 7980 58772 8036
rect 58604 4172 58660 4228
rect 56700 2716 56756 2772
<< metal3 >>
rect 6066 58492 6076 58548
rect 6132 58492 38220 58548
rect 38276 58492 38286 58548
rect 2594 58380 2604 58436
rect 2660 58380 13356 58436
rect 13412 58380 13422 58436
rect 7858 58268 7868 58324
rect 7924 58268 40124 58324
rect 40180 58268 40190 58324
rect 10882 58156 10892 58212
rect 10948 58156 33852 58212
rect 33908 58156 33918 58212
rect 1362 58044 1372 58100
rect 1428 58044 2268 58100
rect 2324 58044 21868 58100
rect 21924 58044 21934 58100
rect 7522 57932 7532 57988
rect 7588 57932 42812 57988
rect 42868 57932 42878 57988
rect 7410 57820 7420 57876
rect 7476 57820 13692 57876
rect 13748 57820 13758 57876
rect 16370 57820 16380 57876
rect 16436 57820 38668 57876
rect 38724 57820 38734 57876
rect 13234 57708 13244 57764
rect 13300 57708 39228 57764
rect 39284 57708 39294 57764
rect 9314 57596 9324 57652
rect 9380 57596 38332 57652
rect 38388 57596 38398 57652
rect 7858 57484 7868 57540
rect 7924 57484 21308 57540
rect 21364 57484 21374 57540
rect 4610 57372 4620 57428
rect 4676 57372 13916 57428
rect 13972 57372 14924 57428
rect 14980 57372 14990 57428
rect 6626 57260 6636 57316
rect 6692 57260 13468 57316
rect 13524 57260 13534 57316
rect 13682 57260 13692 57316
rect 13748 57260 40684 57316
rect 40740 57260 40750 57316
rect 59200 57204 59800 57232
rect 5842 57148 5852 57204
rect 5908 57148 14812 57204
rect 14868 57148 14878 57204
rect 15026 57148 15036 57204
rect 15092 57148 25900 57204
rect 25956 57148 25966 57204
rect 55794 57148 55804 57204
rect 55860 57148 59800 57204
rect 59200 57120 59800 57148
rect 12786 56700 12796 56756
rect 12852 56700 33628 56756
rect 33684 56700 33694 56756
rect 14914 56588 14924 56644
rect 14980 56588 32956 56644
rect 33012 56588 33022 56644
rect 13458 56476 13468 56532
rect 13524 56476 17388 56532
rect 17444 56476 17454 56532
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 21858 56364 21868 56420
rect 21924 56364 30548 56420
rect 31200 56364 31276 56420
rect 31332 56364 36540 56420
rect 36596 56364 38780 56420
rect 38836 56364 38846 56420
rect 30492 56308 30548 56364
rect 9202 56252 9212 56308
rect 9268 56252 26460 56308
rect 26516 56252 26526 56308
rect 27458 56252 27468 56308
rect 27524 56252 28924 56308
rect 28980 56252 30268 56308
rect 30324 56252 30334 56308
rect 30492 56252 31948 56308
rect 33618 56252 33628 56308
rect 33684 56252 39452 56308
rect 39508 56252 39518 56308
rect 31892 56196 31948 56252
rect 5954 56140 5964 56196
rect 6020 56140 14140 56196
rect 14196 56140 14206 56196
rect 22540 56140 26124 56196
rect 26180 56140 26572 56196
rect 26628 56140 26638 56196
rect 31892 56140 43596 56196
rect 43652 56140 43662 56196
rect 46386 56140 46396 56196
rect 46452 56140 47292 56196
rect 47348 56140 47358 56196
rect 22540 56084 22596 56140
rect 6524 56028 10444 56084
rect 10500 56028 10510 56084
rect 10658 56028 10668 56084
rect 10724 56028 14028 56084
rect 14084 56028 17500 56084
rect 17556 56028 17566 56084
rect 18470 56028 18508 56084
rect 18564 56028 18574 56084
rect 21634 56028 21644 56084
rect 21700 56028 22540 56084
rect 22596 56028 22606 56084
rect 24434 56028 24444 56084
rect 24500 56028 25676 56084
rect 25732 56028 25742 56084
rect 31948 56028 34412 56084
rect 34468 56028 34478 56084
rect 47506 56028 47516 56084
rect 47572 56028 52780 56084
rect 52836 56028 52846 56084
rect 6524 55972 6580 56028
rect 1250 55916 1260 55972
rect 1316 55916 3052 55972
rect 3108 55916 3118 55972
rect 5058 55916 5068 55972
rect 5124 55916 5404 55972
rect 5460 55916 5470 55972
rect 5618 55916 5628 55972
rect 5684 55916 6076 55972
rect 6132 55916 6142 55972
rect 6486 55916 6524 55972
rect 6580 55916 6590 55972
rect 10098 55916 10108 55972
rect 10164 55916 10220 55972
rect 10276 55916 10286 55972
rect 11106 55916 11116 55972
rect 11172 55916 15708 55972
rect 15764 55916 15774 55972
rect 18162 55916 18172 55972
rect 18228 55916 19068 55972
rect 19124 55916 19134 55972
rect 25778 55916 25788 55972
rect 25844 55916 29260 55972
rect 29316 55916 29326 55972
rect 200 55860 800 55888
rect 200 55804 1932 55860
rect 1988 55804 1998 55860
rect 8978 55804 8988 55860
rect 9044 55804 11676 55860
rect 11732 55804 11742 55860
rect 14130 55804 14140 55860
rect 14196 55804 16940 55860
rect 16996 55804 17006 55860
rect 17938 55804 17948 55860
rect 18004 55804 18452 55860
rect 22642 55804 22652 55860
rect 22708 55804 24892 55860
rect 24948 55804 24958 55860
rect 200 55776 800 55804
rect 5506 55692 5516 55748
rect 5572 55692 10668 55748
rect 10724 55692 10734 55748
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 18396 55636 18452 55804
rect 31948 55636 32004 56028
rect 32162 55916 32172 55972
rect 32228 55916 33292 55972
rect 33348 55916 36988 55972
rect 37044 55916 37054 55972
rect 39778 55916 39788 55972
rect 39844 55916 40236 55972
rect 40292 55916 42364 55972
rect 42420 55916 42430 55972
rect 51762 55916 51772 55972
rect 51828 55916 53452 55972
rect 53508 55916 53518 55972
rect 5170 55580 5180 55636
rect 5236 55580 17836 55636
rect 17892 55580 17902 55636
rect 18386 55580 18396 55636
rect 18452 55580 19852 55636
rect 19908 55580 19918 55636
rect 26002 55580 26012 55636
rect 26068 55580 32004 55636
rect 32620 55804 43484 55860
rect 43540 55804 43550 55860
rect 32620 55524 32676 55804
rect 37986 55692 37996 55748
rect 38052 55692 41804 55748
rect 41860 55692 41870 55748
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 42802 55580 42812 55636
rect 42868 55580 43932 55636
rect 43988 55580 43998 55636
rect 9762 55468 9772 55524
rect 9828 55468 11732 55524
rect 16818 55468 16828 55524
rect 16884 55468 19516 55524
rect 19572 55468 19582 55524
rect 26562 55468 26572 55524
rect 26628 55468 32676 55524
rect 33058 55468 33068 55524
rect 33124 55468 39116 55524
rect 39172 55468 39182 55524
rect 11676 55412 11732 55468
rect 11676 55356 12908 55412
rect 12964 55356 12974 55412
rect 23538 55356 23548 55412
rect 23604 55356 28476 55412
rect 28532 55356 28542 55412
rect 30594 55356 30604 55412
rect 30660 55356 32172 55412
rect 32228 55356 32238 55412
rect 32386 55356 32396 55412
rect 32452 55356 33964 55412
rect 34020 55356 34030 55412
rect 44594 55356 44604 55412
rect 44660 55356 45836 55412
rect 45892 55356 45902 55412
rect 56018 55356 56028 55412
rect 56084 55356 57148 55412
rect 57204 55356 57214 55412
rect 2790 55244 2828 55300
rect 2884 55244 2894 55300
rect 4162 55244 4172 55300
rect 4228 55244 6860 55300
rect 6916 55244 6926 55300
rect 15138 55244 15148 55300
rect 15204 55244 16156 55300
rect 16212 55244 16222 55300
rect 21074 55244 21084 55300
rect 21140 55244 23884 55300
rect 23940 55244 24220 55300
rect 24276 55244 24286 55300
rect 25218 55244 25228 55300
rect 25284 55244 28252 55300
rect 28308 55244 29932 55300
rect 29988 55244 29998 55300
rect 30146 55244 30156 55300
rect 30212 55244 34300 55300
rect 34356 55244 34366 55300
rect 38882 55244 38892 55300
rect 38948 55244 39564 55300
rect 39620 55244 40012 55300
rect 40068 55244 40078 55300
rect 43138 55244 43148 55300
rect 43204 55244 44492 55300
rect 44548 55244 44558 55300
rect 24220 55188 24276 55244
rect 5058 55132 5068 55188
rect 5124 55132 9436 55188
rect 9492 55132 9884 55188
rect 9940 55132 9950 55188
rect 12114 55132 12124 55188
rect 12180 55132 14924 55188
rect 14980 55132 14990 55188
rect 15082 55132 15092 55188
rect 15148 55132 15596 55188
rect 15652 55132 15662 55188
rect 16594 55132 16604 55188
rect 16660 55132 17276 55188
rect 17332 55132 19180 55188
rect 19236 55132 19246 55188
rect 22194 55132 22204 55188
rect 22260 55132 23436 55188
rect 23492 55132 23502 55188
rect 24220 55132 25340 55188
rect 25396 55132 26236 55188
rect 26292 55132 26302 55188
rect 28476 55132 30156 55188
rect 30212 55132 30222 55188
rect 30594 55132 30604 55188
rect 30660 55132 31164 55188
rect 31220 55132 31230 55188
rect 36082 55132 36092 55188
rect 36148 55132 42476 55188
rect 42532 55132 42542 55188
rect 46610 55132 46620 55188
rect 46676 55132 47180 55188
rect 47236 55132 47246 55188
rect 28476 55076 28532 55132
rect 6738 55020 6748 55076
rect 6804 55020 10108 55076
rect 10164 55020 14140 55076
rect 14196 55020 14206 55076
rect 14802 55020 14812 55076
rect 14868 55020 16380 55076
rect 16436 55020 16446 55076
rect 18386 55020 18396 55076
rect 18452 55020 19404 55076
rect 19460 55020 22092 55076
rect 22148 55020 22158 55076
rect 22306 55020 22316 55076
rect 22372 55020 22410 55076
rect 23202 55020 23212 55076
rect 23268 55020 28476 55076
rect 28532 55020 28542 55076
rect 30034 55020 30044 55076
rect 30100 55020 30716 55076
rect 30772 55020 31388 55076
rect 31444 55020 31454 55076
rect 35186 55020 35196 55076
rect 35252 55020 35868 55076
rect 35924 55020 36988 55076
rect 37044 55020 38444 55076
rect 38500 55020 38510 55076
rect 39890 55020 39900 55076
rect 39956 55020 41244 55076
rect 41300 55020 41310 55076
rect 43026 55020 43036 55076
rect 43092 55020 43372 55076
rect 43428 55020 44716 55076
rect 44772 55020 44782 55076
rect 22316 54964 22372 55020
rect 8642 54908 8652 54964
rect 8708 54908 9772 54964
rect 9828 54908 12796 54964
rect 12852 54908 12862 54964
rect 13122 54908 13132 54964
rect 13188 54908 17164 54964
rect 17220 54908 17230 54964
rect 20850 54908 20860 54964
rect 20916 54908 22764 54964
rect 22820 54908 23324 54964
rect 23380 54908 23548 54964
rect 26842 54908 26852 54964
rect 26908 54908 27916 54964
rect 27972 54908 28588 54964
rect 28644 54908 29708 54964
rect 29764 54908 29774 54964
rect 31154 54908 31164 54964
rect 31220 54908 31612 54964
rect 31668 54908 32172 54964
rect 32228 54908 32620 54964
rect 32676 54908 47068 54964
rect 47124 54908 47134 54964
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 23492 54852 23548 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 6290 54796 6300 54852
rect 6356 54796 8876 54852
rect 8932 54796 18172 54852
rect 18228 54796 18238 54852
rect 23492 54796 23660 54852
rect 23716 54796 27132 54852
rect 27188 54796 27198 54852
rect 3938 54684 3948 54740
rect 4004 54684 8540 54740
rect 8596 54684 11452 54740
rect 11508 54684 11518 54740
rect 12226 54684 12236 54740
rect 12292 54684 13132 54740
rect 13188 54684 13198 54740
rect 14662 54684 14700 54740
rect 14756 54684 14766 54740
rect 15138 54684 15148 54740
rect 15204 54684 20412 54740
rect 20468 54684 20478 54740
rect 22194 54684 22204 54740
rect 22260 54684 26908 54740
rect 27234 54684 27244 54740
rect 27300 54684 30156 54740
rect 30212 54684 30222 54740
rect 30930 54684 30940 54740
rect 30996 54684 31612 54740
rect 31668 54684 31678 54740
rect 36194 54684 36204 54740
rect 36260 54684 39340 54740
rect 39396 54684 40348 54740
rect 40404 54684 40414 54740
rect 42242 54684 42252 54740
rect 42308 54684 45836 54740
rect 45892 54684 45902 54740
rect 10322 54572 10332 54628
rect 10388 54572 11004 54628
rect 11060 54572 11070 54628
rect 12450 54572 12460 54628
rect 12516 54572 18284 54628
rect 18340 54572 18350 54628
rect 19058 54572 19068 54628
rect 19124 54572 24444 54628
rect 24500 54572 24510 54628
rect 25228 54572 26684 54628
rect 26740 54572 26750 54628
rect 26852 54572 26908 54684
rect 26964 54572 27692 54628
rect 27748 54572 27758 54628
rect 28924 54572 34636 54628
rect 34692 54572 34702 54628
rect 37762 54572 37772 54628
rect 37828 54572 38780 54628
rect 38836 54572 38846 54628
rect 42130 54572 42140 54628
rect 42196 54572 43708 54628
rect 43764 54572 44156 54628
rect 44212 54572 44222 54628
rect 3714 54460 3724 54516
rect 3780 54460 12684 54516
rect 12740 54460 12750 54516
rect 14130 54460 14140 54516
rect 14196 54460 15932 54516
rect 15988 54460 15998 54516
rect 16482 54460 16492 54516
rect 16548 54460 20748 54516
rect 20804 54460 20814 54516
rect 22082 54460 22092 54516
rect 22148 54460 23996 54516
rect 24052 54460 24556 54516
rect 24612 54460 25004 54516
rect 25060 54460 25070 54516
rect 15932 54404 15988 54460
rect 25228 54404 25284 54572
rect 26758 54460 26796 54516
rect 26852 54460 26862 54516
rect 2482 54348 2492 54404
rect 2548 54348 3388 54404
rect 3826 54348 3836 54404
rect 3892 54348 8204 54404
rect 8260 54348 8270 54404
rect 9090 54348 9100 54404
rect 9156 54348 9772 54404
rect 9828 54348 9838 54404
rect 11106 54348 11116 54404
rect 11172 54348 13132 54404
rect 13188 54348 13804 54404
rect 13860 54348 14812 54404
rect 14868 54348 14878 54404
rect 15932 54348 16716 54404
rect 16772 54348 16782 54404
rect 17154 54348 17164 54404
rect 17220 54348 19348 54404
rect 21298 54348 21308 54404
rect 21364 54348 21868 54404
rect 21924 54348 25284 54404
rect 26674 54348 26684 54404
rect 26740 54348 28700 54404
rect 28756 54348 28766 54404
rect 3332 54292 3388 54348
rect 19292 54292 19348 54348
rect 28924 54292 28980 54572
rect 33842 54460 33852 54516
rect 33908 54460 34356 54516
rect 39330 54460 39340 54516
rect 39396 54460 42028 54516
rect 42084 54460 43596 54516
rect 43652 54460 43662 54516
rect 34300 54404 34356 54460
rect 29138 54348 29148 54404
rect 29204 54348 29932 54404
rect 29988 54348 30940 54404
rect 30996 54348 31006 54404
rect 31266 54348 31276 54404
rect 31332 54348 34076 54404
rect 34132 54348 34142 54404
rect 34300 54348 40180 54404
rect 40124 54292 40180 54348
rect 3332 54236 9996 54292
rect 10052 54236 10062 54292
rect 13010 54236 13020 54292
rect 13076 54236 15372 54292
rect 15428 54236 15438 54292
rect 17378 54236 17388 54292
rect 17444 54236 17948 54292
rect 18004 54236 18014 54292
rect 18162 54236 18172 54292
rect 18228 54236 18266 54292
rect 18610 54236 18620 54292
rect 18676 54236 19068 54292
rect 19124 54236 19134 54292
rect 19292 54236 28980 54292
rect 30482 54236 30492 54292
rect 30548 54236 34188 54292
rect 34244 54236 34860 54292
rect 34916 54236 34926 54292
rect 35970 54236 35980 54292
rect 36036 54236 36988 54292
rect 37044 54236 37054 54292
rect 40114 54236 40124 54292
rect 40180 54236 40190 54292
rect 41122 54236 41132 54292
rect 41188 54236 43596 54292
rect 43652 54236 44044 54292
rect 44100 54236 44110 54292
rect 17948 54180 18004 54236
rect 5954 54124 5964 54180
rect 6020 54124 6524 54180
rect 6580 54124 13692 54180
rect 13748 54124 13758 54180
rect 17948 54124 21644 54180
rect 21700 54124 21710 54180
rect 41458 54124 41468 54180
rect 41524 54124 43148 54180
rect 43204 54124 43708 54180
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 13692 54068 13748 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 43652 54068 43708 54124
rect 5058 54012 5068 54068
rect 5124 54012 5516 54068
rect 5572 54012 5582 54068
rect 7970 54012 7980 54068
rect 8036 54012 8204 54068
rect 8260 54012 8270 54068
rect 9874 54012 9884 54068
rect 9940 54012 10556 54068
rect 10612 54012 10622 54068
rect 13692 54012 18732 54068
rect 18788 54012 18844 54068
rect 18900 54012 18910 54068
rect 25442 54012 25452 54068
rect 25508 54012 33404 54068
rect 33460 54012 33470 54068
rect 43652 54012 45724 54068
rect 45780 54012 45790 54068
rect 6962 53900 6972 53956
rect 7028 53900 8316 53956
rect 8372 53900 8382 53956
rect 9426 53900 9436 53956
rect 9492 53900 16156 53956
rect 16212 53900 16222 53956
rect 16370 53900 16380 53956
rect 16436 53900 23436 53956
rect 23492 53900 28700 53956
rect 28756 53900 28766 53956
rect 28914 53900 28924 53956
rect 28980 53900 30604 53956
rect 30660 53900 30670 53956
rect 33954 53900 33964 53956
rect 34020 53900 42140 53956
rect 42196 53900 42206 53956
rect 3378 53788 3388 53844
rect 3444 53788 5628 53844
rect 5684 53788 5694 53844
rect 8352 53788 8428 53844
rect 8484 53788 9100 53844
rect 9156 53788 9166 53844
rect 10770 53788 10780 53844
rect 10836 53788 14756 53844
rect 17826 53788 17836 53844
rect 17892 53788 23100 53844
rect 23156 53788 23166 53844
rect 23492 53788 25004 53844
rect 25060 53788 25452 53844
rect 25508 53788 25518 53844
rect 26562 53788 26572 53844
rect 26628 53788 27020 53844
rect 27076 53788 28028 53844
rect 28084 53788 28094 53844
rect 30370 53788 30380 53844
rect 30436 53788 30828 53844
rect 30884 53788 31164 53844
rect 31220 53788 31230 53844
rect 34626 53788 34636 53844
rect 34692 53788 37044 53844
rect 37426 53788 37436 53844
rect 37492 53788 39788 53844
rect 39844 53788 39854 53844
rect 49522 53788 49532 53844
rect 49588 53788 53900 53844
rect 53956 53788 53966 53844
rect 14700 53732 14756 53788
rect 23492 53732 23548 53788
rect 36988 53732 37044 53788
rect 3490 53676 3500 53732
rect 3556 53676 5740 53732
rect 5796 53676 6076 53732
rect 6132 53676 6142 53732
rect 6626 53676 6636 53732
rect 6692 53676 7756 53732
rect 7812 53676 7822 53732
rect 12674 53676 12684 53732
rect 12740 53676 14532 53732
rect 14690 53676 14700 53732
rect 14756 53676 14812 53732
rect 14868 53676 14878 53732
rect 15586 53676 15596 53732
rect 15652 53676 15820 53732
rect 15876 53676 17108 53732
rect 18274 53676 18284 53732
rect 18340 53676 19964 53732
rect 20020 53676 23548 53732
rect 24098 53676 24108 53732
rect 24164 53676 25676 53732
rect 25732 53676 25742 53732
rect 28354 53676 28364 53732
rect 28420 53676 30156 53732
rect 30212 53676 30222 53732
rect 31938 53676 31948 53732
rect 32004 53676 33404 53732
rect 33460 53676 33470 53732
rect 36988 53676 37324 53732
rect 37380 53676 40012 53732
rect 40068 53676 40078 53732
rect 14476 53620 14532 53676
rect 1810 53564 1820 53620
rect 1876 53564 6524 53620
rect 6580 53564 6590 53620
rect 6738 53564 6748 53620
rect 6804 53564 7644 53620
rect 7700 53564 7710 53620
rect 13458 53564 13468 53620
rect 13524 53564 13804 53620
rect 13860 53564 13870 53620
rect 14476 53564 16884 53620
rect 6748 53508 6804 53564
rect 2258 53452 2268 53508
rect 2324 53452 3948 53508
rect 4004 53452 4014 53508
rect 5170 53452 5180 53508
rect 5236 53452 6804 53508
rect 7970 53452 7980 53508
rect 8036 53452 8876 53508
rect 8932 53452 8942 53508
rect 12534 53452 12572 53508
rect 12628 53452 12638 53508
rect 14130 53452 14140 53508
rect 14196 53452 14476 53508
rect 14532 53452 15260 53508
rect 15316 53452 16268 53508
rect 16324 53452 16334 53508
rect 16828 53396 16884 53564
rect 17052 53508 17108 53676
rect 18274 53564 18284 53620
rect 18340 53564 18844 53620
rect 18900 53564 18910 53620
rect 19618 53564 19628 53620
rect 19684 53564 22428 53620
rect 22484 53564 23044 53620
rect 23426 53564 23436 53620
rect 23492 53564 23996 53620
rect 24052 53564 25004 53620
rect 25060 53564 25070 53620
rect 26562 53564 26572 53620
rect 26628 53564 27356 53620
rect 27412 53564 27422 53620
rect 39890 53564 39900 53620
rect 39956 53564 40908 53620
rect 40964 53564 40974 53620
rect 22988 53508 23044 53564
rect 17042 53452 17052 53508
rect 17108 53452 17118 53508
rect 19170 53452 19180 53508
rect 19236 53452 22764 53508
rect 22820 53452 22830 53508
rect 22988 53452 24556 53508
rect 24612 53452 24622 53508
rect 34738 53452 34748 53508
rect 34804 53452 35644 53508
rect 35700 53452 36876 53508
rect 36932 53452 36942 53508
rect 43596 53452 44044 53508
rect 44100 53452 44492 53508
rect 44548 53452 44558 53508
rect 2034 53340 2044 53396
rect 2100 53340 7980 53396
rect 8036 53340 8046 53396
rect 13356 53340 14588 53396
rect 14644 53340 16380 53396
rect 16436 53340 16446 53396
rect 16828 53340 19628 53396
rect 19684 53340 19694 53396
rect 22978 53340 22988 53396
rect 23044 53340 30828 53396
rect 30884 53340 30894 53396
rect 33394 53340 33404 53396
rect 33460 53340 33740 53396
rect 33796 53340 34412 53396
rect 34468 53340 35084 53396
rect 35140 53340 36092 53396
rect 36148 53340 36764 53396
rect 36820 53340 37324 53396
rect 37380 53340 37660 53396
rect 37716 53340 37726 53396
rect 1474 53228 1484 53284
rect 1540 53228 2716 53284
rect 2772 53228 2782 53284
rect 3490 53228 3500 53284
rect 3556 53228 11676 53284
rect 11732 53228 11742 53284
rect 13356 53172 13412 53340
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 43596 53284 43652 53452
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 15138 53228 15148 53284
rect 15204 53228 17500 53284
rect 17556 53228 17566 53284
rect 27906 53228 27916 53284
rect 27972 53228 32452 53284
rect 32722 53228 32732 53284
rect 32788 53228 43036 53284
rect 43092 53228 43596 53284
rect 43652 53228 43662 53284
rect 2482 53116 2492 53172
rect 2548 53116 3612 53172
rect 3668 53116 5628 53172
rect 5684 53116 5694 53172
rect 6178 53116 6188 53172
rect 6244 53116 6300 53172
rect 6356 53116 8092 53172
rect 8148 53116 8158 53172
rect 9986 53116 9996 53172
rect 10052 53116 13356 53172
rect 13412 53116 13422 53172
rect 14354 53116 14364 53172
rect 14420 53116 15036 53172
rect 15092 53116 15102 53172
rect 16818 53116 16828 53172
rect 16884 53116 17948 53172
rect 18004 53116 18396 53172
rect 18452 53116 20524 53172
rect 20580 53116 20590 53172
rect 20962 53116 20972 53172
rect 21028 53116 23548 53172
rect 23604 53116 23996 53172
rect 24052 53116 24062 53172
rect 26786 53116 26796 53172
rect 26852 53116 31948 53172
rect 32004 53116 32014 53172
rect 4274 53004 4284 53060
rect 4340 53004 9884 53060
rect 9940 53004 9950 53060
rect 13010 53004 13020 53060
rect 13076 53004 14588 53060
rect 14644 53004 14654 53060
rect 14802 53004 14812 53060
rect 14868 53004 16716 53060
rect 16772 53004 25340 53060
rect 25396 53004 25406 53060
rect 26114 53004 26124 53060
rect 26180 53004 27916 53060
rect 27972 53004 27982 53060
rect 5954 52892 5964 52948
rect 6020 52892 6972 52948
rect 7028 52892 7196 52948
rect 7252 52892 7262 52948
rect 8194 52892 8204 52948
rect 8260 52892 8876 52948
rect 8932 52892 8942 52948
rect 11218 52892 11228 52948
rect 11284 52892 12572 52948
rect 12628 52892 12638 52948
rect 13094 52892 13132 52948
rect 13188 52892 13198 52948
rect 14690 52892 14700 52948
rect 14756 52892 15148 52948
rect 15204 52892 15214 52948
rect 15708 52892 18564 52948
rect 20626 52892 20636 52948
rect 20692 52892 21196 52948
rect 21252 52892 21262 52948
rect 26674 52892 26684 52948
rect 26740 52892 27804 52948
rect 27860 52892 27870 52948
rect 1362 52780 1372 52836
rect 1428 52780 2156 52836
rect 2212 52780 2222 52836
rect 3154 52780 3164 52836
rect 3220 52780 6300 52836
rect 6356 52780 6366 52836
rect 7746 52780 7756 52836
rect 7812 52780 10220 52836
rect 10276 52780 10286 52836
rect 14354 52780 14364 52836
rect 14420 52780 15148 52836
rect 15204 52780 15214 52836
rect 10220 52724 10276 52780
rect 2940 52668 8540 52724
rect 8596 52668 8606 52724
rect 10220 52668 14700 52724
rect 14756 52668 14766 52724
rect 2940 52612 2996 52668
rect 15708 52612 15764 52892
rect 15922 52780 15932 52836
rect 15988 52780 16156 52836
rect 16212 52780 16222 52836
rect 16454 52780 16492 52836
rect 16548 52780 16558 52836
rect 18508 52724 18564 52892
rect 20178 52780 20188 52836
rect 20244 52780 21420 52836
rect 21476 52780 21486 52836
rect 22418 52780 22428 52836
rect 22484 52780 23100 52836
rect 23156 52780 23166 52836
rect 23314 52780 23324 52836
rect 23380 52780 24780 52836
rect 24836 52780 24846 52836
rect 26450 52780 26460 52836
rect 26516 52780 26796 52836
rect 26852 52780 26862 52836
rect 27010 52780 27020 52836
rect 27076 52780 28476 52836
rect 28532 52780 29372 52836
rect 29428 52780 29438 52836
rect 32396 52724 32452 53228
rect 32610 53116 32620 53172
rect 32676 53116 33740 53172
rect 33796 53116 33806 53172
rect 36754 53116 36764 53172
rect 36820 53116 37772 53172
rect 37828 53116 37838 53172
rect 36530 53004 36540 53060
rect 36596 53004 38220 53060
rect 38276 53004 38286 53060
rect 40786 53004 40796 53060
rect 40852 53004 42476 53060
rect 42532 53004 42542 53060
rect 35970 52892 35980 52948
rect 36036 52892 41580 52948
rect 41636 52892 41646 52948
rect 37426 52780 37436 52836
rect 37492 52780 38668 52836
rect 38724 52780 38734 52836
rect 42354 52780 42364 52836
rect 42420 52780 52892 52836
rect 52948 52780 52958 52836
rect 16604 52668 17500 52724
rect 17556 52668 17566 52724
rect 18498 52668 18508 52724
rect 18564 52668 20300 52724
rect 20356 52668 30268 52724
rect 30324 52668 30334 52724
rect 32396 52668 41580 52724
rect 41636 52668 42476 52724
rect 42532 52668 42542 52724
rect 16604 52612 16660 52668
rect 1810 52556 1820 52612
rect 1876 52556 2940 52612
rect 2996 52556 3006 52612
rect 9986 52556 9996 52612
rect 10052 52556 13244 52612
rect 13300 52556 13310 52612
rect 14802 52556 14812 52612
rect 14868 52556 15764 52612
rect 16594 52556 16604 52612
rect 16660 52556 16670 52612
rect 17154 52556 17164 52612
rect 17220 52556 18172 52612
rect 18228 52556 18238 52612
rect 20514 52556 20524 52612
rect 20580 52556 22316 52612
rect 22372 52556 22382 52612
rect 27132 52556 28924 52612
rect 28980 52556 28990 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 27132 52500 27188 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 7186 52444 7196 52500
rect 7252 52444 15092 52500
rect 15036 52388 15092 52444
rect 15596 52444 17724 52500
rect 17780 52444 17790 52500
rect 17938 52444 17948 52500
rect 18004 52444 18844 52500
rect 18900 52444 18910 52500
rect 20066 52444 20076 52500
rect 20132 52444 24108 52500
rect 24164 52444 24174 52500
rect 25890 52444 25900 52500
rect 25956 52444 26460 52500
rect 26516 52444 27132 52500
rect 27188 52444 27198 52500
rect 27458 52444 27468 52500
rect 27524 52444 33404 52500
rect 33460 52444 33470 52500
rect 15596 52388 15652 52444
rect 8194 52332 8204 52388
rect 8260 52332 11900 52388
rect 11956 52332 11966 52388
rect 12460 52332 12796 52388
rect 12852 52332 12862 52388
rect 13010 52332 13020 52388
rect 13076 52332 13244 52388
rect 13300 52332 13310 52388
rect 15026 52332 15036 52388
rect 15092 52332 15596 52388
rect 15652 52332 15662 52388
rect 16930 52332 16940 52388
rect 16996 52332 18396 52388
rect 18452 52332 18462 52388
rect 19366 52332 19404 52388
rect 19460 52332 19470 52388
rect 25218 52332 25228 52388
rect 25284 52332 26684 52388
rect 26740 52332 26750 52388
rect 30706 52332 30716 52388
rect 30772 52332 37548 52388
rect 37604 52332 37614 52388
rect 44706 52332 44716 52388
rect 44772 52332 46060 52388
rect 46116 52332 46126 52388
rect 12460 52276 12516 52332
rect 1138 52220 1148 52276
rect 1204 52220 2604 52276
rect 2660 52220 2670 52276
rect 5170 52220 5180 52276
rect 5236 52220 5852 52276
rect 5908 52220 6524 52276
rect 6580 52220 6590 52276
rect 6962 52220 6972 52276
rect 7028 52220 9436 52276
rect 9492 52220 10892 52276
rect 10948 52220 10958 52276
rect 12114 52220 12124 52276
rect 12180 52220 12460 52276
rect 12516 52220 12526 52276
rect 12674 52220 12684 52276
rect 12740 52220 12778 52276
rect 12898 52220 12908 52276
rect 12964 52220 20524 52276
rect 20580 52220 20590 52276
rect 23538 52220 23548 52276
rect 23604 52220 29820 52276
rect 29876 52220 29886 52276
rect 32050 52220 32060 52276
rect 32116 52220 33292 52276
rect 33348 52220 34412 52276
rect 34468 52220 34478 52276
rect 35858 52220 35868 52276
rect 35924 52220 42252 52276
rect 42308 52220 42318 52276
rect 3266 52108 3276 52164
rect 3332 52108 6972 52164
rect 7028 52108 7038 52164
rect 7522 52108 7532 52164
rect 7588 52108 8092 52164
rect 8148 52108 8158 52164
rect 9090 52108 9100 52164
rect 9156 52108 14700 52164
rect 14756 52108 14766 52164
rect 16304 52108 16380 52164
rect 16436 52108 20188 52164
rect 20244 52108 20636 52164
rect 20692 52108 20702 52164
rect 20850 52108 20860 52164
rect 20916 52108 23660 52164
rect 23716 52108 23726 52164
rect 24098 52108 24108 52164
rect 24164 52108 24556 52164
rect 24612 52108 24622 52164
rect 24994 52108 25004 52164
rect 25060 52108 26404 52164
rect 26562 52108 26572 52164
rect 26628 52108 27692 52164
rect 27748 52108 27758 52164
rect 28588 52108 35532 52164
rect 35588 52108 36764 52164
rect 36820 52108 36830 52164
rect 40450 52108 40460 52164
rect 40516 52108 41356 52164
rect 41412 52108 41422 52164
rect 43922 52108 43932 52164
rect 43988 52108 45388 52164
rect 45444 52108 45454 52164
rect 48738 52108 48748 52164
rect 48804 52108 54908 52164
rect 54964 52108 54974 52164
rect 26348 52052 26404 52108
rect 2706 51996 2716 52052
rect 2772 51996 5068 52052
rect 5124 51996 5134 52052
rect 6626 51996 6636 52052
rect 6692 51996 8204 52052
rect 8260 51996 8270 52052
rect 11442 51996 11452 52052
rect 11508 51996 12572 52052
rect 12628 51996 16268 52052
rect 16324 51996 16334 52052
rect 16482 51996 16492 52052
rect 16548 51996 16828 52052
rect 16884 51996 17164 52052
rect 17220 51996 17230 52052
rect 19170 51996 19180 52052
rect 19236 51996 19852 52052
rect 19908 51996 19918 52052
rect 22866 51996 22876 52052
rect 22932 51996 24668 52052
rect 24724 51996 24734 52052
rect 24882 51996 24892 52052
rect 24948 51996 25564 52052
rect 25620 51996 26124 52052
rect 26180 51996 26190 52052
rect 26348 51996 27132 52052
rect 27188 51996 27198 52052
rect 28588 51940 28644 52108
rect 31266 51996 31276 52052
rect 31332 51996 31836 52052
rect 31892 51996 32396 52052
rect 32452 51996 32956 52052
rect 33012 51996 33022 52052
rect 37650 51996 37660 52052
rect 37716 51996 38444 52052
rect 38500 51996 38510 52052
rect 41906 51996 41916 52052
rect 41972 51996 42364 52052
rect 42420 51996 42430 52052
rect 44370 51996 44380 52052
rect 44436 51996 46060 52052
rect 46116 51996 46126 52052
rect 1922 51884 1932 51940
rect 1988 51884 2156 51940
rect 2212 51884 2222 51940
rect 5618 51884 5628 51940
rect 5684 51884 6524 51940
rect 6580 51884 7644 51940
rect 7700 51884 12124 51940
rect 12180 51884 12190 51940
rect 12310 51884 12348 51940
rect 12404 51884 12414 51940
rect 15362 51884 15372 51940
rect 15428 51884 15484 51940
rect 15540 51884 16716 51940
rect 16772 51884 16782 51940
rect 18162 51884 18172 51940
rect 18228 51884 22092 51940
rect 22148 51884 22158 51940
rect 23762 51884 23772 51940
rect 23828 51884 28644 51940
rect 38098 51884 38108 51940
rect 38164 51884 38556 51940
rect 38612 51884 38622 51940
rect 43250 51884 43260 51940
rect 43316 51884 44604 51940
rect 44660 51884 45836 51940
rect 45892 51884 45902 51940
rect 59200 51828 59800 51856
rect 5282 51772 5292 51828
rect 5348 51772 5358 51828
rect 7522 51772 7532 51828
rect 7588 51772 9996 51828
rect 10052 51772 10062 51828
rect 11218 51772 11228 51828
rect 11284 51772 13692 51828
rect 13748 51772 13758 51828
rect 14018 51772 14028 51828
rect 14084 51772 14924 51828
rect 14980 51772 14990 51828
rect 15250 51772 15260 51828
rect 15316 51772 15708 51828
rect 15764 51772 16492 51828
rect 16548 51772 16558 51828
rect 18274 51772 18284 51828
rect 18340 51772 19292 51828
rect 19348 51772 19358 51828
rect 21410 51772 21420 51828
rect 21476 51772 21756 51828
rect 21812 51772 22764 51828
rect 22820 51772 23436 51828
rect 23492 51772 23502 51828
rect 25330 51772 25340 51828
rect 25396 51772 26124 51828
rect 26180 51772 26190 51828
rect 27010 51772 27020 51828
rect 27076 51772 27244 51828
rect 27300 51772 27310 51828
rect 32386 51772 32396 51828
rect 32452 51772 33068 51828
rect 33124 51772 33740 51828
rect 33796 51772 33806 51828
rect 56018 51772 56028 51828
rect 56084 51772 59800 51828
rect 5292 51716 5348 51772
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 59200 51744 59800 51772
rect 5292 51660 5628 51716
rect 5684 51660 5694 51716
rect 6850 51660 6860 51716
rect 6916 51660 7868 51716
rect 7924 51660 7934 51716
rect 9174 51660 9212 51716
rect 9268 51660 9278 51716
rect 11330 51660 11340 51716
rect 11396 51660 13916 51716
rect 13972 51660 13982 51716
rect 16370 51660 16380 51716
rect 16436 51660 16446 51716
rect 20738 51660 20748 51716
rect 20804 51660 31276 51716
rect 31332 51660 31342 51716
rect 33730 51660 33740 51716
rect 33796 51660 40572 51716
rect 40628 51660 40638 51716
rect 4162 51548 4172 51604
rect 4228 51548 5404 51604
rect 5460 51548 5470 51604
rect 5730 51548 5740 51604
rect 5796 51548 6524 51604
rect 6580 51548 6590 51604
rect 7298 51548 7308 51604
rect 7364 51548 9884 51604
rect 9940 51548 9950 51604
rect 11666 51548 11676 51604
rect 11732 51548 11742 51604
rect 12012 51548 12628 51604
rect 11676 51492 11732 51548
rect 12012 51492 12068 51548
rect 12572 51492 12628 51548
rect 16380 51492 16436 51660
rect 16706 51548 16716 51604
rect 16772 51548 17948 51604
rect 18004 51548 18014 51604
rect 18946 51548 18956 51604
rect 19012 51548 20524 51604
rect 20580 51548 20972 51604
rect 21028 51548 21038 51604
rect 21270 51548 21308 51604
rect 21364 51548 21374 51604
rect 23874 51548 23884 51604
rect 23940 51548 24836 51604
rect 25666 51548 25676 51604
rect 25732 51548 26236 51604
rect 26292 51548 26302 51604
rect 26786 51548 26796 51604
rect 26852 51548 31052 51604
rect 31108 51548 31118 51604
rect 31602 51548 31612 51604
rect 31668 51548 37212 51604
rect 37268 51548 37278 51604
rect 39778 51548 39788 51604
rect 39844 51548 44380 51604
rect 44436 51548 44446 51604
rect 24780 51492 24836 51548
rect 4050 51436 4060 51492
rect 4116 51436 4126 51492
rect 4834 51436 4844 51492
rect 4900 51436 5852 51492
rect 5908 51436 7420 51492
rect 7476 51436 7486 51492
rect 7942 51436 7980 51492
rect 8036 51436 8046 51492
rect 8540 51436 12068 51492
rect 12198 51436 12236 51492
rect 12292 51436 12302 51492
rect 12572 51436 14252 51492
rect 14308 51436 14318 51492
rect 16380 51436 23660 51492
rect 23716 51436 23726 51492
rect 24770 51436 24780 51492
rect 24836 51436 25564 51492
rect 25620 51436 25630 51492
rect 28130 51436 28140 51492
rect 28196 51436 29708 51492
rect 29764 51436 30380 51492
rect 30436 51436 30446 51492
rect 4060 51380 4116 51436
rect 4060 51324 8316 51380
rect 8372 51324 8382 51380
rect 8540 51268 8596 51436
rect 31052 51380 31108 51548
rect 33394 51436 33404 51492
rect 33460 51436 33852 51492
rect 33908 51436 34524 51492
rect 34580 51436 34590 51492
rect 9314 51324 9324 51380
rect 9380 51324 10444 51380
rect 10500 51324 10510 51380
rect 12086 51324 12124 51380
rect 12180 51324 12190 51380
rect 12450 51324 12460 51380
rect 12516 51324 13692 51380
rect 13748 51324 13758 51380
rect 16342 51324 16380 51380
rect 16436 51324 16446 51380
rect 16930 51324 16940 51380
rect 16996 51324 17612 51380
rect 17668 51324 17678 51380
rect 18162 51324 18172 51380
rect 18228 51324 20860 51380
rect 20916 51324 20926 51380
rect 22418 51324 22428 51380
rect 22484 51324 23212 51380
rect 23268 51324 23548 51380
rect 23604 51324 23614 51380
rect 23874 51324 23884 51380
rect 23940 51324 24108 51380
rect 24164 51324 24174 51380
rect 27122 51324 27132 51380
rect 27188 51324 28364 51380
rect 28420 51324 28430 51380
rect 31052 51324 31612 51380
rect 31668 51324 31678 51380
rect 32498 51324 32508 51380
rect 32564 51324 33740 51380
rect 33796 51324 33806 51380
rect 34066 51324 34076 51380
rect 34132 51324 35644 51380
rect 35700 51324 35710 51380
rect 38210 51324 38220 51380
rect 38276 51324 39676 51380
rect 39732 51324 39742 51380
rect 43586 51324 43596 51380
rect 43652 51324 44828 51380
rect 44884 51324 44894 51380
rect 3042 51212 3052 51268
rect 3108 51212 4340 51268
rect 4834 51212 4844 51268
rect 4900 51212 4956 51268
rect 5012 51212 5022 51268
rect 5170 51212 5180 51268
rect 5236 51212 8596 51268
rect 8838 51212 8876 51268
rect 8932 51212 8942 51268
rect 10098 51212 10108 51268
rect 10164 51212 12236 51268
rect 12292 51212 12302 51268
rect 14354 51212 14364 51268
rect 14420 51212 21868 51268
rect 21924 51212 21934 51268
rect 22642 51212 22652 51268
rect 22708 51212 29820 51268
rect 29876 51212 29886 51268
rect 30146 51212 30156 51268
rect 30212 51212 33740 51268
rect 33796 51212 33806 51268
rect 33954 51212 33964 51268
rect 34020 51212 34860 51268
rect 34916 51212 36652 51268
rect 36708 51212 36718 51268
rect 45042 51212 45052 51268
rect 45108 51212 45724 51268
rect 45780 51212 45790 51268
rect 4284 51156 4340 51212
rect 4284 51100 5292 51156
rect 5348 51100 5358 51156
rect 7970 51100 7980 51156
rect 8036 51100 11564 51156
rect 11620 51100 11630 51156
rect 13010 51100 13020 51156
rect 13076 51100 13356 51156
rect 13412 51100 13422 51156
rect 14914 51100 14924 51156
rect 14980 51100 18956 51156
rect 19012 51100 23324 51156
rect 23380 51100 23390 51156
rect 26852 51100 31388 51156
rect 31444 51100 31454 51156
rect 32722 51100 32732 51156
rect 32788 51100 36092 51156
rect 36148 51100 36158 51156
rect 36866 51100 36876 51156
rect 36932 51100 41580 51156
rect 41636 51100 41646 51156
rect 3714 50988 3724 51044
rect 3780 50988 3948 51044
rect 4004 50988 4014 51044
rect 5058 50988 5068 51044
rect 5124 50988 7644 51044
rect 7700 50988 13468 51044
rect 13524 50988 13534 51044
rect 16482 50988 16492 51044
rect 16548 50988 24780 51044
rect 24836 50988 24846 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 3574 50876 3612 50932
rect 3668 50876 3678 50932
rect 5506 50876 5516 50932
rect 5572 50876 8764 50932
rect 8820 50876 9660 50932
rect 9716 50876 10724 50932
rect 11330 50876 11340 50932
rect 11396 50876 12124 50932
rect 12180 50876 12190 50932
rect 13234 50876 13244 50932
rect 13300 50876 13580 50932
rect 13636 50876 13646 50932
rect 16258 50876 16268 50932
rect 16324 50876 19180 50932
rect 19236 50876 20188 50932
rect 20244 50876 20254 50932
rect 21746 50876 21756 50932
rect 21812 50876 22764 50932
rect 22820 50876 22830 50932
rect 23426 50876 23436 50932
rect 23492 50876 23996 50932
rect 24052 50876 24062 50932
rect 10668 50820 10724 50876
rect 26852 50820 26908 51100
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 38098 50876 38108 50932
rect 38164 50876 38174 50932
rect 2258 50764 2268 50820
rect 2324 50764 5796 50820
rect 6402 50764 6412 50820
rect 6468 50764 8204 50820
rect 8260 50764 10444 50820
rect 10500 50764 10510 50820
rect 10668 50764 13804 50820
rect 13860 50764 13870 50820
rect 14354 50764 14364 50820
rect 14420 50764 21532 50820
rect 21588 50764 21598 50820
rect 22306 50764 22316 50820
rect 22372 50764 26908 50820
rect 31938 50764 31948 50820
rect 32004 50764 34188 50820
rect 34244 50764 34254 50820
rect 34514 50764 34524 50820
rect 34580 50764 36540 50820
rect 36596 50764 36606 50820
rect 5740 50708 5796 50764
rect 2370 50652 2380 50708
rect 2436 50652 5516 50708
rect 5572 50652 5582 50708
rect 5740 50652 12012 50708
rect 12068 50652 12078 50708
rect 13010 50652 13020 50708
rect 13076 50652 16940 50708
rect 16996 50652 17006 50708
rect 17826 50652 17836 50708
rect 17892 50652 18396 50708
rect 18452 50652 19404 50708
rect 19460 50652 20076 50708
rect 20132 50652 25340 50708
rect 25396 50652 25406 50708
rect 27570 50652 27580 50708
rect 27636 50652 28812 50708
rect 28868 50652 29932 50708
rect 29988 50652 29998 50708
rect 35522 50652 35532 50708
rect 35588 50652 36428 50708
rect 36484 50652 37436 50708
rect 37492 50652 37502 50708
rect 3014 50540 3052 50596
rect 3108 50540 3118 50596
rect 4274 50540 4284 50596
rect 4340 50540 14028 50596
rect 14084 50540 14094 50596
rect 14242 50540 14252 50596
rect 14308 50540 16156 50596
rect 16212 50540 16222 50596
rect 19618 50540 19628 50596
rect 19684 50540 21644 50596
rect 21700 50540 21710 50596
rect 23548 50540 27356 50596
rect 27412 50540 27422 50596
rect 34514 50540 34524 50596
rect 34580 50540 35196 50596
rect 35252 50540 36204 50596
rect 36260 50540 37324 50596
rect 37380 50540 37390 50596
rect 200 50484 800 50512
rect 23548 50484 23604 50540
rect 38108 50484 38164 50876
rect 200 50428 1932 50484
rect 1988 50428 1998 50484
rect 3154 50428 3164 50484
rect 3220 50428 3836 50484
rect 3892 50428 3902 50484
rect 4284 50428 4396 50484
rect 4452 50428 4462 50484
rect 4992 50428 5068 50484
rect 5124 50428 5796 50484
rect 5954 50428 5964 50484
rect 6020 50428 6748 50484
rect 6804 50428 6814 50484
rect 7410 50428 7420 50484
rect 7476 50428 8092 50484
rect 8148 50428 8158 50484
rect 9090 50428 9100 50484
rect 9156 50428 10108 50484
rect 10164 50428 13356 50484
rect 13412 50428 13422 50484
rect 13570 50428 13580 50484
rect 13636 50428 14252 50484
rect 14308 50428 14318 50484
rect 14578 50428 14588 50484
rect 14644 50428 16212 50484
rect 16930 50428 16940 50484
rect 16996 50428 17388 50484
rect 17444 50428 17454 50484
rect 18246 50428 18284 50484
rect 18340 50428 18350 50484
rect 21298 50428 21308 50484
rect 21364 50428 22540 50484
rect 22596 50428 22876 50484
rect 22932 50428 23604 50484
rect 23874 50428 23884 50484
rect 23940 50428 24892 50484
rect 24948 50428 24958 50484
rect 26982 50428 27020 50484
rect 27076 50428 27086 50484
rect 27794 50428 27804 50484
rect 27860 50428 28476 50484
rect 28532 50428 28542 50484
rect 30594 50428 30604 50484
rect 30660 50428 32172 50484
rect 32228 50428 32238 50484
rect 36530 50428 36540 50484
rect 36596 50428 38332 50484
rect 38388 50428 38398 50484
rect 200 50400 800 50428
rect 4284 50372 4340 50428
rect 5740 50372 5796 50428
rect 16156 50372 16212 50428
rect 3602 50316 3612 50372
rect 3668 50316 4172 50372
rect 4228 50316 4340 50372
rect 4498 50316 4508 50372
rect 4564 50316 4956 50372
rect 5012 50316 5022 50372
rect 5740 50316 5852 50372
rect 5908 50316 5918 50372
rect 7074 50316 7084 50372
rect 7140 50316 7532 50372
rect 7588 50316 7598 50372
rect 8306 50316 8316 50372
rect 8372 50316 9436 50372
rect 9492 50316 9502 50372
rect 11442 50316 11452 50372
rect 11508 50316 14924 50372
rect 14980 50316 14990 50372
rect 15092 50260 15148 50372
rect 15204 50316 15214 50372
rect 16146 50316 16156 50372
rect 16212 50316 16222 50372
rect 16818 50316 16828 50372
rect 16884 50316 17724 50372
rect 17780 50316 17790 50372
rect 18620 50316 25620 50372
rect 25778 50316 25788 50372
rect 25844 50316 26236 50372
rect 26292 50316 28364 50372
rect 28420 50316 29372 50372
rect 29428 50316 29438 50372
rect 31154 50316 31164 50372
rect 31220 50316 31724 50372
rect 31780 50316 32620 50372
rect 32676 50316 32686 50372
rect 4274 50204 4284 50260
rect 4340 50204 4452 50260
rect 6850 50204 6860 50260
rect 6916 50204 8652 50260
rect 8708 50204 11452 50260
rect 11508 50204 11518 50260
rect 11666 50204 11676 50260
rect 11732 50204 15484 50260
rect 15540 50204 15550 50260
rect 4396 50036 4452 50204
rect 16828 50148 16884 50316
rect 4946 50092 4956 50148
rect 5012 50092 9324 50148
rect 9380 50092 9390 50148
rect 12338 50092 12348 50148
rect 12404 50092 14700 50148
rect 14756 50092 14766 50148
rect 15026 50092 15036 50148
rect 15092 50092 16884 50148
rect 18620 50036 18676 50316
rect 25564 50260 25620 50316
rect 23174 50204 23212 50260
rect 23268 50204 23278 50260
rect 25564 50204 25900 50260
rect 25956 50204 25966 50260
rect 37884 50204 38780 50260
rect 38836 50204 39228 50260
rect 39284 50204 39564 50260
rect 39620 50204 39630 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 26114 50092 26124 50148
rect 26180 50092 30156 50148
rect 30212 50092 30222 50148
rect 31266 50092 31276 50148
rect 31332 50092 32060 50148
rect 32116 50092 33292 50148
rect 33348 50092 33358 50148
rect 37884 50036 37940 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 3714 49980 3724 50036
rect 3780 49980 3790 50036
rect 3938 49980 3948 50036
rect 4004 49980 4172 50036
rect 4228 49980 4238 50036
rect 4396 49980 9772 50036
rect 9828 49980 9838 50036
rect 10322 49980 10332 50036
rect 10388 49980 15036 50036
rect 15092 49980 15102 50036
rect 15362 49980 15372 50036
rect 15428 49980 15820 50036
rect 15876 49980 15886 50036
rect 16482 49980 16492 50036
rect 16548 49980 16604 50036
rect 16660 49980 16716 50036
rect 16772 49980 18676 50036
rect 18834 49980 18844 50036
rect 18900 49980 19852 50036
rect 19908 49980 19918 50036
rect 22306 49980 22316 50036
rect 22372 49980 23324 50036
rect 23380 49980 23390 50036
rect 28242 49980 28252 50036
rect 28308 49980 37884 50036
rect 37940 49980 37950 50036
rect 38210 49980 38220 50036
rect 38276 49980 39564 50036
rect 39620 49980 39630 50036
rect 3724 49924 3780 49980
rect 9772 49924 9828 49980
rect 3724 49868 5628 49924
rect 5684 49868 5694 49924
rect 6850 49868 6860 49924
rect 6916 49868 8204 49924
rect 8260 49868 8596 49924
rect 9314 49868 9324 49924
rect 9380 49868 9436 49924
rect 9492 49868 9502 49924
rect 9772 49868 14140 49924
rect 14196 49868 14206 49924
rect 15922 49868 15932 49924
rect 15988 49868 17388 49924
rect 17444 49868 17454 49924
rect 17602 49868 17612 49924
rect 17668 49868 18956 49924
rect 19012 49868 19022 49924
rect 19394 49868 19404 49924
rect 19460 49868 19516 49924
rect 19572 49868 20188 49924
rect 20244 49868 20254 49924
rect 20402 49868 20412 49924
rect 20468 49868 23212 49924
rect 23268 49868 23772 49924
rect 23828 49868 23838 49924
rect 24322 49868 24332 49924
rect 24388 49868 24892 49924
rect 24948 49868 24958 49924
rect 26450 49868 26460 49924
rect 26516 49868 27804 49924
rect 27860 49868 27870 49924
rect 30818 49868 30828 49924
rect 30884 49868 36316 49924
rect 36372 49868 36382 49924
rect 38612 49868 40908 49924
rect 40964 49868 41804 49924
rect 41860 49868 42252 49924
rect 42308 49868 42476 49924
rect 42532 49868 42542 49924
rect 8540 49812 8596 49868
rect 38612 49812 38668 49868
rect 3332 49756 3948 49812
rect 4004 49756 4956 49812
rect 5012 49756 7084 49812
rect 7140 49756 7150 49812
rect 7522 49756 7532 49812
rect 7588 49756 8316 49812
rect 8372 49756 8382 49812
rect 8540 49756 12908 49812
rect 12964 49756 13356 49812
rect 13412 49756 13422 49812
rect 15474 49756 15484 49812
rect 15540 49756 16380 49812
rect 16436 49756 16446 49812
rect 16818 49756 16828 49812
rect 16884 49756 16940 49812
rect 16996 49756 17006 49812
rect 18498 49756 18508 49812
rect 18564 49756 19628 49812
rect 19684 49756 20076 49812
rect 20132 49756 20142 49812
rect 21970 49756 21980 49812
rect 22036 49756 22652 49812
rect 22708 49756 22718 49812
rect 24546 49756 24556 49812
rect 24612 49756 26908 49812
rect 28354 49756 28364 49812
rect 28420 49756 38668 49812
rect 3332 49700 3388 49756
rect 16828 49700 16884 49756
rect 26852 49700 26908 49756
rect 3154 49644 3164 49700
rect 3220 49644 3388 49700
rect 3612 49644 4060 49700
rect 4116 49644 8652 49700
rect 8708 49644 8718 49700
rect 9090 49644 9100 49700
rect 9156 49644 9548 49700
rect 9604 49644 9614 49700
rect 9958 49644 9996 49700
rect 10052 49644 10062 49700
rect 10630 49644 10668 49700
rect 10724 49644 10734 49700
rect 11554 49644 11564 49700
rect 11620 49644 11676 49700
rect 11732 49644 11742 49700
rect 13990 49644 14028 49700
rect 14084 49644 14094 49700
rect 15092 49644 16884 49700
rect 18610 49644 18620 49700
rect 18676 49644 18844 49700
rect 18900 49644 20748 49700
rect 20804 49644 20814 49700
rect 26852 49644 31836 49700
rect 31892 49644 32732 49700
rect 32788 49644 32798 49700
rect 33926 49644 33964 49700
rect 34020 49644 38220 49700
rect 38276 49644 38286 49700
rect 40226 49644 40236 49700
rect 40292 49644 42812 49700
rect 42868 49644 43484 49700
rect 43540 49644 43550 49700
rect 3612 49588 3668 49644
rect 15092 49588 15148 49644
rect 3378 49532 3388 49588
rect 3444 49532 3668 49588
rect 4060 49532 4620 49588
rect 4676 49532 15148 49588
rect 15698 49532 15708 49588
rect 15764 49532 18620 49588
rect 18676 49532 19628 49588
rect 19684 49532 25564 49588
rect 25620 49532 25630 49588
rect 26852 49532 39452 49588
rect 39508 49532 39518 49588
rect 4060 49476 4116 49532
rect 4050 49420 4060 49476
rect 4116 49420 4126 49476
rect 6962 49420 6972 49476
rect 7028 49420 7084 49476
rect 7140 49420 7150 49476
rect 8642 49420 8652 49476
rect 8708 49420 11900 49476
rect 11956 49420 17556 49476
rect 19058 49420 19068 49476
rect 19124 49420 21420 49476
rect 21476 49420 21486 49476
rect 22194 49420 22204 49476
rect 22260 49420 22876 49476
rect 22932 49420 22942 49476
rect 23090 49420 23100 49476
rect 23156 49420 23212 49476
rect 23268 49420 23278 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 17500 49364 17556 49420
rect 5618 49308 5628 49364
rect 5684 49308 11340 49364
rect 11396 49308 11406 49364
rect 14130 49308 14140 49364
rect 14196 49308 16268 49364
rect 16324 49308 16334 49364
rect 17500 49308 18508 49364
rect 18564 49308 18574 49364
rect 19170 49308 19180 49364
rect 19236 49308 19628 49364
rect 19684 49308 21868 49364
rect 21924 49308 21934 49364
rect 22082 49308 22092 49364
rect 22148 49308 24556 49364
rect 24612 49308 24622 49364
rect 3238 49196 3276 49252
rect 3332 49196 3342 49252
rect 3826 49196 3836 49252
rect 3892 49196 4956 49252
rect 5012 49196 5022 49252
rect 6178 49196 6188 49252
rect 6244 49196 6860 49252
rect 6916 49196 6926 49252
rect 7634 49196 7644 49252
rect 7700 49196 8204 49252
rect 8260 49196 8270 49252
rect 9398 49196 9436 49252
rect 9492 49196 9502 49252
rect 10658 49196 10668 49252
rect 10724 49196 12236 49252
rect 12292 49196 12302 49252
rect 14242 49196 14252 49252
rect 14308 49196 21084 49252
rect 21140 49196 21150 49252
rect 22194 49196 22204 49252
rect 22260 49196 25116 49252
rect 25172 49196 25182 49252
rect 26852 49140 26908 49532
rect 28242 49420 28252 49476
rect 28308 49420 28924 49476
rect 28980 49420 28990 49476
rect 36726 49420 36764 49476
rect 36820 49420 36830 49476
rect 38658 49420 38668 49476
rect 38724 49420 40684 49476
rect 40740 49420 40750 49476
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 31126 49196 31164 49252
rect 31220 49196 31230 49252
rect 2818 49084 2828 49140
rect 2884 49084 5964 49140
rect 6020 49084 6076 49140
rect 6132 49084 6142 49140
rect 7942 49084 7980 49140
rect 8036 49084 8046 49140
rect 8978 49084 8988 49140
rect 9044 49084 10108 49140
rect 10164 49084 10174 49140
rect 10322 49084 10332 49140
rect 10388 49084 10780 49140
rect 10836 49084 10846 49140
rect 11330 49084 11340 49140
rect 11396 49084 14364 49140
rect 14420 49084 14430 49140
rect 15092 49084 15596 49140
rect 15652 49084 15662 49140
rect 16930 49084 16940 49140
rect 16996 49084 18620 49140
rect 18676 49084 18686 49140
rect 19394 49084 19404 49140
rect 19460 49084 19964 49140
rect 20020 49084 20030 49140
rect 20178 49084 20188 49140
rect 20244 49084 20282 49140
rect 21522 49084 21532 49140
rect 21588 49084 24108 49140
rect 24164 49084 24174 49140
rect 24630 49084 24668 49140
rect 24724 49084 24734 49140
rect 25340 49084 26908 49140
rect 28242 49084 28252 49140
rect 28308 49084 29036 49140
rect 29092 49084 29102 49140
rect 32722 49084 32732 49140
rect 32788 49084 33852 49140
rect 33908 49084 33918 49140
rect 34962 49084 34972 49140
rect 35028 49084 37100 49140
rect 37156 49084 37166 49140
rect 15092 49028 15148 49084
rect 25340 49028 25396 49084
rect 2706 48972 2716 49028
rect 2772 48972 4060 49028
rect 4116 48972 4844 49028
rect 4900 48972 4910 49028
rect 7074 48972 7084 49028
rect 7140 48972 7644 49028
rect 7700 48972 7710 49028
rect 8306 48972 8316 49028
rect 8372 48972 14140 49028
rect 14196 48972 15148 49028
rect 15698 48972 15708 49028
rect 15764 48972 16156 49028
rect 16212 48972 16222 49028
rect 17714 48972 17724 49028
rect 17780 48972 18508 49028
rect 18564 48972 18574 49028
rect 18834 48972 18844 49028
rect 18900 48972 25340 49028
rect 25396 48972 25406 49028
rect 28914 48972 28924 49028
rect 28980 48972 29372 49028
rect 29428 48972 30604 49028
rect 30660 48972 30670 49028
rect 30930 48972 30940 49028
rect 30996 48972 31836 49028
rect 31892 48972 33068 49028
rect 33124 48972 33516 49028
rect 33572 48972 33582 49028
rect 34178 48972 34188 49028
rect 34244 48972 35084 49028
rect 35140 48972 35150 49028
rect 36306 48972 36316 49028
rect 36372 48972 37772 49028
rect 37828 48972 38108 49028
rect 38164 48972 38174 49028
rect 39778 48972 39788 49028
rect 39844 48972 40124 49028
rect 40180 48972 40460 49028
rect 40516 48972 40526 49028
rect 30604 48916 30660 48972
rect 1810 48860 1820 48916
rect 1876 48860 2044 48916
rect 2100 48860 4732 48916
rect 4788 48860 4798 48916
rect 4956 48860 5068 48916
rect 5124 48860 5134 48916
rect 8530 48860 8540 48916
rect 8596 48860 10556 48916
rect 10612 48860 10622 48916
rect 11638 48860 11676 48916
rect 11732 48860 11742 48916
rect 14354 48860 14364 48916
rect 14420 48860 14924 48916
rect 14980 48860 14990 48916
rect 15810 48860 15820 48916
rect 15876 48860 20748 48916
rect 20804 48860 20814 48916
rect 22306 48860 22316 48916
rect 22372 48860 22652 48916
rect 22708 48860 22718 48916
rect 23090 48860 23100 48916
rect 23156 48860 23212 48916
rect 23268 48860 23436 48916
rect 23492 48860 23502 48916
rect 27010 48860 27020 48916
rect 27076 48860 27468 48916
rect 27524 48860 27534 48916
rect 30604 48860 31500 48916
rect 31556 48860 31566 48916
rect 32610 48860 32620 48916
rect 32676 48860 33180 48916
rect 33236 48860 33246 48916
rect 36978 48860 36988 48916
rect 37044 48860 40236 48916
rect 40292 48860 40302 48916
rect 41122 48860 41132 48916
rect 41188 48860 42700 48916
rect 42756 48860 43484 48916
rect 43540 48860 43550 48916
rect 45154 48860 45164 48916
rect 45220 48860 45612 48916
rect 45668 48860 45678 48916
rect 47394 48860 47404 48916
rect 47460 48860 58156 48916
rect 58212 48860 58222 48916
rect 4956 48804 5012 48860
rect 3042 48748 3052 48804
rect 3108 48748 3220 48804
rect 3686 48748 3724 48804
rect 3780 48748 3790 48804
rect 4610 48748 4620 48804
rect 4676 48748 5012 48804
rect 5068 48748 10780 48804
rect 10836 48748 10846 48804
rect 12450 48748 12460 48804
rect 12516 48748 16044 48804
rect 16100 48748 16110 48804
rect 18610 48748 18620 48804
rect 18676 48748 20300 48804
rect 20356 48748 20366 48804
rect 22502 48748 22540 48804
rect 22596 48748 22606 48804
rect 23202 48748 23212 48804
rect 23268 48748 24668 48804
rect 24724 48748 24734 48804
rect 26114 48748 26124 48804
rect 26180 48748 26348 48804
rect 26404 48748 26414 48804
rect 35522 48748 35532 48804
rect 35588 48748 35756 48804
rect 35812 48748 35822 48804
rect 42130 48748 42140 48804
rect 42196 48748 43372 48804
rect 43428 48748 43438 48804
rect 43698 48748 43708 48804
rect 43764 48748 44716 48804
rect 44772 48748 45500 48804
rect 45556 48748 45566 48804
rect 3164 48692 3220 48748
rect 5068 48692 5124 48748
rect 22540 48692 22596 48748
rect 3164 48636 3388 48692
rect 3444 48636 3454 48692
rect 5058 48636 5068 48692
rect 5124 48636 5134 48692
rect 5852 48636 6916 48692
rect 11666 48636 11676 48692
rect 11732 48636 17220 48692
rect 17378 48636 17388 48692
rect 17444 48636 19292 48692
rect 19348 48636 19358 48692
rect 19506 48636 19516 48692
rect 19572 48636 19610 48692
rect 20178 48636 20188 48692
rect 20244 48636 23548 48692
rect 23604 48636 23614 48692
rect 24770 48636 24780 48692
rect 24836 48636 26908 48692
rect 32274 48636 32284 48692
rect 32340 48636 32844 48692
rect 32900 48636 33852 48692
rect 33908 48636 33918 48692
rect 37874 48636 37884 48692
rect 37940 48636 40012 48692
rect 40068 48636 40078 48692
rect 5852 48580 5908 48636
rect 6860 48580 6916 48636
rect 17164 48580 17220 48636
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 26852 48580 26908 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 3332 48524 5908 48580
rect 6850 48524 6860 48580
rect 6916 48524 15148 48580
rect 15204 48524 15280 48580
rect 17164 48524 18284 48580
rect 18340 48524 18350 48580
rect 18498 48524 18508 48580
rect 18564 48524 19628 48580
rect 19684 48524 19694 48580
rect 20514 48524 20524 48580
rect 20580 48524 20972 48580
rect 21028 48524 21038 48580
rect 26852 48524 33964 48580
rect 34020 48524 34860 48580
rect 34916 48524 34926 48580
rect 36866 48524 36876 48580
rect 36932 48524 36942 48580
rect 3332 48468 3388 48524
rect 1474 48412 1484 48468
rect 1540 48412 3388 48468
rect 4274 48412 4284 48468
rect 4340 48412 4844 48468
rect 4900 48412 4910 48468
rect 5404 48412 6636 48468
rect 6692 48412 6702 48468
rect 8082 48412 8092 48468
rect 8148 48412 12348 48468
rect 12404 48412 12414 48468
rect 12786 48412 12796 48468
rect 12852 48412 13804 48468
rect 13860 48412 13870 48468
rect 15250 48412 15260 48468
rect 15316 48412 21644 48468
rect 21700 48412 22092 48468
rect 22148 48412 22988 48468
rect 23044 48412 23100 48468
rect 23156 48412 23166 48468
rect 26002 48412 26012 48468
rect 26068 48412 29932 48468
rect 29988 48412 29998 48468
rect 30930 48412 30940 48468
rect 30996 48412 35868 48468
rect 35924 48412 36428 48468
rect 36484 48412 36494 48468
rect 5404 48356 5460 48412
rect 1586 48300 1596 48356
rect 1652 48300 5404 48356
rect 5460 48300 5470 48356
rect 6402 48300 6412 48356
rect 6468 48300 6972 48356
rect 7028 48300 7420 48356
rect 7476 48300 7486 48356
rect 9762 48300 9772 48356
rect 9828 48300 9884 48356
rect 9940 48300 9996 48356
rect 10052 48300 10062 48356
rect 10322 48300 10332 48356
rect 10388 48300 11228 48356
rect 11284 48300 12908 48356
rect 12964 48300 12974 48356
rect 13234 48300 13244 48356
rect 13300 48300 16492 48356
rect 16548 48300 16604 48356
rect 16660 48300 16670 48356
rect 16818 48300 16828 48356
rect 16884 48300 16922 48356
rect 17826 48300 17836 48356
rect 17892 48300 18172 48356
rect 18228 48300 19068 48356
rect 19124 48300 19134 48356
rect 19954 48300 19964 48356
rect 20020 48300 20860 48356
rect 20916 48300 20926 48356
rect 21746 48300 21756 48356
rect 21812 48300 23436 48356
rect 23492 48300 23660 48356
rect 23716 48300 23726 48356
rect 31826 48300 31836 48356
rect 31892 48300 32284 48356
rect 32340 48300 32350 48356
rect 4274 48188 4284 48244
rect 4340 48188 5068 48244
rect 5124 48188 5134 48244
rect 6514 48188 6524 48244
rect 6580 48188 6636 48244
rect 6692 48188 6860 48244
rect 6916 48188 6926 48244
rect 8642 48188 8652 48244
rect 8708 48188 11116 48244
rect 11172 48188 11182 48244
rect 11442 48188 11452 48244
rect 11508 48188 11676 48244
rect 11732 48188 11742 48244
rect 12450 48188 12460 48244
rect 12516 48188 12572 48244
rect 12628 48188 12638 48244
rect 17266 48188 17276 48244
rect 17332 48188 17724 48244
rect 17780 48188 17790 48244
rect 18386 48188 18396 48244
rect 18452 48188 23212 48244
rect 23268 48188 23278 48244
rect 26338 48188 26348 48244
rect 26404 48188 27132 48244
rect 27188 48188 27198 48244
rect 29922 48188 29932 48244
rect 29988 48188 31164 48244
rect 31220 48188 31230 48244
rect 32610 48188 32620 48244
rect 32676 48188 33628 48244
rect 33684 48188 33694 48244
rect 6524 48132 6580 48188
rect 11452 48132 11508 48188
rect 36876 48132 36932 48524
rect 38098 48412 38108 48468
rect 38164 48412 38892 48468
rect 38948 48412 38958 48468
rect 38546 48300 38556 48356
rect 38612 48300 39788 48356
rect 39844 48300 39854 48356
rect 43026 48300 43036 48356
rect 43092 48300 43932 48356
rect 43988 48300 44268 48356
rect 44324 48300 44334 48356
rect 44482 48300 44492 48356
rect 44548 48300 45388 48356
rect 45444 48300 45454 48356
rect 2146 48076 2156 48132
rect 2212 48076 6580 48132
rect 8530 48076 8540 48132
rect 8596 48076 8764 48132
rect 8820 48076 8830 48132
rect 10994 48076 11004 48132
rect 11060 48076 11508 48132
rect 11778 48076 11788 48132
rect 11844 48076 12124 48132
rect 12180 48076 17836 48132
rect 17892 48076 17902 48132
rect 18610 48076 18620 48132
rect 18676 48076 18732 48132
rect 18788 48076 18798 48132
rect 19282 48076 19292 48132
rect 19348 48076 20076 48132
rect 20132 48076 21644 48132
rect 21700 48076 21710 48132
rect 24882 48076 24892 48132
rect 24948 48076 26684 48132
rect 26740 48076 26908 48132
rect 26964 48076 26974 48132
rect 35298 48076 35308 48132
rect 35364 48076 35644 48132
rect 35700 48076 35710 48132
rect 36876 48076 36988 48132
rect 37044 48076 37548 48132
rect 37604 48076 37614 48132
rect 40338 48076 40348 48132
rect 40404 48076 41692 48132
rect 41748 48076 41758 48132
rect 43698 48076 43708 48132
rect 43764 48076 45276 48132
rect 45332 48076 45342 48132
rect 3910 47964 3948 48020
rect 4004 47964 4014 48020
rect 4172 47964 4900 48020
rect 5394 47964 5404 48020
rect 5460 47964 11452 48020
rect 11508 47964 11518 48020
rect 14130 47964 14140 48020
rect 14196 47964 18732 48020
rect 18788 47964 18798 48020
rect 19842 47964 19852 48020
rect 19908 47964 20524 48020
rect 20580 47964 20590 48020
rect 25218 47964 25228 48020
rect 25284 47964 26012 48020
rect 26068 47964 26078 48020
rect 26562 47964 26572 48020
rect 26628 47964 27916 48020
rect 27972 47964 28644 48020
rect 30930 47964 30940 48020
rect 30996 47964 39228 48020
rect 39284 47964 39294 48020
rect 4172 47908 4228 47964
rect 2818 47852 2828 47908
rect 2884 47852 2894 47908
rect 3490 47852 3500 47908
rect 3556 47852 4228 47908
rect 2828 47684 2884 47852
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 4844 47796 4900 47964
rect 28588 47908 28644 47964
rect 7970 47852 7980 47908
rect 8036 47852 21308 47908
rect 21364 47852 21374 47908
rect 23538 47852 23548 47908
rect 23604 47852 24108 47908
rect 24164 47852 24174 47908
rect 28578 47852 28588 47908
rect 28644 47852 28654 47908
rect 36726 47852 36764 47908
rect 36820 47852 36830 47908
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 4844 47740 10108 47796
rect 10164 47740 13020 47796
rect 13076 47740 13086 47796
rect 13346 47740 13356 47796
rect 13412 47740 15148 47796
rect 15204 47740 15260 47796
rect 15316 47740 15326 47796
rect 18946 47740 18956 47796
rect 19012 47740 20860 47796
rect 20916 47740 21196 47796
rect 21252 47740 21262 47796
rect 23650 47740 23660 47796
rect 23716 47740 23996 47796
rect 24052 47740 24062 47796
rect 28466 47740 28476 47796
rect 28532 47740 34300 47796
rect 34356 47740 34366 47796
rect 41010 47740 41020 47796
rect 41076 47740 41804 47796
rect 41860 47740 41870 47796
rect 2828 47628 3052 47684
rect 3108 47628 3276 47684
rect 3332 47628 6860 47684
rect 6916 47628 6926 47684
rect 8866 47628 8876 47684
rect 8932 47628 9212 47684
rect 9268 47628 9884 47684
rect 9940 47628 9950 47684
rect 13122 47628 13132 47684
rect 13188 47628 14028 47684
rect 14084 47628 14094 47684
rect 14466 47628 14476 47684
rect 14532 47628 15036 47684
rect 15092 47628 15102 47684
rect 17154 47628 17164 47684
rect 17220 47628 18172 47684
rect 18228 47628 18238 47684
rect 19282 47628 19292 47684
rect 19348 47628 19852 47684
rect 19908 47628 19918 47684
rect 20178 47628 20188 47684
rect 20244 47628 20524 47684
rect 20580 47628 20590 47684
rect 21074 47628 21084 47684
rect 21140 47628 22540 47684
rect 22596 47628 22606 47684
rect 23314 47628 23324 47684
rect 23380 47628 30156 47684
rect 30212 47628 30222 47684
rect 34290 47628 34300 47684
rect 34356 47628 34860 47684
rect 34916 47628 34926 47684
rect 2146 47516 2156 47572
rect 2212 47516 4060 47572
rect 4116 47516 4508 47572
rect 4564 47516 4574 47572
rect 7308 47516 9996 47572
rect 10052 47516 10556 47572
rect 10612 47516 10622 47572
rect 10882 47516 10892 47572
rect 10948 47516 10958 47572
rect 12002 47516 12012 47572
rect 12068 47516 17444 47572
rect 17602 47516 17612 47572
rect 17668 47516 25452 47572
rect 25508 47516 26572 47572
rect 26628 47516 26638 47572
rect 29810 47516 29820 47572
rect 29876 47516 30268 47572
rect 30324 47516 30334 47572
rect 31938 47516 31948 47572
rect 32004 47516 32396 47572
rect 32452 47516 33068 47572
rect 33124 47516 33134 47572
rect 36530 47516 36540 47572
rect 36596 47516 37884 47572
rect 37940 47516 39004 47572
rect 39060 47516 39070 47572
rect 2034 47404 2044 47460
rect 2100 47404 3164 47460
rect 3220 47404 3230 47460
rect 4162 47404 4172 47460
rect 4228 47404 4732 47460
rect 4788 47404 4798 47460
rect 6402 47404 6412 47460
rect 6468 47404 6860 47460
rect 6916 47404 6926 47460
rect 7308 47348 7364 47516
rect 10892 47460 10948 47516
rect 17388 47460 17444 47516
rect 7970 47404 7980 47460
rect 8036 47404 8428 47460
rect 8484 47404 9436 47460
rect 9492 47404 9884 47460
rect 9940 47404 10948 47460
rect 14466 47404 14476 47460
rect 14532 47404 17164 47460
rect 17220 47404 17230 47460
rect 17388 47404 17500 47460
rect 17556 47404 17566 47460
rect 18274 47404 18284 47460
rect 18340 47404 19628 47460
rect 19684 47404 19694 47460
rect 23426 47404 23436 47460
rect 23492 47404 24444 47460
rect 24500 47404 24510 47460
rect 24882 47404 24892 47460
rect 24948 47404 25004 47460
rect 25060 47404 25070 47460
rect 27234 47404 27244 47460
rect 27300 47404 28140 47460
rect 28196 47404 28206 47460
rect 32806 47404 32844 47460
rect 32900 47404 32910 47460
rect 33842 47404 33852 47460
rect 33908 47404 35196 47460
rect 35252 47404 35262 47460
rect 35522 47404 35532 47460
rect 35588 47404 36652 47460
rect 36708 47404 37212 47460
rect 37268 47404 38108 47460
rect 38164 47404 38174 47460
rect 44594 47404 44604 47460
rect 44660 47404 46060 47460
rect 46116 47404 46126 47460
rect 17500 47348 17556 47404
rect 5618 47292 5628 47348
rect 5684 47292 7308 47348
rect 7364 47292 7374 47348
rect 8082 47292 8092 47348
rect 8148 47292 8988 47348
rect 9044 47292 9054 47348
rect 9202 47292 9212 47348
rect 9268 47292 9306 47348
rect 9650 47292 9660 47348
rect 9716 47292 10332 47348
rect 10388 47292 12236 47348
rect 12292 47292 12302 47348
rect 17500 47292 19964 47348
rect 20020 47292 22988 47348
rect 23044 47292 23054 47348
rect 23762 47292 23772 47348
rect 23828 47292 26012 47348
rect 26068 47292 26078 47348
rect 33170 47292 33180 47348
rect 33236 47292 33628 47348
rect 33684 47292 34076 47348
rect 34132 47292 34142 47348
rect 34290 47292 34300 47348
rect 34356 47292 38108 47348
rect 38164 47292 39676 47348
rect 39732 47292 40572 47348
rect 40628 47292 40638 47348
rect 43334 47292 43372 47348
rect 43428 47292 43438 47348
rect 1138 47180 1148 47236
rect 1204 47180 1484 47236
rect 1540 47180 3052 47236
rect 3108 47180 11340 47236
rect 11396 47180 11406 47236
rect 12786 47180 12796 47236
rect 12852 47180 14812 47236
rect 14868 47180 14878 47236
rect 15138 47180 15148 47236
rect 15204 47180 16044 47236
rect 16100 47180 16110 47236
rect 16594 47180 16604 47236
rect 16660 47180 17500 47236
rect 17556 47180 17566 47236
rect 19730 47180 19740 47236
rect 19796 47180 26124 47236
rect 26180 47180 29484 47236
rect 29540 47180 30156 47236
rect 30212 47180 31500 47236
rect 31556 47180 31566 47236
rect 35410 47180 35420 47236
rect 35476 47180 35980 47236
rect 36036 47180 36046 47236
rect 44146 47180 44156 47236
rect 44212 47180 44940 47236
rect 44996 47180 45724 47236
rect 45780 47180 45790 47236
rect 1698 47068 1708 47124
rect 1764 47068 5628 47124
rect 5684 47068 5694 47124
rect 5842 47068 5852 47124
rect 5908 47068 6636 47124
rect 6692 47068 6702 47124
rect 8082 47068 8092 47124
rect 8148 47068 9212 47124
rect 9268 47068 9278 47124
rect 9538 47068 9548 47124
rect 9604 47068 12572 47124
rect 12628 47068 12638 47124
rect 15250 47068 15260 47124
rect 15316 47068 15708 47124
rect 15764 47068 15774 47124
rect 24882 47068 24892 47124
rect 24948 47068 25004 47124
rect 25060 47068 25070 47124
rect 27570 47068 27580 47124
rect 27636 47068 27646 47124
rect 32834 47068 32844 47124
rect 32900 47068 32938 47124
rect 33058 47068 33068 47124
rect 33124 47068 33162 47124
rect 33618 47068 33628 47124
rect 33684 47068 34300 47124
rect 34356 47068 34366 47124
rect 36642 47068 36652 47124
rect 36708 47068 36988 47124
rect 37044 47068 37054 47124
rect 37874 47068 37884 47124
rect 37940 47068 38220 47124
rect 38276 47068 38556 47124
rect 38612 47068 38622 47124
rect 39218 47068 39228 47124
rect 39284 47068 40124 47124
rect 40180 47068 40190 47124
rect 41906 47068 41916 47124
rect 41972 47068 44492 47124
rect 44548 47068 44558 47124
rect 2492 47012 2548 47068
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 27580 47012 27636 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 2482 46956 2492 47012
rect 2548 46956 2558 47012
rect 4834 46956 4844 47012
rect 4900 46956 5404 47012
rect 5460 46956 10164 47012
rect 10658 46956 10668 47012
rect 10724 46956 16436 47012
rect 21746 46956 21756 47012
rect 21812 46956 21868 47012
rect 21924 46956 22764 47012
rect 22820 46956 22830 47012
rect 25106 46956 25116 47012
rect 25172 46956 28140 47012
rect 28196 46956 28206 47012
rect 32498 46956 32508 47012
rect 32564 46956 33180 47012
rect 33236 46956 35084 47012
rect 35140 46956 35150 47012
rect 37426 46956 37436 47012
rect 37492 46956 37772 47012
rect 37828 46956 38332 47012
rect 38388 46956 38398 47012
rect 2258 46844 2268 46900
rect 2324 46844 2334 46900
rect 2594 46844 2604 46900
rect 2660 46844 2828 46900
rect 2884 46844 3612 46900
rect 3668 46844 3678 46900
rect 4946 46844 4956 46900
rect 5012 46844 8092 46900
rect 8148 46844 8158 46900
rect 8866 46844 8876 46900
rect 8932 46844 9660 46900
rect 9716 46844 9726 46900
rect 2268 46788 2324 46844
rect 10108 46788 10164 46956
rect 16380 46900 16436 46956
rect 13458 46844 13468 46900
rect 13524 46844 14028 46900
rect 14084 46844 14094 46900
rect 16370 46844 16380 46900
rect 16436 46844 17052 46900
rect 17108 46844 17388 46900
rect 17444 46844 17454 46900
rect 17602 46844 17612 46900
rect 17668 46844 18060 46900
rect 18116 46844 18126 46900
rect 19058 46844 19068 46900
rect 19124 46844 19964 46900
rect 20020 46844 20188 46900
rect 20244 46844 20254 46900
rect 21298 46844 21308 46900
rect 21364 46844 22540 46900
rect 22596 46844 23212 46900
rect 23268 46844 25452 46900
rect 25508 46844 25518 46900
rect 31378 46844 31388 46900
rect 31444 46844 34412 46900
rect 34468 46844 34478 46900
rect 34626 46844 34636 46900
rect 34692 46844 38668 46900
rect 38724 46844 38734 46900
rect 2268 46732 3052 46788
rect 3108 46732 3118 46788
rect 4246 46732 4284 46788
rect 4340 46732 4350 46788
rect 5618 46732 5628 46788
rect 5684 46732 6524 46788
rect 6580 46732 6590 46788
rect 10108 46732 12460 46788
rect 12516 46732 14140 46788
rect 14196 46732 14206 46788
rect 15092 46732 15708 46788
rect 15764 46732 15774 46788
rect 15922 46732 15932 46788
rect 15988 46732 16828 46788
rect 16884 46732 16894 46788
rect 19618 46732 19628 46788
rect 19684 46732 26908 46788
rect 27346 46732 27356 46788
rect 27412 46732 28028 46788
rect 28084 46732 28094 46788
rect 35746 46732 35756 46788
rect 35812 46732 36876 46788
rect 36932 46732 36942 46788
rect 13468 46676 13524 46732
rect 2930 46620 2940 46676
rect 2996 46620 3724 46676
rect 3780 46620 3836 46676
rect 3892 46620 5740 46676
rect 5796 46620 6412 46676
rect 6468 46620 6478 46676
rect 11218 46620 11228 46676
rect 11284 46620 12124 46676
rect 12180 46620 13244 46676
rect 13300 46620 13310 46676
rect 13458 46620 13468 46676
rect 13524 46620 13534 46676
rect 14018 46620 14028 46676
rect 14084 46620 14094 46676
rect 14028 46564 14084 46620
rect 15092 46564 15148 46732
rect 26852 46676 26908 46732
rect 15586 46620 15596 46676
rect 15652 46620 16940 46676
rect 16996 46620 17006 46676
rect 18358 46620 18396 46676
rect 18452 46620 18462 46676
rect 18946 46620 18956 46676
rect 19012 46620 19628 46676
rect 19684 46620 19694 46676
rect 20626 46620 20636 46676
rect 20692 46620 24332 46676
rect 24388 46620 24398 46676
rect 26852 46620 31276 46676
rect 31332 46620 38780 46676
rect 38836 46620 38846 46676
rect 5058 46508 5068 46564
rect 5124 46508 7420 46564
rect 7476 46508 7486 46564
rect 11526 46508 11564 46564
rect 11620 46508 11630 46564
rect 14028 46508 14924 46564
rect 14980 46508 15148 46564
rect 15362 46508 15372 46564
rect 15428 46508 15820 46564
rect 15876 46508 18284 46564
rect 18340 46508 18350 46564
rect 19730 46508 19740 46564
rect 19796 46508 20972 46564
rect 21028 46508 21038 46564
rect 32022 46508 32060 46564
rect 32116 46508 32126 46564
rect 32722 46508 32732 46564
rect 32788 46508 35308 46564
rect 35364 46508 35374 46564
rect 59200 46452 59800 46480
rect 3462 46396 3500 46452
rect 3556 46396 3566 46452
rect 4162 46396 4172 46452
rect 4228 46396 6468 46452
rect 6598 46396 6636 46452
rect 6692 46396 6702 46452
rect 6962 46396 6972 46452
rect 7028 46396 8092 46452
rect 8148 46396 8652 46452
rect 8708 46396 8718 46452
rect 13682 46396 13692 46452
rect 13748 46396 14476 46452
rect 14532 46396 14542 46452
rect 14690 46396 14700 46452
rect 14756 46396 16156 46452
rect 16212 46396 16222 46452
rect 16818 46396 16828 46452
rect 16884 46396 18620 46452
rect 18676 46396 18686 46452
rect 19506 46396 19516 46452
rect 19572 46396 20076 46452
rect 20132 46396 24780 46452
rect 24836 46396 24846 46452
rect 27010 46396 27020 46452
rect 27076 46396 28364 46452
rect 28420 46396 28430 46452
rect 31714 46396 31724 46452
rect 31780 46396 35588 46452
rect 38070 46396 38108 46452
rect 38164 46396 38174 46452
rect 38612 46396 42364 46452
rect 42420 46396 42430 46452
rect 55346 46396 55356 46452
rect 55412 46396 59800 46452
rect 6412 46340 6468 46396
rect 35532 46340 35588 46396
rect 38612 46340 38668 46396
rect 59200 46368 59800 46396
rect 3714 46284 3724 46340
rect 3780 46284 3836 46340
rect 3892 46284 3902 46340
rect 5954 46284 5964 46340
rect 6020 46284 6030 46340
rect 6412 46284 9436 46340
rect 9492 46284 9996 46340
rect 10052 46284 10062 46340
rect 10322 46284 10332 46340
rect 10388 46284 10892 46340
rect 10948 46284 10958 46340
rect 13794 46284 13804 46340
rect 13860 46284 15484 46340
rect 15540 46284 15550 46340
rect 15820 46284 16604 46340
rect 16660 46284 16670 46340
rect 16930 46284 16940 46340
rect 16996 46284 17500 46340
rect 17556 46284 17566 46340
rect 24658 46284 24668 46340
rect 24724 46284 27244 46340
rect 27300 46284 27310 46340
rect 35532 46284 38668 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 5964 46228 6020 46284
rect 15820 46228 15876 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 2594 46172 2604 46228
rect 2660 46172 3948 46228
rect 4004 46172 4014 46228
rect 5964 46172 6412 46228
rect 6468 46172 6478 46228
rect 6738 46172 6748 46228
rect 6804 46172 6860 46228
rect 6916 46172 15820 46228
rect 15876 46172 15886 46228
rect 16034 46172 16044 46228
rect 16100 46172 29484 46228
rect 29540 46172 29550 46228
rect 3714 46060 3724 46116
rect 3780 46060 3836 46116
rect 3892 46060 3902 46116
rect 4610 46060 4620 46116
rect 4676 46060 5292 46116
rect 5348 46060 6188 46116
rect 6244 46060 6254 46116
rect 8530 46060 8540 46116
rect 8596 46060 11340 46116
rect 11396 46060 11406 46116
rect 13458 46060 13468 46116
rect 13524 46060 15596 46116
rect 15652 46060 15662 46116
rect 17938 46060 17948 46116
rect 18004 46060 19180 46116
rect 19236 46060 20300 46116
rect 20356 46060 20366 46116
rect 1922 45948 1932 46004
rect 1988 45948 4060 46004
rect 4116 45948 4126 46004
rect 4274 45948 4284 46004
rect 4340 45948 4508 46004
rect 4564 45948 7980 46004
rect 8036 45948 8046 46004
rect 10098 45948 10108 46004
rect 10164 45948 12684 46004
rect 12740 45948 12796 46004
rect 12852 45948 13580 46004
rect 13636 45948 13646 46004
rect 14018 45948 14028 46004
rect 14084 45948 25116 46004
rect 25172 45948 25676 46004
rect 25732 45948 25742 46004
rect 32946 45948 32956 46004
rect 33012 45948 33404 46004
rect 33460 45948 33470 46004
rect 33730 45948 33740 46004
rect 33796 45948 34860 46004
rect 34916 45948 34926 46004
rect 39666 45948 39676 46004
rect 39732 45948 40348 46004
rect 40404 45948 40414 46004
rect 3378 45836 3388 45892
rect 3444 45836 3520 45892
rect 3602 45836 3612 45892
rect 3668 45836 4396 45892
rect 4452 45836 4462 45892
rect 4620 45836 8428 45892
rect 8484 45836 8494 45892
rect 8642 45836 8652 45892
rect 8708 45836 8988 45892
rect 9044 45836 9054 45892
rect 11228 45836 15372 45892
rect 15428 45836 15438 45892
rect 16118 45836 16156 45892
rect 16212 45836 16222 45892
rect 16930 45836 16940 45892
rect 16996 45836 17052 45892
rect 17108 45836 18396 45892
rect 18452 45836 18462 45892
rect 20076 45836 23100 45892
rect 23156 45836 23166 45892
rect 23426 45836 23436 45892
rect 23492 45836 23884 45892
rect 23940 45836 23950 45892
rect 31602 45836 31612 45892
rect 31668 45836 31724 45892
rect 31780 45836 31790 45892
rect 36418 45836 36428 45892
rect 36484 45836 36988 45892
rect 37044 45836 37054 45892
rect 56690 45836 56700 45892
rect 56756 45836 57372 45892
rect 57428 45836 57438 45892
rect 3388 45556 3444 45836
rect 4620 45780 4676 45836
rect 11228 45780 11284 45836
rect 20076 45780 20132 45836
rect 3938 45724 3948 45780
rect 4004 45724 4060 45780
rect 4116 45724 4676 45780
rect 5394 45724 5404 45780
rect 5460 45724 10108 45780
rect 10164 45724 10174 45780
rect 10434 45724 10444 45780
rect 10500 45724 10780 45780
rect 10836 45724 11228 45780
rect 11284 45724 11294 45780
rect 12450 45724 12460 45780
rect 12516 45724 13804 45780
rect 13860 45724 13870 45780
rect 15026 45724 15036 45780
rect 15092 45724 15372 45780
rect 15428 45724 15438 45780
rect 15810 45724 15820 45780
rect 15876 45724 20132 45780
rect 20486 45724 20524 45780
rect 20580 45724 20590 45780
rect 35298 45724 35308 45780
rect 35364 45724 41132 45780
rect 41188 45724 41198 45780
rect 44370 45724 44380 45780
rect 44436 45724 45500 45780
rect 45556 45724 45566 45780
rect 56130 45724 56140 45780
rect 56196 45724 57148 45780
rect 57204 45724 57214 45780
rect 20524 45668 20580 45724
rect 4050 45612 4060 45668
rect 4116 45612 4452 45668
rect 5506 45612 5516 45668
rect 5572 45612 6972 45668
rect 7028 45612 7308 45668
rect 7364 45612 7374 45668
rect 7858 45612 7868 45668
rect 7924 45612 8652 45668
rect 8708 45612 8718 45668
rect 10098 45612 10108 45668
rect 10164 45612 17948 45668
rect 18004 45612 18014 45668
rect 19506 45612 19516 45668
rect 19572 45612 20580 45668
rect 25442 45612 25452 45668
rect 25508 45612 26236 45668
rect 26292 45612 26302 45668
rect 27010 45612 27020 45668
rect 27076 45612 31052 45668
rect 31108 45612 31388 45668
rect 31444 45612 31454 45668
rect 33842 45612 33852 45668
rect 33908 45612 36372 45668
rect 36530 45612 36540 45668
rect 36596 45612 37548 45668
rect 37604 45612 37614 45668
rect 4396 45556 4452 45612
rect 3388 45500 3948 45556
rect 4004 45500 4172 45556
rect 4228 45500 4238 45556
rect 4396 45500 6020 45556
rect 6738 45500 6748 45556
rect 6804 45500 7196 45556
rect 7252 45500 7262 45556
rect 7410 45500 7420 45556
rect 7476 45500 12796 45556
rect 12852 45500 14588 45556
rect 14644 45500 15372 45556
rect 15428 45500 15932 45556
rect 15988 45500 15998 45556
rect 18274 45500 18284 45556
rect 18340 45500 18844 45556
rect 18900 45500 18910 45556
rect 20178 45500 20188 45556
rect 20244 45500 20748 45556
rect 20804 45500 20814 45556
rect 28242 45500 28252 45556
rect 28308 45500 29484 45556
rect 29540 45500 30044 45556
rect 30100 45500 31164 45556
rect 31220 45500 31230 45556
rect 5964 45444 6020 45500
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 36316 45444 36372 45612
rect 39442 45500 39452 45556
rect 39508 45500 39788 45556
rect 39844 45500 39854 45556
rect 39452 45444 39508 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 2706 45388 2716 45444
rect 2772 45388 5740 45444
rect 5796 45388 5806 45444
rect 5964 45388 8540 45444
rect 8596 45388 8606 45444
rect 9202 45388 9212 45444
rect 9268 45388 9772 45444
rect 9828 45388 9838 45444
rect 10182 45388 10220 45444
rect 10276 45388 10286 45444
rect 12114 45388 12124 45444
rect 12180 45388 15148 45444
rect 15586 45388 15596 45444
rect 15652 45388 15708 45444
rect 15764 45388 16716 45444
rect 16772 45388 16782 45444
rect 22754 45388 22764 45444
rect 22820 45388 23660 45444
rect 23716 45388 24108 45444
rect 24164 45388 24174 45444
rect 33170 45388 33180 45444
rect 33236 45388 33404 45444
rect 33460 45388 33470 45444
rect 33842 45388 33852 45444
rect 33908 45388 34636 45444
rect 34692 45388 34702 45444
rect 36316 45388 36652 45444
rect 36708 45388 39508 45444
rect 15092 45332 15148 45388
rect 4498 45276 4508 45332
rect 4564 45276 6300 45332
rect 6356 45276 6366 45332
rect 7522 45276 7532 45332
rect 7588 45276 11788 45332
rect 13010 45276 13020 45332
rect 13076 45276 14252 45332
rect 14308 45276 14318 45332
rect 15092 45276 15596 45332
rect 15652 45276 15662 45332
rect 16034 45276 16044 45332
rect 16100 45276 21532 45332
rect 21588 45276 21598 45332
rect 26674 45276 26684 45332
rect 26740 45276 28140 45332
rect 28196 45276 28206 45332
rect 34514 45276 34524 45332
rect 34580 45276 35756 45332
rect 35812 45276 35822 45332
rect 38322 45276 38332 45332
rect 38388 45276 38892 45332
rect 38948 45276 41244 45332
rect 41300 45276 41310 45332
rect 11732 45220 11788 45276
rect 3602 45164 3612 45220
rect 3668 45164 6748 45220
rect 6804 45164 6814 45220
rect 6962 45164 6972 45220
rect 7028 45164 8204 45220
rect 8260 45164 8270 45220
rect 8530 45164 8540 45220
rect 8596 45164 9212 45220
rect 9268 45164 9278 45220
rect 9548 45164 9772 45220
rect 9828 45164 9838 45220
rect 11732 45164 13468 45220
rect 13524 45164 13534 45220
rect 14924 45164 15148 45220
rect 15204 45164 15214 45220
rect 15362 45164 15372 45220
rect 15428 45164 16716 45220
rect 16772 45164 16782 45220
rect 17490 45164 17500 45220
rect 17556 45164 18620 45220
rect 18676 45164 18686 45220
rect 19394 45164 19404 45220
rect 19460 45164 21868 45220
rect 21924 45164 21934 45220
rect 22418 45164 22428 45220
rect 22484 45164 22764 45220
rect 22820 45164 22830 45220
rect 24444 45164 26012 45220
rect 26068 45164 26078 45220
rect 27346 45164 27356 45220
rect 27412 45164 28028 45220
rect 28084 45164 28094 45220
rect 34524 45164 34860 45220
rect 34916 45164 34926 45220
rect 9548 45108 9604 45164
rect 2146 45052 2156 45108
rect 2212 45052 2828 45108
rect 2884 45052 2894 45108
rect 3266 45052 3276 45108
rect 3332 45052 3948 45108
rect 4004 45052 4014 45108
rect 6066 45052 6076 45108
rect 6132 45052 6860 45108
rect 6916 45052 6926 45108
rect 7494 45052 7532 45108
rect 7588 45052 7598 45108
rect 8614 45052 8652 45108
rect 8708 45052 8718 45108
rect 9202 45052 9212 45108
rect 9268 45052 9604 45108
rect 9772 45052 14364 45108
rect 14420 45052 14430 45108
rect 7532 44996 7588 45052
rect 9772 44996 9828 45052
rect 14924 44996 14980 45164
rect 24444 45108 24500 45164
rect 34524 45108 34580 45164
rect 39228 45108 39284 45276
rect 2034 44940 2044 44996
rect 2100 44940 3388 44996
rect 7532 44940 9828 44996
rect 11890 44940 11900 44996
rect 11956 44940 12012 44996
rect 12068 44940 12078 44996
rect 13356 44940 14980 44996
rect 15092 45052 16940 45108
rect 16996 45052 17006 45108
rect 18834 45052 18844 45108
rect 18900 45052 19740 45108
rect 19796 45052 19806 45108
rect 20626 45052 20636 45108
rect 20692 45052 24444 45108
rect 24500 45052 24510 45108
rect 26114 45052 26124 45108
rect 26180 45052 27132 45108
rect 27188 45052 28140 45108
rect 28196 45052 28206 45108
rect 33618 45052 33628 45108
rect 33684 45052 33964 45108
rect 34020 45052 34524 45108
rect 34580 45052 34590 45108
rect 34962 45052 34972 45108
rect 35028 45052 35532 45108
rect 35588 45052 35598 45108
rect 39218 45052 39228 45108
rect 39284 45052 39294 45108
rect 40002 45052 40012 45108
rect 40068 45052 40078 45108
rect 3332 44884 3388 44940
rect 3332 44828 4172 44884
rect 4228 44828 4844 44884
rect 4900 44828 11788 44884
rect 11844 44828 11854 44884
rect 12226 44828 12236 44884
rect 12292 44828 12796 44884
rect 12852 44828 12862 44884
rect 13356 44772 13412 44940
rect 15092 44884 15148 45052
rect 40012 44996 40068 45052
rect 15586 44940 15596 44996
rect 15652 44940 16716 44996
rect 16772 44940 16782 44996
rect 18050 44940 18060 44996
rect 18116 44940 19236 44996
rect 26898 44940 26908 44996
rect 26964 44940 38668 44996
rect 38994 44940 39004 44996
rect 39060 44940 40068 44996
rect 19180 44884 19236 44940
rect 5954 44716 5964 44772
rect 6020 44716 7532 44772
rect 7588 44716 7598 44772
rect 7746 44716 7756 44772
rect 7812 44716 8204 44772
rect 8260 44716 8270 44772
rect 11330 44716 11340 44772
rect 11396 44716 13412 44772
rect 13468 44828 15148 44884
rect 18498 44828 18508 44884
rect 18564 44828 18844 44884
rect 18900 44828 18910 44884
rect 19170 44828 19180 44884
rect 19236 44828 19628 44884
rect 19684 44828 20188 44884
rect 20244 44828 20254 44884
rect 20486 44828 20524 44884
rect 20580 44828 20590 44884
rect 24770 44828 24780 44884
rect 24836 44828 31276 44884
rect 31332 44828 31836 44884
rect 31892 44828 31902 44884
rect 36082 44828 36092 44884
rect 36148 44828 38332 44884
rect 38388 44828 38398 44884
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 13468 44660 13524 44828
rect 13682 44716 13692 44772
rect 13748 44716 18844 44772
rect 18900 44716 19068 44772
rect 19124 44716 19134 44772
rect 24546 44716 24556 44772
rect 24612 44716 29148 44772
rect 29204 44716 29214 44772
rect 31574 44716 31612 44772
rect 31668 44716 31678 44772
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 38612 44660 38668 44940
rect 6290 44604 6300 44660
rect 6356 44604 6860 44660
rect 6916 44604 8428 44660
rect 8484 44604 13524 44660
rect 14466 44604 14476 44660
rect 14532 44604 25340 44660
rect 25396 44604 25900 44660
rect 25956 44604 26460 44660
rect 26516 44604 27132 44660
rect 27188 44604 27692 44660
rect 27748 44604 27758 44660
rect 35634 44604 35644 44660
rect 35700 44604 35868 44660
rect 35924 44604 35934 44660
rect 38612 44604 42364 44660
rect 42420 44604 42430 44660
rect 1586 44492 1596 44548
rect 1652 44492 2492 44548
rect 2548 44492 2558 44548
rect 4498 44492 4508 44548
rect 4564 44492 8204 44548
rect 8260 44492 9324 44548
rect 9380 44492 9390 44548
rect 11890 44492 11900 44548
rect 11956 44492 12012 44548
rect 12068 44492 12078 44548
rect 12562 44492 12572 44548
rect 12628 44492 13468 44548
rect 13524 44492 13534 44548
rect 14018 44492 14028 44548
rect 14084 44492 15260 44548
rect 15316 44492 15326 44548
rect 18918 44492 18956 44548
rect 19012 44492 19022 44548
rect 20178 44492 20188 44548
rect 20244 44492 21308 44548
rect 21364 44492 21374 44548
rect 32946 44492 32956 44548
rect 33012 44492 33516 44548
rect 33572 44492 33582 44548
rect 38994 44492 39004 44548
rect 39060 44492 42700 44548
rect 42756 44492 42766 44548
rect 200 44436 800 44464
rect 200 44380 1932 44436
rect 1988 44380 1998 44436
rect 6822 44380 6860 44436
rect 6916 44380 7980 44436
rect 8036 44380 8046 44436
rect 14130 44380 14140 44436
rect 14196 44380 17500 44436
rect 17556 44380 17566 44436
rect 17714 44380 17724 44436
rect 17780 44380 19068 44436
rect 19124 44380 19134 44436
rect 25890 44380 25900 44436
rect 25956 44380 26684 44436
rect 26740 44380 26750 44436
rect 35634 44380 35644 44436
rect 35700 44380 36988 44436
rect 37044 44380 37054 44436
rect 38546 44380 38556 44436
rect 38612 44380 39452 44436
rect 39508 44380 39518 44436
rect 43474 44380 43484 44436
rect 43540 44380 44156 44436
rect 44212 44380 44222 44436
rect 200 44352 800 44380
rect 2930 44268 2940 44324
rect 2996 44268 3948 44324
rect 4004 44268 4014 44324
rect 6626 44268 6636 44324
rect 6692 44268 8428 44324
rect 8484 44268 8494 44324
rect 9314 44268 9324 44324
rect 9380 44268 9660 44324
rect 9716 44268 9726 44324
rect 11442 44268 11452 44324
rect 11508 44268 14252 44324
rect 14308 44268 14318 44324
rect 21858 44268 21868 44324
rect 21924 44268 23212 44324
rect 23268 44268 23278 44324
rect 23426 44268 23436 44324
rect 23492 44268 24108 44324
rect 24164 44268 24174 44324
rect 30482 44268 30492 44324
rect 30548 44268 36764 44324
rect 36820 44268 36830 44324
rect 37314 44268 37324 44324
rect 37380 44268 39676 44324
rect 39732 44268 39742 44324
rect 41794 44268 41804 44324
rect 41860 44268 43932 44324
rect 43988 44268 44268 44324
rect 44324 44268 44334 44324
rect 44706 44268 44716 44324
rect 44772 44268 45052 44324
rect 45108 44268 45500 44324
rect 45556 44268 45566 44324
rect 36764 44212 36820 44268
rect 3266 44156 3276 44212
rect 3332 44156 8988 44212
rect 9044 44156 9054 44212
rect 9398 44156 9436 44212
rect 9492 44156 9502 44212
rect 9734 44156 9772 44212
rect 9828 44156 11676 44212
rect 11732 44156 11742 44212
rect 13654 44156 13692 44212
rect 13748 44156 13758 44212
rect 15698 44156 15708 44212
rect 15764 44156 24220 44212
rect 24276 44156 24286 44212
rect 26450 44156 26460 44212
rect 26516 44156 26684 44212
rect 26740 44156 26750 44212
rect 32274 44156 32284 44212
rect 32340 44156 33292 44212
rect 33348 44156 33358 44212
rect 36764 44156 38556 44212
rect 38612 44156 38622 44212
rect 43138 44156 43148 44212
rect 43204 44156 44044 44212
rect 44100 44156 44110 44212
rect 5618 44044 5628 44100
rect 5684 44044 5964 44100
rect 6020 44044 7532 44100
rect 7588 44044 7598 44100
rect 9136 44044 9212 44100
rect 9268 44044 9884 44100
rect 9940 44044 9950 44100
rect 13458 44044 13468 44100
rect 13524 44044 14140 44100
rect 14196 44044 14206 44100
rect 15138 44044 15148 44100
rect 15204 44044 16604 44100
rect 16660 44044 17388 44100
rect 17444 44044 17724 44100
rect 17780 44044 17790 44100
rect 18274 44044 18284 44100
rect 18340 44044 22092 44100
rect 22148 44044 22158 44100
rect 23062 44044 23100 44100
rect 23156 44044 24556 44100
rect 24612 44044 24622 44100
rect 29362 44044 29372 44100
rect 29428 44044 29596 44100
rect 29652 44044 29708 44100
rect 29764 44044 30716 44100
rect 30772 44044 30782 44100
rect 32162 44044 32172 44100
rect 32228 44044 33516 44100
rect 33572 44044 33582 44100
rect 3154 43932 3164 43988
rect 3220 43932 6972 43988
rect 7028 43932 7644 43988
rect 7700 43932 7710 43988
rect 7858 43932 7868 43988
rect 7924 43932 11788 43988
rect 11844 43932 12460 43988
rect 12516 43932 12526 43988
rect 12674 43932 12684 43988
rect 12740 43932 16044 43988
rect 16100 43932 16110 43988
rect 16706 43932 16716 43988
rect 16772 43932 17164 43988
rect 17220 43932 17230 43988
rect 18806 43932 18844 43988
rect 18900 43932 18910 43988
rect 21298 43932 21308 43988
rect 21364 43932 23996 43988
rect 24052 43932 24062 43988
rect 27682 43932 27692 43988
rect 27748 43932 28252 43988
rect 28308 43932 28318 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 6626 43820 6636 43876
rect 6692 43820 6748 43876
rect 6804 43820 8092 43876
rect 8148 43820 8158 43876
rect 8978 43820 8988 43876
rect 9044 43820 9772 43876
rect 9828 43820 10332 43876
rect 10388 43820 10398 43876
rect 12310 43820 12348 43876
rect 12404 43820 12414 43876
rect 17490 43820 17500 43876
rect 17556 43820 18620 43876
rect 18676 43820 18686 43876
rect 20402 43820 20412 43876
rect 20468 43820 23324 43876
rect 23380 43820 23390 43876
rect 28690 43820 28700 43876
rect 28756 43820 29708 43876
rect 29764 43820 36652 43876
rect 36708 43820 36718 43876
rect 8092 43764 8148 43820
rect 2706 43708 2716 43764
rect 2772 43708 5292 43764
rect 5348 43708 5852 43764
rect 5908 43708 5918 43764
rect 8092 43708 12572 43764
rect 12628 43708 12638 43764
rect 13234 43708 13244 43764
rect 13300 43708 13692 43764
rect 13748 43708 15596 43764
rect 15652 43708 15662 43764
rect 16930 43708 16940 43764
rect 16996 43708 19740 43764
rect 19796 43708 21420 43764
rect 21476 43708 21980 43764
rect 22036 43708 22046 43764
rect 28914 43708 28924 43764
rect 28980 43708 29372 43764
rect 29428 43708 30156 43764
rect 30212 43708 30222 43764
rect 37202 43708 37212 43764
rect 37268 43708 37996 43764
rect 38052 43708 39228 43764
rect 39284 43708 40460 43764
rect 40516 43708 40526 43764
rect 42354 43708 42364 43764
rect 42420 43708 43372 43764
rect 43428 43708 43438 43764
rect 2818 43596 2828 43652
rect 2884 43596 6748 43652
rect 6804 43596 6814 43652
rect 8082 43596 8092 43652
rect 8148 43596 8540 43652
rect 8596 43596 9100 43652
rect 9156 43596 9166 43652
rect 12226 43596 12236 43652
rect 12292 43596 13580 43652
rect 13636 43596 13646 43652
rect 15138 43596 15148 43652
rect 15204 43596 15260 43652
rect 15316 43596 15326 43652
rect 15810 43596 15820 43652
rect 15876 43596 16716 43652
rect 16772 43596 16782 43652
rect 16940 43596 18508 43652
rect 18564 43596 18574 43652
rect 18806 43596 18844 43652
rect 18900 43596 18910 43652
rect 19394 43596 19404 43652
rect 19460 43596 20636 43652
rect 20692 43596 20702 43652
rect 22082 43596 22092 43652
rect 22148 43596 23548 43652
rect 23604 43596 23614 43652
rect 26674 43596 26684 43652
rect 26740 43596 27020 43652
rect 27076 43596 27244 43652
rect 27300 43596 27310 43652
rect 31714 43596 31724 43652
rect 31780 43596 32620 43652
rect 32676 43596 34412 43652
rect 34468 43596 34478 43652
rect 40114 43596 40124 43652
rect 40180 43596 40796 43652
rect 40852 43596 40862 43652
rect 42802 43596 42812 43652
rect 42868 43596 43708 43652
rect 43764 43596 43774 43652
rect 16940 43540 16996 43596
rect 2258 43484 2268 43540
rect 2324 43484 2940 43540
rect 2996 43484 4172 43540
rect 4228 43484 4238 43540
rect 5516 43484 5852 43540
rect 5908 43484 7420 43540
rect 7476 43484 7486 43540
rect 7858 43484 7868 43540
rect 7924 43484 10108 43540
rect 10164 43484 10174 43540
rect 10994 43484 11004 43540
rect 11060 43484 12348 43540
rect 12404 43484 13356 43540
rect 13412 43484 13422 43540
rect 14018 43484 14028 43540
rect 14084 43484 14812 43540
rect 14868 43484 15260 43540
rect 15316 43484 15326 43540
rect 16930 43484 16940 43540
rect 16996 43484 17006 43540
rect 17686 43484 17724 43540
rect 17780 43484 17790 43540
rect 18274 43484 18284 43540
rect 18340 43484 19964 43540
rect 20020 43484 20030 43540
rect 20290 43484 20300 43540
rect 20356 43484 21532 43540
rect 21588 43484 22316 43540
rect 22372 43484 22382 43540
rect 34626 43484 34636 43540
rect 34692 43484 34972 43540
rect 35028 43484 35038 43540
rect 37650 43484 37660 43540
rect 37716 43484 37884 43540
rect 37940 43484 38444 43540
rect 38500 43484 40572 43540
rect 40628 43484 40638 43540
rect 41794 43484 41804 43540
rect 41860 43484 42364 43540
rect 42420 43484 42430 43540
rect 43250 43484 43260 43540
rect 43316 43484 44156 43540
rect 44212 43484 44222 43540
rect 44370 43484 44380 43540
rect 44436 43484 44828 43540
rect 44884 43484 45948 43540
rect 46004 43484 46014 43540
rect 5516 43428 5572 43484
rect 1810 43372 1820 43428
rect 1876 43372 5516 43428
rect 5572 43372 5582 43428
rect 6066 43372 6076 43428
rect 6132 43372 7756 43428
rect 7812 43372 7822 43428
rect 8306 43372 8316 43428
rect 8372 43372 8988 43428
rect 9044 43372 9212 43428
rect 9268 43372 9660 43428
rect 9716 43372 9726 43428
rect 9986 43372 9996 43428
rect 10052 43372 10780 43428
rect 10836 43372 13692 43428
rect 13748 43372 13758 43428
rect 14130 43372 14140 43428
rect 14196 43372 21084 43428
rect 21140 43372 22540 43428
rect 22596 43372 22606 43428
rect 24994 43372 25004 43428
rect 25060 43372 25900 43428
rect 25956 43372 26348 43428
rect 26404 43372 26414 43428
rect 30594 43372 30604 43428
rect 30660 43372 31500 43428
rect 31556 43372 31836 43428
rect 31892 43372 32284 43428
rect 32340 43372 32350 43428
rect 32610 43372 32620 43428
rect 32676 43372 34188 43428
rect 34244 43372 34524 43428
rect 34580 43372 34590 43428
rect 39330 43372 39340 43428
rect 39396 43372 42700 43428
rect 42756 43372 42766 43428
rect 1922 43260 1932 43316
rect 1988 43260 3724 43316
rect 3780 43260 8428 43316
rect 8484 43260 8494 43316
rect 14354 43260 14364 43316
rect 14420 43260 14588 43316
rect 14644 43260 14654 43316
rect 15586 43260 15596 43316
rect 15652 43260 18844 43316
rect 18900 43260 20412 43316
rect 20468 43260 20478 43316
rect 21634 43260 21644 43316
rect 21700 43260 27020 43316
rect 27076 43260 27086 43316
rect 34850 43260 34860 43316
rect 34916 43260 35868 43316
rect 35924 43260 35934 43316
rect 36194 43260 36204 43316
rect 36260 43260 39900 43316
rect 39956 43260 39966 43316
rect 43138 43260 43148 43316
rect 43204 43260 44156 43316
rect 44212 43260 44222 43316
rect 39116 43204 39172 43260
rect 3490 43148 3500 43204
rect 3556 43148 3612 43204
rect 3668 43148 3678 43204
rect 4834 43148 4844 43204
rect 4900 43148 11900 43204
rect 11956 43148 11966 43204
rect 15698 43148 15708 43204
rect 15764 43148 19852 43204
rect 19908 43148 19918 43204
rect 21522 43148 21532 43204
rect 21588 43148 22428 43204
rect 22484 43148 22494 43204
rect 36082 43148 36092 43204
rect 36148 43148 36652 43204
rect 36708 43148 36718 43204
rect 39106 43148 39116 43204
rect 39172 43148 39182 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 3266 43036 3276 43092
rect 3332 43036 3388 43092
rect 3444 43036 3454 43092
rect 5282 43036 5292 43092
rect 5348 43036 6524 43092
rect 6580 43036 9548 43092
rect 9604 43036 9614 43092
rect 10882 43036 10892 43092
rect 10948 43036 18732 43092
rect 18788 43036 19404 43092
rect 19460 43036 20524 43092
rect 20580 43036 20590 43092
rect 1362 42924 1372 42980
rect 1428 42924 5404 42980
rect 5460 42924 6076 42980
rect 6132 42924 6142 42980
rect 6402 42924 6412 42980
rect 6468 42924 6524 42980
rect 6580 42924 6590 42980
rect 6738 42924 6748 42980
rect 6804 42924 11900 42980
rect 11956 42924 15260 42980
rect 15316 42924 15326 42980
rect 15474 42924 15484 42980
rect 15540 42924 17500 42980
rect 17556 42924 18060 42980
rect 18116 42924 18126 42980
rect 18386 42924 18396 42980
rect 18452 42924 18956 42980
rect 19012 42924 19628 42980
rect 19684 42924 19694 42980
rect 22642 42924 22652 42980
rect 22708 42924 29484 42980
rect 29540 42924 29932 42980
rect 29988 42924 30716 42980
rect 30772 42924 32060 42980
rect 32116 42924 33516 42980
rect 33572 42924 33582 42980
rect 35186 42924 35196 42980
rect 35252 42924 36316 42980
rect 36372 42924 36382 42980
rect 2594 42812 2604 42868
rect 2660 42812 3836 42868
rect 3892 42812 3902 42868
rect 6290 42812 6300 42868
rect 6356 42812 6412 42868
rect 6468 42812 10220 42868
rect 10276 42812 10286 42868
rect 14018 42812 14028 42868
rect 14084 42812 16268 42868
rect 16324 42812 16334 42868
rect 16930 42812 16940 42868
rect 16996 42812 19516 42868
rect 19572 42812 19582 42868
rect 19730 42812 19740 42868
rect 19796 42812 26012 42868
rect 26068 42812 26078 42868
rect 2258 42700 2268 42756
rect 2324 42700 3612 42756
rect 3668 42700 3678 42756
rect 6178 42700 6188 42756
rect 6244 42700 6748 42756
rect 6804 42700 6814 42756
rect 9874 42700 9884 42756
rect 9940 42700 11228 42756
rect 11284 42700 12124 42756
rect 12180 42700 12190 42756
rect 14354 42700 14364 42756
rect 14420 42700 19180 42756
rect 19236 42700 19246 42756
rect 22642 42700 22652 42756
rect 22708 42700 23100 42756
rect 23156 42700 23166 42756
rect 23650 42700 23660 42756
rect 23716 42700 25676 42756
rect 25732 42700 26796 42756
rect 26852 42700 26862 42756
rect 34626 42700 34636 42756
rect 34692 42700 34860 42756
rect 34916 42700 34926 42756
rect 38098 42700 38108 42756
rect 38164 42700 38892 42756
rect 38948 42700 39564 42756
rect 39620 42700 40124 42756
rect 40180 42700 40190 42756
rect 44258 42700 44268 42756
rect 44324 42700 46172 42756
rect 46228 42700 46238 42756
rect 6188 42644 6244 42700
rect 2146 42588 2156 42644
rect 2212 42588 2828 42644
rect 2884 42588 2894 42644
rect 3714 42588 3724 42644
rect 3780 42588 6244 42644
rect 6626 42588 6636 42644
rect 6692 42588 7308 42644
rect 7364 42588 10444 42644
rect 10500 42588 10510 42644
rect 11330 42588 11340 42644
rect 11396 42588 11452 42644
rect 11508 42588 11518 42644
rect 13458 42588 13468 42644
rect 13524 42588 13692 42644
rect 13748 42588 13758 42644
rect 13906 42588 13916 42644
rect 13972 42588 14812 42644
rect 14868 42588 14878 42644
rect 15782 42588 15820 42644
rect 15876 42588 15886 42644
rect 17938 42588 17948 42644
rect 18004 42588 18620 42644
rect 18676 42588 18686 42644
rect 20066 42588 20076 42644
rect 20132 42588 23548 42644
rect 23604 42588 23614 42644
rect 30146 42588 30156 42644
rect 30212 42588 30492 42644
rect 30548 42588 30558 42644
rect 34402 42588 34412 42644
rect 34468 42588 35756 42644
rect 35812 42588 35822 42644
rect 35970 42588 35980 42644
rect 36036 42588 36046 42644
rect 3378 42476 3388 42532
rect 3444 42476 8316 42532
rect 8372 42476 8382 42532
rect 8530 42476 8540 42532
rect 8596 42476 8634 42532
rect 13122 42476 13132 42532
rect 13188 42476 15932 42532
rect 15988 42476 15998 42532
rect 16146 42476 16156 42532
rect 16212 42476 16492 42532
rect 16548 42476 16558 42532
rect 17378 42476 17388 42532
rect 17444 42476 18396 42532
rect 18452 42476 18462 42532
rect 18946 42476 18956 42532
rect 19012 42476 22204 42532
rect 22260 42476 22270 42532
rect 22502 42476 22540 42532
rect 22596 42476 22606 42532
rect 23090 42476 23100 42532
rect 23156 42476 24444 42532
rect 24500 42476 24510 42532
rect 34822 42476 34860 42532
rect 34916 42476 34926 42532
rect 35980 42420 36036 42588
rect 38434 42476 38444 42532
rect 38500 42476 39004 42532
rect 39060 42476 39070 42532
rect 2146 42364 2156 42420
rect 2212 42364 10108 42420
rect 10164 42364 10780 42420
rect 10836 42364 10846 42420
rect 11554 42364 11564 42420
rect 11620 42364 12124 42420
rect 12180 42364 13692 42420
rect 13748 42364 13758 42420
rect 15110 42364 15148 42420
rect 15204 42364 15214 42420
rect 16034 42364 16044 42420
rect 16100 42364 19684 42420
rect 28018 42364 28028 42420
rect 28084 42364 29596 42420
rect 29652 42364 29662 42420
rect 32498 42364 32508 42420
rect 32564 42364 34972 42420
rect 35028 42364 36036 42420
rect 3798 42252 3836 42308
rect 3892 42252 3902 42308
rect 7746 42252 7756 42308
rect 7812 42252 13132 42308
rect 13188 42252 13198 42308
rect 13356 42252 14588 42308
rect 14644 42252 15372 42308
rect 15428 42252 16268 42308
rect 16324 42252 16334 42308
rect 18610 42252 18620 42308
rect 18676 42252 19292 42308
rect 19348 42252 19358 42308
rect 13356 42196 13412 42252
rect 19628 42196 19684 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 26786 42252 26796 42308
rect 26852 42252 26862 42308
rect 34178 42252 34188 42308
rect 34244 42252 37436 42308
rect 37492 42252 37772 42308
rect 37828 42252 37838 42308
rect 26796 42196 26852 42252
rect 2818 42140 2828 42196
rect 2884 42140 7420 42196
rect 7476 42140 8204 42196
rect 8260 42140 8270 42196
rect 9510 42140 9548 42196
rect 9604 42140 9614 42196
rect 10892 42140 13412 42196
rect 14130 42140 14140 42196
rect 14196 42140 16604 42196
rect 16660 42140 16670 42196
rect 19628 42140 21644 42196
rect 21700 42140 21710 42196
rect 22418 42140 22428 42196
rect 22484 42140 23324 42196
rect 23380 42140 23390 42196
rect 25218 42140 25228 42196
rect 25284 42140 25452 42196
rect 25508 42140 25518 42196
rect 26450 42140 26460 42196
rect 26516 42140 27580 42196
rect 27636 42140 27646 42196
rect 29474 42140 29484 42196
rect 29540 42140 35756 42196
rect 35812 42140 35822 42196
rect 37650 42140 37660 42196
rect 37716 42140 38892 42196
rect 38948 42140 38958 42196
rect 10892 42084 10948 42140
rect 3154 42028 3164 42084
rect 3220 42028 3388 42084
rect 3444 42028 3454 42084
rect 4806 42028 4844 42084
rect 4900 42028 4910 42084
rect 5478 42028 5516 42084
rect 5572 42028 5582 42084
rect 7410 42028 7420 42084
rect 7476 42028 7756 42084
rect 7812 42028 7822 42084
rect 8530 42028 8540 42084
rect 8596 42028 9324 42084
rect 9380 42028 10948 42084
rect 12674 42028 12684 42084
rect 12740 42028 17724 42084
rect 17780 42028 17790 42084
rect 18050 42028 18060 42084
rect 18116 42028 21420 42084
rect 21476 42028 21486 42084
rect 22642 42028 22652 42084
rect 22708 42028 23772 42084
rect 23828 42028 23838 42084
rect 24444 42028 25004 42084
rect 25060 42028 25228 42084
rect 25284 42028 25294 42084
rect 26002 42028 26012 42084
rect 26068 42028 26684 42084
rect 26740 42028 26750 42084
rect 26898 42028 26908 42084
rect 26964 42028 29820 42084
rect 29876 42028 29886 42084
rect 30594 42028 30604 42084
rect 30660 42028 31948 42084
rect 32004 42028 32014 42084
rect 32386 42028 32396 42084
rect 32452 42028 33964 42084
rect 34020 42028 34030 42084
rect 34290 42028 34300 42084
rect 34356 42028 35420 42084
rect 35476 42028 35486 42084
rect 35634 42028 35644 42084
rect 35700 42028 35868 42084
rect 35924 42028 36316 42084
rect 36372 42028 36540 42084
rect 36596 42028 36606 42084
rect 40674 42028 40684 42084
rect 40740 42028 43708 42084
rect 43764 42028 43932 42084
rect 43988 42028 43998 42084
rect 24444 41972 24500 42028
rect 4162 41916 4172 41972
rect 4228 41916 4620 41972
rect 4676 41916 6300 41972
rect 6356 41916 9772 41972
rect 9828 41916 10332 41972
rect 10388 41916 10398 41972
rect 10658 41916 10668 41972
rect 10724 41916 11788 41972
rect 11844 41916 11854 41972
rect 13010 41916 13020 41972
rect 13076 41916 13580 41972
rect 13636 41916 13646 41972
rect 15026 41916 15036 41972
rect 15092 41916 16044 41972
rect 16100 41916 16110 41972
rect 16482 41916 16492 41972
rect 16548 41916 16772 41972
rect 16930 41916 16940 41972
rect 16996 41916 17500 41972
rect 17556 41916 18844 41972
rect 18900 41916 18910 41972
rect 19058 41916 19068 41972
rect 19124 41916 24500 41972
rect 24658 41916 24668 41972
rect 24724 41916 25452 41972
rect 25508 41916 25676 41972
rect 25732 41916 25742 41972
rect 27010 41916 27020 41972
rect 27076 41916 27916 41972
rect 27972 41916 28588 41972
rect 28644 41916 28654 41972
rect 32834 41916 32844 41972
rect 32900 41916 33740 41972
rect 33796 41916 33806 41972
rect 38210 41916 38220 41972
rect 38276 41916 38668 41972
rect 38724 41916 39228 41972
rect 39284 41916 39294 41972
rect 40450 41916 40460 41972
rect 40516 41916 41468 41972
rect 41524 41916 41534 41972
rect 16716 41860 16772 41916
rect 2342 41804 2380 41860
rect 2436 41804 2446 41860
rect 4722 41804 4732 41860
rect 4788 41804 5292 41860
rect 5348 41804 5358 41860
rect 5506 41804 5516 41860
rect 5572 41804 5964 41860
rect 6020 41804 6188 41860
rect 6244 41804 7084 41860
rect 7140 41804 7150 41860
rect 8978 41804 8988 41860
rect 9044 41804 11452 41860
rect 11508 41804 11518 41860
rect 13570 41804 13580 41860
rect 13636 41804 14308 41860
rect 14252 41748 14308 41804
rect 15036 41804 15708 41860
rect 15764 41804 15774 41860
rect 16716 41804 20300 41860
rect 20356 41804 20366 41860
rect 21158 41804 21196 41860
rect 21252 41804 21262 41860
rect 23314 41804 23324 41860
rect 23380 41804 23660 41860
rect 23716 41804 23726 41860
rect 28242 41804 28252 41860
rect 28308 41804 36876 41860
rect 36932 41804 36942 41860
rect 1922 41692 1932 41748
rect 1988 41692 4900 41748
rect 5058 41692 5068 41748
rect 5124 41692 5740 41748
rect 5796 41692 5806 41748
rect 6738 41692 6748 41748
rect 6804 41692 10668 41748
rect 10724 41692 10734 41748
rect 13234 41692 13244 41748
rect 13300 41692 13916 41748
rect 13972 41692 13982 41748
rect 14242 41692 14252 41748
rect 14308 41692 14318 41748
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 4844 41524 4900 41692
rect 15036 41636 15092 41804
rect 16594 41692 16604 41748
rect 16660 41692 17612 41748
rect 17668 41692 17678 41748
rect 20738 41692 20748 41748
rect 20804 41692 23100 41748
rect 23156 41692 23166 41748
rect 39778 41692 39788 41748
rect 39844 41692 40572 41748
rect 40628 41692 40638 41748
rect 6514 41580 6524 41636
rect 6580 41580 15092 41636
rect 17276 41580 20524 41636
rect 20580 41580 22540 41636
rect 22596 41580 22606 41636
rect 23202 41580 23212 41636
rect 23268 41580 24556 41636
rect 24612 41580 24622 41636
rect 24994 41580 25004 41636
rect 25060 41580 28364 41636
rect 28420 41580 28430 41636
rect 4844 41468 6076 41524
rect 6132 41468 8428 41524
rect 8484 41468 8494 41524
rect 11442 41468 11452 41524
rect 11508 41468 14084 41524
rect 14028 41412 14084 41468
rect 6402 41356 6412 41412
rect 6468 41356 12124 41412
rect 12180 41356 12190 41412
rect 14018 41356 14028 41412
rect 14084 41356 14364 41412
rect 14420 41356 14430 41412
rect 17276 41300 17332 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 18946 41468 18956 41524
rect 19012 41468 19404 41524
rect 19460 41468 19852 41524
rect 19908 41468 19918 41524
rect 21074 41468 21084 41524
rect 21140 41468 21308 41524
rect 21364 41468 21868 41524
rect 21924 41468 21934 41524
rect 24098 41468 24108 41524
rect 24164 41468 31052 41524
rect 31108 41468 31836 41524
rect 31892 41468 32172 41524
rect 32228 41468 32844 41524
rect 32900 41468 32910 41524
rect 17602 41356 17612 41412
rect 17668 41356 18956 41412
rect 19012 41356 19022 41412
rect 19954 41356 19964 41412
rect 20020 41356 20748 41412
rect 20804 41356 22204 41412
rect 22260 41356 22876 41412
rect 22932 41356 22942 41412
rect 27010 41356 27020 41412
rect 27076 41356 27086 41412
rect 27020 41300 27076 41356
rect 3378 41244 3388 41300
rect 3444 41244 3724 41300
rect 3780 41244 4956 41300
rect 5012 41244 5964 41300
rect 6020 41244 6860 41300
rect 6916 41244 6926 41300
rect 7942 41244 7980 41300
rect 8036 41244 8046 41300
rect 13122 41244 13132 41300
rect 13188 41244 17332 41300
rect 20626 41244 20636 41300
rect 20692 41244 25228 41300
rect 25284 41244 25788 41300
rect 25844 41244 25854 41300
rect 26338 41244 26348 41300
rect 26404 41244 27076 41300
rect 27906 41244 27916 41300
rect 27972 41244 38668 41300
rect 38724 41244 39004 41300
rect 39060 41244 39340 41300
rect 39396 41244 39676 41300
rect 39732 41244 39742 41300
rect 3826 41132 3836 41188
rect 3892 41132 4620 41188
rect 4676 41132 4686 41188
rect 6598 41132 6636 41188
rect 6692 41132 6702 41188
rect 7298 41132 7308 41188
rect 7364 41132 7644 41188
rect 7700 41132 7710 41188
rect 9762 41132 9772 41188
rect 9828 41132 12012 41188
rect 12068 41132 12078 41188
rect 13570 41132 13580 41188
rect 13636 41132 14252 41188
rect 14308 41132 14318 41188
rect 17126 41132 17164 41188
rect 17220 41132 17230 41188
rect 19282 41132 19292 41188
rect 19348 41132 20412 41188
rect 20468 41132 20478 41188
rect 21186 41132 21196 41188
rect 21252 41132 23772 41188
rect 23828 41132 23838 41188
rect 28914 41132 28924 41188
rect 28980 41132 28990 41188
rect 42914 41132 42924 41188
rect 42980 41132 43820 41188
rect 43876 41132 45724 41188
rect 45780 41132 45790 41188
rect 28924 41076 28980 41132
rect 4050 41020 4060 41076
rect 4116 41020 4732 41076
rect 4788 41020 4798 41076
rect 4946 41020 4956 41076
rect 5012 41020 7532 41076
rect 7588 41020 7598 41076
rect 10658 41020 10668 41076
rect 10724 41020 14308 41076
rect 14914 41020 14924 41076
rect 14980 41020 15596 41076
rect 15652 41020 17724 41076
rect 17780 41020 17836 41076
rect 17892 41020 19516 41076
rect 19572 41020 21644 41076
rect 21700 41020 22540 41076
rect 22596 41020 22606 41076
rect 25190 41020 25228 41076
rect 25284 41020 25294 41076
rect 25778 41020 25788 41076
rect 25844 41020 28476 41076
rect 28532 41020 28542 41076
rect 28924 41020 40012 41076
rect 40068 41020 40348 41076
rect 40404 41020 40414 41076
rect 14252 40964 14308 41020
rect 1810 40908 1820 40964
rect 1876 40908 2828 40964
rect 2884 40908 3052 40964
rect 3108 40908 4508 40964
rect 4564 40908 4574 40964
rect 6850 40908 6860 40964
rect 6916 40908 11564 40964
rect 11620 40908 11630 40964
rect 12002 40908 12012 40964
rect 12068 40908 14028 40964
rect 14084 40908 14094 40964
rect 14252 40908 14812 40964
rect 14868 40908 14878 40964
rect 17938 40908 17948 40964
rect 18004 40908 18508 40964
rect 18564 40908 18574 40964
rect 19516 40908 19740 40964
rect 19796 40908 19806 40964
rect 21970 40908 21980 40964
rect 22036 40908 22204 40964
rect 22260 40908 22270 40964
rect 29362 40908 29372 40964
rect 29428 40908 29596 40964
rect 29652 40908 29662 40964
rect 30034 40908 30044 40964
rect 30100 40908 30380 40964
rect 30436 40908 30604 40964
rect 30660 40908 31052 40964
rect 31108 40908 37100 40964
rect 37156 40908 37166 40964
rect 39890 40908 39900 40964
rect 39956 40908 40460 40964
rect 40516 40908 40684 40964
rect 40740 40908 40750 40964
rect 43250 40908 43260 40964
rect 43316 40908 43820 40964
rect 43876 40908 45164 40964
rect 45220 40908 45230 40964
rect 19516 40852 19572 40908
rect 10322 40796 10332 40852
rect 10388 40796 12236 40852
rect 12292 40796 15036 40852
rect 15092 40796 15102 40852
rect 16566 40796 16604 40852
rect 16660 40796 16670 40852
rect 19506 40796 19516 40852
rect 19572 40796 19582 40852
rect 23538 40796 23548 40852
rect 23604 40796 24108 40852
rect 24164 40796 24174 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 4274 40684 4284 40740
rect 4340 40684 4956 40740
rect 5012 40684 5022 40740
rect 8418 40684 8428 40740
rect 8484 40684 8494 40740
rect 11666 40684 11676 40740
rect 11732 40684 16940 40740
rect 16996 40684 17006 40740
rect 17154 40684 17164 40740
rect 17220 40684 17388 40740
rect 17444 40684 17454 40740
rect 23426 40684 23436 40740
rect 23492 40684 25452 40740
rect 25508 40684 26124 40740
rect 26180 40684 26190 40740
rect 27346 40684 27356 40740
rect 27412 40684 33852 40740
rect 33908 40684 33918 40740
rect 1810 40572 1820 40628
rect 1876 40572 3724 40628
rect 3780 40572 3790 40628
rect 2482 40460 2492 40516
rect 2548 40460 6412 40516
rect 6468 40460 7084 40516
rect 7140 40460 7150 40516
rect 8428 40404 8484 40684
rect 8866 40572 8876 40628
rect 8932 40572 9884 40628
rect 9940 40572 9950 40628
rect 11106 40572 11116 40628
rect 11172 40572 25900 40628
rect 25956 40572 26348 40628
rect 26404 40572 26414 40628
rect 26758 40572 26796 40628
rect 26852 40572 26862 40628
rect 28018 40572 28028 40628
rect 28084 40572 28252 40628
rect 28308 40572 28318 40628
rect 34850 40572 34860 40628
rect 34916 40572 36540 40628
rect 36596 40572 36606 40628
rect 40002 40572 40012 40628
rect 40068 40572 40796 40628
rect 40852 40572 42140 40628
rect 42196 40572 42206 40628
rect 43922 40572 43932 40628
rect 43988 40572 45500 40628
rect 45556 40572 45566 40628
rect 11554 40460 11564 40516
rect 11620 40460 12908 40516
rect 12964 40460 13580 40516
rect 13636 40460 13646 40516
rect 15138 40460 15148 40516
rect 15204 40460 16380 40516
rect 16436 40460 16446 40516
rect 16594 40460 16604 40516
rect 16660 40460 20076 40516
rect 20132 40460 20142 40516
rect 28914 40460 28924 40516
rect 28980 40460 29372 40516
rect 29428 40460 29438 40516
rect 31126 40460 31164 40516
rect 31220 40460 31230 40516
rect 33954 40460 33964 40516
rect 34020 40460 34636 40516
rect 34692 40460 34702 40516
rect 41682 40460 41692 40516
rect 41748 40460 43708 40516
rect 43764 40460 44492 40516
rect 44548 40460 44558 40516
rect 45602 40460 45612 40516
rect 45668 40460 47852 40516
rect 47908 40460 47918 40516
rect 59200 40404 59800 40432
rect 8428 40348 8876 40404
rect 8932 40348 9772 40404
rect 9828 40348 9838 40404
rect 13906 40348 13916 40404
rect 13972 40348 13982 40404
rect 15698 40348 15708 40404
rect 15764 40348 15820 40404
rect 15876 40348 15886 40404
rect 16930 40348 16940 40404
rect 16996 40348 20412 40404
rect 20468 40348 20860 40404
rect 20916 40348 20926 40404
rect 21410 40348 21420 40404
rect 21476 40348 21868 40404
rect 21924 40348 21934 40404
rect 22082 40348 22092 40404
rect 22148 40348 22652 40404
rect 22708 40348 22718 40404
rect 23538 40348 23548 40404
rect 23604 40348 34244 40404
rect 36866 40348 36876 40404
rect 36932 40348 37436 40404
rect 37492 40348 37502 40404
rect 42802 40348 42812 40404
rect 42868 40348 43596 40404
rect 43652 40348 44380 40404
rect 44436 40348 44446 40404
rect 45378 40348 45388 40404
rect 45444 40348 46844 40404
rect 46900 40348 46910 40404
rect 55346 40348 55356 40404
rect 55412 40348 59800 40404
rect 13916 40292 13972 40348
rect 34188 40292 34244 40348
rect 59200 40320 59800 40348
rect 2370 40236 2380 40292
rect 2436 40236 4284 40292
rect 4340 40236 4350 40292
rect 7186 40236 7196 40292
rect 7252 40236 10780 40292
rect 10836 40236 10846 40292
rect 13244 40236 13356 40292
rect 13412 40236 13972 40292
rect 14802 40236 14812 40292
rect 14868 40236 15036 40292
rect 15092 40236 15148 40292
rect 15204 40236 15214 40292
rect 18722 40236 18732 40292
rect 18788 40236 19068 40292
rect 19124 40236 20804 40292
rect 20962 40236 20972 40292
rect 21028 40236 23660 40292
rect 23716 40236 23726 40292
rect 34178 40236 34188 40292
rect 34244 40236 34254 40292
rect 40898 40236 40908 40292
rect 40964 40236 41804 40292
rect 41860 40236 41870 40292
rect 13244 40180 13300 40236
rect 20748 40180 20804 40236
rect 7270 40124 7308 40180
rect 7364 40124 7374 40180
rect 9090 40124 9100 40180
rect 9156 40124 13300 40180
rect 19516 40124 20524 40180
rect 20580 40124 20590 40180
rect 20748 40124 22092 40180
rect 22148 40124 22158 40180
rect 19516 40068 19572 40124
rect 4834 40012 4844 40068
rect 4900 40012 11564 40068
rect 11620 40012 12460 40068
rect 12516 40012 12526 40068
rect 13346 40012 13356 40068
rect 13412 40012 13580 40068
rect 13636 40012 13692 40068
rect 13748 40012 13758 40068
rect 13906 40012 13916 40068
rect 13972 40012 13982 40068
rect 19506 40012 19516 40068
rect 19572 40012 19582 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 4844 39900 10052 39956
rect 4844 39844 4900 39900
rect 9996 39844 10052 39900
rect 3714 39788 3724 39844
rect 3780 39788 4900 39844
rect 6850 39788 6860 39844
rect 6916 39788 8540 39844
rect 8596 39788 8606 39844
rect 9986 39788 9996 39844
rect 10052 39788 10668 39844
rect 10724 39788 10734 39844
rect 11666 39788 11676 39844
rect 11732 39788 11742 39844
rect 11676 39732 11732 39788
rect 13916 39732 13972 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 14466 39900 14476 39956
rect 14532 39900 20972 39956
rect 21028 39900 21038 39956
rect 21410 39900 21420 39956
rect 21476 39900 24556 39956
rect 24612 39900 24622 39956
rect 16930 39788 16940 39844
rect 16996 39788 18228 39844
rect 19842 39788 19852 39844
rect 19908 39788 21756 39844
rect 21812 39788 22428 39844
rect 22484 39788 23660 39844
rect 23716 39788 23726 39844
rect 30930 39788 30940 39844
rect 30996 39788 31500 39844
rect 31556 39788 32620 39844
rect 32676 39788 32686 39844
rect 36866 39788 36876 39844
rect 36932 39788 37660 39844
rect 37716 39788 37884 39844
rect 37940 39788 37950 39844
rect 40786 39788 40796 39844
rect 40852 39788 42028 39844
rect 42084 39788 42094 39844
rect 18172 39732 18228 39788
rect 2930 39676 2940 39732
rect 2996 39676 3836 39732
rect 3892 39676 3902 39732
rect 4162 39676 4172 39732
rect 4228 39676 5180 39732
rect 5236 39676 6748 39732
rect 6804 39676 6814 39732
rect 7980 39676 12908 39732
rect 12964 39676 13580 39732
rect 13636 39676 13972 39732
rect 16146 39676 16156 39732
rect 16212 39676 17052 39732
rect 17108 39676 17118 39732
rect 18162 39676 18172 39732
rect 18228 39676 21420 39732
rect 21476 39676 21486 39732
rect 22194 39676 22204 39732
rect 22260 39676 41356 39732
rect 41412 39676 41422 39732
rect 7980 39620 8036 39676
rect 1586 39564 1596 39620
rect 1652 39564 2828 39620
rect 2884 39564 2894 39620
rect 3490 39564 3500 39620
rect 3556 39564 3948 39620
rect 4004 39564 4014 39620
rect 7074 39564 7084 39620
rect 7140 39564 7980 39620
rect 8036 39564 8046 39620
rect 8978 39564 8988 39620
rect 9044 39564 9548 39620
rect 9604 39564 10836 39620
rect 13458 39564 13468 39620
rect 13524 39564 14252 39620
rect 14308 39564 21868 39620
rect 21924 39564 21934 39620
rect 22530 39564 22540 39620
rect 22596 39564 22988 39620
rect 23044 39564 23054 39620
rect 39330 39564 39340 39620
rect 39396 39564 40572 39620
rect 40628 39564 41692 39620
rect 41748 39564 41758 39620
rect 56690 39564 56700 39620
rect 56756 39564 57372 39620
rect 57428 39564 57438 39620
rect 10780 39508 10836 39564
rect 5170 39452 5180 39508
rect 5236 39452 9100 39508
rect 9156 39452 9166 39508
rect 10210 39452 10220 39508
rect 10276 39452 10444 39508
rect 10500 39452 10510 39508
rect 10770 39452 10780 39508
rect 10836 39452 10846 39508
rect 15922 39452 15932 39508
rect 15988 39452 19628 39508
rect 19684 39452 19694 39508
rect 21634 39452 21644 39508
rect 21700 39452 22316 39508
rect 22372 39452 22382 39508
rect 22642 39452 22652 39508
rect 22708 39452 24780 39508
rect 24836 39452 24846 39508
rect 25890 39452 25900 39508
rect 25956 39452 27692 39508
rect 27748 39452 27758 39508
rect 31826 39452 31836 39508
rect 31892 39452 32284 39508
rect 32340 39452 32956 39508
rect 33012 39452 33022 39508
rect 56130 39452 56140 39508
rect 56196 39452 57148 39508
rect 57204 39452 57214 39508
rect 3602 39340 3612 39396
rect 3668 39340 8204 39396
rect 8260 39340 8270 39396
rect 8418 39340 8428 39396
rect 8484 39340 12348 39396
rect 12404 39340 13692 39396
rect 13748 39340 13758 39396
rect 17826 39340 17836 39396
rect 17892 39340 23100 39396
rect 23156 39340 23166 39396
rect 8204 39284 8260 39340
rect 4946 39228 4956 39284
rect 5012 39228 5022 39284
rect 7634 39228 7644 39284
rect 7700 39228 7756 39284
rect 7812 39228 7980 39284
rect 8036 39228 8046 39284
rect 8204 39228 8876 39284
rect 8932 39228 9772 39284
rect 9828 39228 9838 39284
rect 10098 39228 10108 39284
rect 10164 39228 10220 39284
rect 10276 39228 10556 39284
rect 10612 39228 10622 39284
rect 11218 39228 11228 39284
rect 11284 39228 15484 39284
rect 15540 39228 19628 39284
rect 19684 39228 19694 39284
rect 4956 39172 5012 39228
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 3154 39116 3164 39172
rect 3220 39116 3836 39172
rect 3892 39116 3902 39172
rect 4956 39116 7924 39172
rect 8306 39116 8316 39172
rect 8372 39116 9996 39172
rect 10052 39116 10062 39172
rect 10434 39116 10444 39172
rect 10500 39116 12572 39172
rect 12628 39116 12638 39172
rect 18582 39116 18620 39172
rect 18676 39116 18686 39172
rect 32498 39116 32508 39172
rect 32564 39116 32574 39172
rect 36978 39116 36988 39172
rect 37044 39116 37772 39172
rect 37828 39116 38108 39172
rect 38164 39116 38174 39172
rect 200 39060 800 39088
rect 200 39004 1932 39060
rect 1988 39004 1998 39060
rect 2594 39004 2604 39060
rect 2660 39004 4172 39060
rect 4228 39004 7084 39060
rect 7140 39004 7150 39060
rect 200 38976 800 39004
rect 7868 38948 7924 39116
rect 32508 39060 32564 39116
rect 8082 39004 8092 39060
rect 8148 39004 15708 39060
rect 15764 39004 15774 39060
rect 16482 39004 16492 39060
rect 16548 39004 17724 39060
rect 17780 39004 17790 39060
rect 25330 39004 25340 39060
rect 25396 39004 25676 39060
rect 25732 39004 25742 39060
rect 28354 39004 28364 39060
rect 28420 39004 28430 39060
rect 30034 39004 30044 39060
rect 30100 39004 30380 39060
rect 30436 39004 30884 39060
rect 32162 39004 32172 39060
rect 32228 39004 32564 39060
rect 36866 39004 36876 39060
rect 36932 39004 37828 39060
rect 28364 38948 28420 39004
rect 1810 38892 1820 38948
rect 1876 38892 3612 38948
rect 3668 38892 3678 38948
rect 3826 38892 3836 38948
rect 3892 38892 7196 38948
rect 7252 38892 7262 38948
rect 7868 38892 9884 38948
rect 9940 38892 9950 38948
rect 10098 38892 10108 38948
rect 10164 38892 11116 38948
rect 11172 38892 13468 38948
rect 13524 38892 14252 38948
rect 14308 38892 14318 38948
rect 14578 38892 14588 38948
rect 14644 38892 14924 38948
rect 14980 38892 14990 38948
rect 16342 38892 16380 38948
rect 16436 38892 16446 38948
rect 20962 38892 20972 38948
rect 21028 38892 23212 38948
rect 23268 38892 23278 38948
rect 25788 38892 26012 38948
rect 26068 38892 26684 38948
rect 26740 38892 27580 38948
rect 27636 38892 28700 38948
rect 28756 38892 28766 38948
rect 25788 38836 25844 38892
rect 1922 38780 1932 38836
rect 1988 38780 3164 38836
rect 3220 38780 3230 38836
rect 4274 38780 4284 38836
rect 4340 38780 5740 38836
rect 5796 38780 5806 38836
rect 8642 38780 8652 38836
rect 8708 38780 12684 38836
rect 12740 38780 12750 38836
rect 16930 38780 16940 38836
rect 16996 38780 20748 38836
rect 20804 38780 20814 38836
rect 21634 38780 21644 38836
rect 21700 38780 25788 38836
rect 25844 38780 25854 38836
rect 26450 38780 26460 38836
rect 26516 38780 26526 38836
rect 27346 38780 27356 38836
rect 27412 38780 28476 38836
rect 28532 38780 28542 38836
rect 26460 38724 26516 38780
rect 30828 38724 30884 39004
rect 32498 38892 32508 38948
rect 32564 38892 33740 38948
rect 33796 38892 34972 38948
rect 35028 38892 35532 38948
rect 35588 38892 35598 38948
rect 37772 38724 37828 39004
rect 38556 38780 40012 38836
rect 40068 38780 40078 38836
rect 2370 38668 2380 38724
rect 2436 38668 5012 38724
rect 5170 38668 5180 38724
rect 5236 38668 9884 38724
rect 9940 38668 9950 38724
rect 12002 38668 12012 38724
rect 12068 38668 14140 38724
rect 14196 38668 14206 38724
rect 16716 38668 17724 38724
rect 17780 38668 17790 38724
rect 20626 38668 20636 38724
rect 20692 38668 21420 38724
rect 21476 38668 21486 38724
rect 22642 38668 22652 38724
rect 22708 38668 23212 38724
rect 23268 38668 23278 38724
rect 24658 38668 24668 38724
rect 24724 38668 25564 38724
rect 25620 38668 26516 38724
rect 28130 38668 28140 38724
rect 28196 38668 28812 38724
rect 28868 38668 28878 38724
rect 30818 38668 30828 38724
rect 30884 38668 30894 38724
rect 31014 38668 31052 38724
rect 31108 38668 31118 38724
rect 37762 38668 37772 38724
rect 37828 38668 37838 38724
rect 4956 38500 5012 38668
rect 16716 38612 16772 38668
rect 38556 38612 38612 38780
rect 39554 38668 39564 38724
rect 39620 38668 40460 38724
rect 40516 38668 40526 38724
rect 6000 38556 6076 38612
rect 6132 38556 7420 38612
rect 7476 38556 9380 38612
rect 9986 38556 9996 38612
rect 10052 38556 16044 38612
rect 16100 38556 16772 38612
rect 38546 38556 38556 38612
rect 38612 38556 38622 38612
rect 9324 38500 9380 38556
rect 2146 38444 2156 38500
rect 2212 38444 2716 38500
rect 2772 38444 3500 38500
rect 3556 38444 3566 38500
rect 4956 38444 5180 38500
rect 5236 38444 7868 38500
rect 7924 38444 7980 38500
rect 8036 38444 9100 38500
rect 9156 38444 9166 38500
rect 9324 38444 13468 38500
rect 13524 38444 13534 38500
rect 14690 38444 14700 38500
rect 14756 38444 28812 38500
rect 28868 38444 29820 38500
rect 29876 38444 31052 38500
rect 31108 38444 31276 38500
rect 31332 38444 32284 38500
rect 32340 38444 33516 38500
rect 33572 38444 33582 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 5954 38332 5964 38388
rect 6020 38332 8204 38388
rect 8260 38332 8270 38388
rect 12674 38332 12684 38388
rect 12740 38332 22540 38388
rect 22596 38332 23660 38388
rect 23716 38332 23726 38388
rect 26002 38332 26012 38388
rect 26068 38332 26572 38388
rect 26628 38332 26638 38388
rect 39330 38332 39340 38388
rect 39396 38332 42364 38388
rect 42420 38332 42430 38388
rect 7186 38220 7196 38276
rect 7252 38220 7308 38276
rect 7364 38220 7374 38276
rect 12338 38220 12348 38276
rect 12404 38220 16940 38276
rect 16996 38220 17006 38276
rect 19058 38220 19068 38276
rect 19124 38220 23716 38276
rect 26674 38220 26684 38276
rect 26740 38220 27244 38276
rect 27300 38220 28364 38276
rect 28420 38220 28430 38276
rect 38612 38220 39452 38276
rect 39508 38220 39518 38276
rect 23660 38164 23716 38220
rect 38612 38164 38668 38220
rect 3266 38108 3276 38164
rect 3332 38108 5404 38164
rect 5460 38108 7420 38164
rect 7476 38108 7486 38164
rect 8194 38108 8204 38164
rect 8260 38108 12796 38164
rect 12852 38108 12862 38164
rect 13570 38108 13580 38164
rect 13636 38108 15372 38164
rect 15428 38108 15438 38164
rect 18722 38108 18732 38164
rect 18788 38108 20300 38164
rect 20356 38108 22204 38164
rect 22260 38108 23436 38164
rect 23492 38108 23502 38164
rect 23660 38108 29316 38164
rect 29474 38108 29484 38164
rect 29540 38108 36764 38164
rect 36820 38108 38668 38164
rect 41906 38108 41916 38164
rect 41972 38108 42588 38164
rect 42644 38108 42654 38164
rect 12796 38052 12852 38108
rect 29260 38052 29316 38108
rect 7046 37996 7084 38052
rect 7140 37996 7150 38052
rect 7522 37996 7532 38052
rect 7588 37996 8540 38052
rect 8596 37996 11788 38052
rect 11844 37996 12236 38052
rect 12292 37996 12302 38052
rect 12796 37996 14028 38052
rect 14084 37996 14094 38052
rect 15586 37996 15596 38052
rect 15652 37996 15662 38052
rect 16594 37996 16604 38052
rect 16660 37996 17500 38052
rect 17556 37996 17566 38052
rect 23650 37996 23660 38052
rect 23716 37996 24444 38052
rect 24500 37996 24510 38052
rect 26562 37996 26572 38052
rect 26628 37996 27356 38052
rect 27412 37996 27422 38052
rect 29260 37996 29596 38052
rect 29652 37996 30044 38052
rect 30100 37996 30604 38052
rect 30660 37996 31052 38052
rect 31108 37996 33068 38052
rect 33124 37996 33964 38052
rect 34020 37996 34030 38052
rect 41682 37996 41692 38052
rect 41748 37996 42364 38052
rect 42420 37996 42430 38052
rect 15596 37940 15652 37996
rect 2370 37884 2380 37940
rect 2436 37884 3388 37940
rect 5730 37884 5740 37940
rect 5796 37884 5852 37940
rect 5908 37884 7364 37940
rect 9202 37884 9212 37940
rect 9268 37884 11676 37940
rect 11732 37884 13692 37940
rect 13748 37884 13758 37940
rect 15148 37884 16044 37940
rect 16100 37884 16492 37940
rect 16548 37884 16940 37940
rect 16996 37884 18900 37940
rect 19254 37884 19292 37940
rect 19348 37884 19358 37940
rect 19618 37884 19628 37940
rect 19684 37884 20636 37940
rect 20692 37884 20702 37940
rect 20850 37884 20860 37940
rect 20916 37884 21644 37940
rect 21700 37884 21710 37940
rect 30818 37884 30828 37940
rect 30884 37884 31388 37940
rect 31444 37884 32060 37940
rect 32116 37884 32126 37940
rect 3332 37716 3388 37884
rect 7308 37828 7364 37884
rect 15148 37828 15204 37884
rect 18844 37828 18900 37884
rect 20860 37828 20916 37884
rect 3938 37772 3948 37828
rect 4004 37772 4956 37828
rect 5012 37772 5022 37828
rect 5170 37772 5180 37828
rect 5236 37772 5852 37828
rect 5908 37772 5918 37828
rect 7298 37772 7308 37828
rect 7364 37772 10108 37828
rect 10164 37772 10174 37828
rect 12310 37772 12348 37828
rect 12404 37772 12414 37828
rect 15138 37772 15148 37828
rect 15204 37772 15214 37828
rect 15596 37772 16604 37828
rect 16660 37772 16670 37828
rect 18844 37772 18956 37828
rect 19012 37772 20916 37828
rect 23314 37772 23324 37828
rect 23380 37772 24892 37828
rect 24948 37772 24958 37828
rect 25778 37772 25788 37828
rect 25844 37772 26684 37828
rect 26740 37772 26750 37828
rect 15596 37716 15652 37772
rect 3332 37660 6972 37716
rect 7028 37660 7038 37716
rect 9874 37660 9884 37716
rect 9940 37660 11228 37716
rect 11284 37660 11564 37716
rect 11620 37660 15652 37716
rect 15810 37660 15820 37716
rect 15876 37660 19628 37716
rect 19684 37660 19694 37716
rect 22530 37660 22540 37716
rect 22596 37660 23996 37716
rect 24052 37660 24276 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 24220 37604 24276 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 24210 37548 24220 37604
rect 24276 37548 24286 37604
rect 28242 37548 28252 37604
rect 28308 37548 37548 37604
rect 37604 37548 37996 37604
rect 38052 37548 38332 37604
rect 38388 37548 38398 37604
rect 6962 37436 6972 37492
rect 7028 37436 9884 37492
rect 9940 37436 12572 37492
rect 12628 37436 13020 37492
rect 13076 37436 13086 37492
rect 15586 37436 15596 37492
rect 15652 37436 16716 37492
rect 16772 37436 16940 37492
rect 16996 37436 17006 37492
rect 17490 37436 17500 37492
rect 17556 37436 21700 37492
rect 23762 37436 23772 37492
rect 23828 37436 29932 37492
rect 29988 37436 29998 37492
rect 21644 37380 21700 37436
rect 1698 37324 1708 37380
rect 1764 37324 2716 37380
rect 2772 37324 3500 37380
rect 3556 37324 3566 37380
rect 5954 37324 5964 37380
rect 6020 37324 7196 37380
rect 7252 37324 7262 37380
rect 8978 37324 8988 37380
rect 9044 37324 10444 37380
rect 10500 37324 10510 37380
rect 20626 37324 20636 37380
rect 20692 37324 21420 37380
rect 21476 37324 21486 37380
rect 21634 37324 21644 37380
rect 21700 37324 23324 37380
rect 23380 37324 23390 37380
rect 3266 37212 3276 37268
rect 3332 37212 4508 37268
rect 4564 37212 4956 37268
rect 5012 37212 5022 37268
rect 6710 37212 6748 37268
rect 6804 37212 6814 37268
rect 6962 37212 6972 37268
rect 7028 37212 7644 37268
rect 7700 37212 13356 37268
rect 13412 37212 14252 37268
rect 14308 37212 14318 37268
rect 17826 37212 17836 37268
rect 17892 37212 18620 37268
rect 18676 37212 18686 37268
rect 19394 37212 19404 37268
rect 19460 37212 20076 37268
rect 20132 37212 21980 37268
rect 22036 37212 22046 37268
rect 26226 37212 26236 37268
rect 26292 37212 28140 37268
rect 28196 37212 28206 37268
rect 35074 37212 35084 37268
rect 35140 37212 35644 37268
rect 35700 37212 35710 37268
rect 10518 37100 10556 37156
rect 10612 37100 11900 37156
rect 11956 37100 11966 37156
rect 26674 37100 26684 37156
rect 26740 37100 27468 37156
rect 27524 37100 28476 37156
rect 28532 37100 29148 37156
rect 29204 37100 29214 37156
rect 4284 36988 4900 37044
rect 6290 36988 6300 37044
rect 6356 36988 15820 37044
rect 15876 36988 16884 37044
rect 22642 36988 22652 37044
rect 22708 36988 23212 37044
rect 23268 36988 23278 37044
rect 26450 36988 26460 37044
rect 26516 36988 27244 37044
rect 27300 36988 27916 37044
rect 27972 36988 27982 37044
rect 34972 36988 35868 37044
rect 35924 36988 35934 37044
rect 43026 36988 43036 37044
rect 43092 36988 54908 37044
rect 54964 36988 54974 37044
rect 4284 36932 4340 36988
rect 3332 36876 4340 36932
rect 4844 36932 4900 36988
rect 16828 36932 16884 36988
rect 34972 36932 35028 36988
rect 4844 36876 6076 36932
rect 6132 36876 6142 36932
rect 7382 36876 7420 36932
rect 7476 36876 7486 36932
rect 10658 36876 10668 36932
rect 10724 36876 16604 36932
rect 16660 36876 16670 36932
rect 16828 36876 19068 36932
rect 19124 36876 19134 36932
rect 26226 36876 26236 36932
rect 26292 36876 26908 36932
rect 26964 36876 26974 36932
rect 27468 36876 35028 36932
rect 41122 36876 41132 36932
rect 41188 36876 41804 36932
rect 41860 36876 42476 36932
rect 42532 36876 42542 36932
rect 3332 36708 3388 36876
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 6934 36764 6972 36820
rect 7028 36764 7038 36820
rect 17714 36764 17724 36820
rect 17780 36764 19852 36820
rect 19908 36764 19918 36820
rect 1922 36652 1932 36708
rect 1988 36652 3388 36708
rect 4050 36652 4060 36708
rect 4116 36652 6860 36708
rect 6916 36652 6926 36708
rect 16146 36652 16156 36708
rect 16212 36652 21868 36708
rect 21924 36652 21934 36708
rect 4060 36596 4116 36652
rect 1810 36540 1820 36596
rect 1876 36540 4116 36596
rect 6066 36540 6076 36596
rect 6132 36540 7532 36596
rect 7588 36540 7598 36596
rect 9202 36540 9212 36596
rect 9268 36540 11900 36596
rect 11956 36540 12236 36596
rect 12292 36540 17164 36596
rect 17220 36540 17230 36596
rect 17714 36540 17724 36596
rect 17780 36540 20972 36596
rect 21028 36540 21038 36596
rect 25666 36540 25676 36596
rect 25732 36540 26236 36596
rect 26292 36540 26302 36596
rect 27468 36484 27524 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 28690 36764 28700 36820
rect 28756 36764 29596 36820
rect 29652 36764 31276 36820
rect 31332 36764 31342 36820
rect 27682 36652 27692 36708
rect 27748 36652 33964 36708
rect 34020 36652 34860 36708
rect 34916 36652 34926 36708
rect 35084 36652 36988 36708
rect 37044 36652 37054 36708
rect 35084 36596 35140 36652
rect 30818 36540 30828 36596
rect 30884 36540 31948 36596
rect 32004 36540 35140 36596
rect 35746 36540 35756 36596
rect 35812 36540 38668 36596
rect 38724 36540 38734 36596
rect 43138 36540 43148 36596
rect 43204 36540 45612 36596
rect 45668 36540 45678 36596
rect 6402 36428 6412 36484
rect 6468 36428 6748 36484
rect 6804 36428 8092 36484
rect 8148 36428 8158 36484
rect 8306 36428 8316 36484
rect 8372 36428 10220 36484
rect 10276 36428 10556 36484
rect 10612 36428 10622 36484
rect 12898 36428 12908 36484
rect 12964 36428 15036 36484
rect 15092 36428 16268 36484
rect 16324 36428 16334 36484
rect 16482 36428 16492 36484
rect 16548 36428 27524 36484
rect 28802 36428 28812 36484
rect 28868 36428 30492 36484
rect 30548 36428 30558 36484
rect 32834 36428 32844 36484
rect 32900 36428 33628 36484
rect 33684 36428 35420 36484
rect 35476 36428 35486 36484
rect 40114 36428 40124 36484
rect 40180 36428 41356 36484
rect 41412 36428 41422 36484
rect 2370 36316 2380 36372
rect 2436 36316 2940 36372
rect 2996 36316 3006 36372
rect 3266 36316 3276 36372
rect 3332 36316 4172 36372
rect 4228 36316 4508 36372
rect 4564 36316 4574 36372
rect 6290 36316 6300 36372
rect 6356 36316 10668 36372
rect 10724 36316 10734 36372
rect 14018 36316 14028 36372
rect 14084 36316 15484 36372
rect 15540 36316 15550 36372
rect 15698 36316 15708 36372
rect 15764 36316 16156 36372
rect 16212 36316 16222 36372
rect 18498 36316 18508 36372
rect 18564 36316 19180 36372
rect 19236 36316 19246 36372
rect 19618 36316 19628 36372
rect 19684 36316 23100 36372
rect 23156 36316 23166 36372
rect 23650 36316 23660 36372
rect 23716 36316 24556 36372
rect 24612 36316 24622 36372
rect 29026 36316 29036 36372
rect 29092 36316 29708 36372
rect 29764 36316 29774 36372
rect 33170 36316 33180 36372
rect 33236 36316 33740 36372
rect 33796 36316 34748 36372
rect 34804 36316 34814 36372
rect 36754 36316 36764 36372
rect 36820 36316 39228 36372
rect 39284 36316 42140 36372
rect 42196 36316 42364 36372
rect 42420 36316 42430 36372
rect 6300 36260 6356 36316
rect 3938 36204 3948 36260
rect 4004 36204 6356 36260
rect 7074 36204 7084 36260
rect 7140 36204 17164 36260
rect 17220 36204 18284 36260
rect 18340 36204 18350 36260
rect 19030 36204 19068 36260
rect 19124 36204 19134 36260
rect 19628 36204 19852 36260
rect 19908 36204 20524 36260
rect 20580 36204 20590 36260
rect 20850 36204 20860 36260
rect 20916 36204 21644 36260
rect 21700 36204 21710 36260
rect 22642 36204 22652 36260
rect 22708 36204 25452 36260
rect 25508 36204 25518 36260
rect 28130 36204 28140 36260
rect 28196 36204 28812 36260
rect 28868 36204 28878 36260
rect 29558 36204 29596 36260
rect 29652 36204 29662 36260
rect 30594 36204 30604 36260
rect 30660 36204 38444 36260
rect 38500 36204 38510 36260
rect 38658 36204 38668 36260
rect 38724 36204 41468 36260
rect 41524 36204 41804 36260
rect 41860 36204 41870 36260
rect 2482 36092 2492 36148
rect 2548 36092 3052 36148
rect 3108 36092 3118 36148
rect 5254 36092 5292 36148
rect 5348 36092 5358 36148
rect 7084 36036 7140 36204
rect 19628 36148 19684 36204
rect 12450 36092 12460 36148
rect 12516 36092 13020 36148
rect 13076 36092 13086 36148
rect 13458 36092 13468 36148
rect 13524 36092 14364 36148
rect 14420 36092 14430 36148
rect 14998 36092 15036 36148
rect 15092 36092 15102 36148
rect 16258 36092 16268 36148
rect 16324 36092 17388 36148
rect 17444 36092 17454 36148
rect 19618 36092 19628 36148
rect 19684 36092 19694 36148
rect 21858 36092 21868 36148
rect 21924 36092 33068 36148
rect 33124 36092 33134 36148
rect 33702 36092 33740 36148
rect 33796 36092 33806 36148
rect 33954 36092 33964 36148
rect 34020 36092 34636 36148
rect 34692 36092 34702 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 2268 35980 7140 36036
rect 11666 35980 11676 36036
rect 11732 35980 12012 36036
rect 12068 35980 12908 36036
rect 12964 35980 12974 36036
rect 13234 35980 13244 36036
rect 13300 35980 18844 36036
rect 18900 35980 18910 36036
rect 38434 35980 38444 36036
rect 38500 35980 39004 36036
rect 39060 35980 41132 36036
rect 41188 35980 41198 36036
rect 2268 35924 2324 35980
rect 1474 35868 1484 35924
rect 1540 35868 2268 35924
rect 2324 35868 2334 35924
rect 4722 35868 4732 35924
rect 4788 35868 5740 35924
rect 5796 35868 6748 35924
rect 6804 35868 6814 35924
rect 9986 35868 9996 35924
rect 10052 35868 11564 35924
rect 11620 35868 15148 35924
rect 15092 35812 15148 35868
rect 16716 35868 17276 35924
rect 17332 35868 17342 35924
rect 21634 35868 21644 35924
rect 21700 35868 21756 35924
rect 21812 35868 21822 35924
rect 35410 35868 35420 35924
rect 35476 35868 36092 35924
rect 36148 35868 36158 35924
rect 47842 35868 47852 35924
rect 47908 35868 54348 35924
rect 54404 35868 54908 35924
rect 54964 35868 54974 35924
rect 6514 35756 6524 35812
rect 6580 35756 8428 35812
rect 8484 35756 8876 35812
rect 8932 35756 9548 35812
rect 9604 35756 9614 35812
rect 9762 35756 9772 35812
rect 9828 35756 11004 35812
rect 11060 35756 11070 35812
rect 11890 35756 11900 35812
rect 11956 35756 13132 35812
rect 13188 35756 14084 35812
rect 15092 35756 16268 35812
rect 16324 35756 16334 35812
rect 9772 35700 9828 35756
rect 14028 35700 14084 35756
rect 8642 35644 8652 35700
rect 8708 35644 9100 35700
rect 9156 35644 9828 35700
rect 11442 35644 11452 35700
rect 11508 35644 12124 35700
rect 12180 35644 12190 35700
rect 14018 35644 14028 35700
rect 14084 35644 14812 35700
rect 14868 35644 14878 35700
rect 16716 35588 16772 35868
rect 17042 35756 17052 35812
rect 17108 35756 17724 35812
rect 17780 35756 17790 35812
rect 19058 35756 19068 35812
rect 19124 35756 21532 35812
rect 21588 35756 21598 35812
rect 32722 35756 32732 35812
rect 32788 35756 33628 35812
rect 33684 35756 33694 35812
rect 43652 35756 52780 35812
rect 52836 35756 52846 35812
rect 16930 35644 16940 35700
rect 16996 35644 18172 35700
rect 18228 35644 18844 35700
rect 18900 35644 19404 35700
rect 19460 35644 19470 35700
rect 32050 35644 32060 35700
rect 32116 35644 32620 35700
rect 32676 35644 33852 35700
rect 33908 35644 33918 35700
rect 34066 35644 34076 35700
rect 34132 35644 38668 35700
rect 7970 35532 7980 35588
rect 8036 35532 8764 35588
rect 8820 35532 8830 35588
rect 11330 35532 11340 35588
rect 11396 35532 15596 35588
rect 15652 35532 19180 35588
rect 19236 35532 19246 35588
rect 28578 35532 28588 35588
rect 28644 35532 28924 35588
rect 28980 35532 28990 35588
rect 30034 35532 30044 35588
rect 30100 35532 30268 35588
rect 30324 35532 30716 35588
rect 30772 35532 31388 35588
rect 31444 35532 31454 35588
rect 33954 35532 33964 35588
rect 34020 35532 34412 35588
rect 34468 35532 34972 35588
rect 35028 35532 35868 35588
rect 35924 35532 35934 35588
rect 38612 35476 38668 35644
rect 43652 35476 43708 35756
rect 3490 35420 3500 35476
rect 3556 35420 5628 35476
rect 5684 35420 5694 35476
rect 8866 35420 8876 35476
rect 8932 35420 9660 35476
rect 9716 35420 12460 35476
rect 12516 35420 12526 35476
rect 16034 35420 16044 35476
rect 16100 35420 17556 35476
rect 19954 35420 19964 35476
rect 20020 35420 23548 35476
rect 23604 35420 23614 35476
rect 24658 35420 24668 35476
rect 24724 35420 25004 35476
rect 25060 35420 25564 35476
rect 25620 35420 27692 35476
rect 27748 35420 34076 35476
rect 34132 35420 34142 35476
rect 34850 35420 34860 35476
rect 34916 35420 35644 35476
rect 35700 35420 36316 35476
rect 36372 35420 36382 35476
rect 38612 35420 43708 35476
rect 17500 35364 17556 35420
rect 4834 35308 4844 35364
rect 4900 35308 4956 35364
rect 5012 35308 10332 35364
rect 10388 35308 10398 35364
rect 10556 35308 15260 35364
rect 15316 35308 15596 35364
rect 15652 35308 16492 35364
rect 16548 35308 16558 35364
rect 16706 35308 16716 35364
rect 16772 35308 16940 35364
rect 16996 35308 17006 35364
rect 17490 35308 17500 35364
rect 17556 35308 18396 35364
rect 18452 35308 18462 35364
rect 21746 35308 21756 35364
rect 21812 35308 22092 35364
rect 22148 35308 23436 35364
rect 23492 35308 23502 35364
rect 28588 35308 29932 35364
rect 29988 35308 29998 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 10556 35252 10612 35308
rect 28588 35252 28644 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 2818 35196 2828 35252
rect 2884 35196 2940 35252
rect 2996 35196 3006 35252
rect 5058 35196 5068 35252
rect 5124 35196 5516 35252
rect 5572 35196 5582 35252
rect 10210 35196 10220 35252
rect 10276 35196 10612 35252
rect 12898 35196 12908 35252
rect 12964 35196 18732 35252
rect 18788 35196 20524 35252
rect 20580 35196 20590 35252
rect 21074 35196 21084 35252
rect 21140 35196 21868 35252
rect 21924 35196 22652 35252
rect 22708 35196 22718 35252
rect 23986 35196 23996 35252
rect 24052 35196 24780 35252
rect 24836 35196 26348 35252
rect 26404 35196 26414 35252
rect 28578 35196 28588 35252
rect 28644 35196 28654 35252
rect 2706 35084 2716 35140
rect 2772 35084 3164 35140
rect 3220 35084 7308 35140
rect 7364 35084 7644 35140
rect 7700 35084 8092 35140
rect 8148 35084 8988 35140
rect 9044 35084 9324 35140
rect 9380 35084 9884 35140
rect 9940 35084 9950 35140
rect 12572 35084 35756 35140
rect 35812 35084 35822 35140
rect 12572 35028 12628 35084
rect 59200 35028 59800 35056
rect 3490 34972 3500 35028
rect 3556 34972 5292 35028
rect 5348 34972 9716 35028
rect 9874 34972 9884 35028
rect 9940 34972 12572 35028
rect 12628 34972 12638 35028
rect 14914 34972 14924 35028
rect 14980 34972 15708 35028
rect 15764 34972 15774 35028
rect 26002 34972 26012 35028
rect 26068 34972 26908 35028
rect 26964 34972 26974 35028
rect 56018 34972 56028 35028
rect 56084 34972 59800 35028
rect 9660 34916 9716 34972
rect 59200 34944 59800 34972
rect 2146 34860 2156 34916
rect 2212 34860 3388 34916
rect 4722 34860 4732 34916
rect 4788 34860 5852 34916
rect 5908 34860 6188 34916
rect 6244 34860 6254 34916
rect 9660 34860 10780 34916
rect 10836 34860 11116 34916
rect 11172 34860 11182 34916
rect 11330 34860 11340 34916
rect 11396 34860 11676 34916
rect 11732 34860 11742 34916
rect 14018 34860 14028 34916
rect 14084 34860 16380 34916
rect 16436 34860 16446 34916
rect 22754 34860 22764 34916
rect 22820 34860 24668 34916
rect 24724 34860 24734 34916
rect 32498 34860 32508 34916
rect 32564 34860 47068 34916
rect 47124 34860 47134 34916
rect 3332 34804 3388 34860
rect 3332 34748 5852 34804
rect 5908 34748 5918 34804
rect 8194 34748 8204 34804
rect 8260 34748 9100 34804
rect 9156 34748 9166 34804
rect 10546 34748 10556 34804
rect 10612 34748 11452 34804
rect 11508 34748 12796 34804
rect 12852 34748 12862 34804
rect 15810 34748 15820 34804
rect 15876 34748 16044 34804
rect 16100 34748 16110 34804
rect 16258 34748 16268 34804
rect 16324 34748 16604 34804
rect 16660 34748 16670 34804
rect 18386 34748 18396 34804
rect 18452 34748 20076 34804
rect 20132 34748 20142 34804
rect 23874 34748 23884 34804
rect 23940 34748 24556 34804
rect 24612 34748 24622 34804
rect 1810 34636 1820 34692
rect 1876 34636 2604 34692
rect 2660 34636 5740 34692
rect 5796 34636 6860 34692
rect 6916 34636 12572 34692
rect 12628 34636 12638 34692
rect 31714 34636 31724 34692
rect 31780 34636 32732 34692
rect 32788 34636 32798 34692
rect 34178 34636 34188 34692
rect 34244 34636 39004 34692
rect 39060 34636 40460 34692
rect 40516 34636 40526 34692
rect 52882 34636 52892 34692
rect 52948 34636 54796 34692
rect 54852 34636 54862 34692
rect 4918 34524 4956 34580
rect 5012 34524 5022 34580
rect 14690 34524 14700 34580
rect 14756 34524 16156 34580
rect 16212 34524 16940 34580
rect 16996 34524 18732 34580
rect 18788 34524 19292 34580
rect 19348 34524 19358 34580
rect 43586 34524 43596 34580
rect 43652 34524 49532 34580
rect 49588 34524 50092 34580
rect 50148 34524 50158 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 4956 34412 5180 34468
rect 5236 34412 5246 34468
rect 5506 34412 5516 34468
rect 5572 34412 6188 34468
rect 6244 34412 11676 34468
rect 11732 34412 13804 34468
rect 13860 34412 13870 34468
rect 21634 34412 21644 34468
rect 21700 34412 23212 34468
rect 23268 34412 24444 34468
rect 24500 34412 24510 34468
rect 30482 34412 30492 34468
rect 30548 34412 36764 34468
rect 36820 34412 37100 34468
rect 37156 34412 37166 34468
rect 4956 34356 5012 34412
rect 3602 34300 3612 34356
rect 3668 34300 4396 34356
rect 4452 34300 4462 34356
rect 4946 34300 4956 34356
rect 5012 34300 5022 34356
rect 5366 34300 5404 34356
rect 5460 34300 5470 34356
rect 6262 34300 6300 34356
rect 6356 34300 6366 34356
rect 9874 34300 9884 34356
rect 9940 34300 10556 34356
rect 10612 34300 10622 34356
rect 12562 34300 12572 34356
rect 12628 34300 14028 34356
rect 14084 34300 14094 34356
rect 15698 34300 15708 34356
rect 15764 34300 18284 34356
rect 18340 34300 18350 34356
rect 24658 34300 24668 34356
rect 24724 34300 25228 34356
rect 25284 34300 25564 34356
rect 25620 34300 25630 34356
rect 28242 34300 28252 34356
rect 28308 34300 30940 34356
rect 30996 34300 31276 34356
rect 31332 34300 31342 34356
rect 32722 34300 32732 34356
rect 32788 34300 37212 34356
rect 37268 34300 37772 34356
rect 37828 34300 37838 34356
rect 5506 34188 5516 34244
rect 5572 34188 5740 34244
rect 5796 34188 5806 34244
rect 7634 34188 7644 34244
rect 7700 34188 17948 34244
rect 18004 34188 18620 34244
rect 18676 34188 22932 34244
rect 23090 34188 23100 34244
rect 23156 34188 23996 34244
rect 24052 34188 24062 34244
rect 24546 34188 24556 34244
rect 24612 34188 39340 34244
rect 39396 34188 39406 34244
rect 22876 34132 22932 34188
rect 3378 34076 3388 34132
rect 3444 34076 4172 34132
rect 4228 34076 4238 34132
rect 11554 34076 11564 34132
rect 11620 34076 13468 34132
rect 13524 34076 13534 34132
rect 13794 34076 13804 34132
rect 13860 34076 14364 34132
rect 14420 34076 16044 34132
rect 16100 34076 19740 34132
rect 19796 34076 19806 34132
rect 20178 34076 20188 34132
rect 20244 34076 21868 34132
rect 21924 34076 22428 34132
rect 22484 34076 22494 34132
rect 22876 34076 23884 34132
rect 23940 34076 23950 34132
rect 26898 34076 26908 34132
rect 26964 34076 27804 34132
rect 27860 34076 28364 34132
rect 28420 34076 29932 34132
rect 29988 34076 29998 34132
rect 30370 34076 30380 34132
rect 30436 34076 31836 34132
rect 31892 34076 31902 34132
rect 19740 34020 19796 34076
rect 3938 33964 3948 34020
rect 4004 33964 13020 34020
rect 13076 33964 14252 34020
rect 14308 33964 14588 34020
rect 14644 33964 14654 34020
rect 19740 33964 20412 34020
rect 20468 33964 20748 34020
rect 20804 33964 21532 34020
rect 21588 33964 21598 34020
rect 22530 33964 22540 34020
rect 22596 33964 24220 34020
rect 24276 33964 28700 34020
rect 28756 33964 29372 34020
rect 29428 33964 29438 34020
rect 31126 33964 31164 34020
rect 31220 33964 31230 34020
rect 36754 33964 36764 34020
rect 36820 33964 38220 34020
rect 38276 33964 42364 34020
rect 42420 33964 42430 34020
rect 2370 33852 2380 33908
rect 2436 33852 2828 33908
rect 2884 33852 6636 33908
rect 6692 33852 7308 33908
rect 7364 33852 7756 33908
rect 7812 33852 8876 33908
rect 8932 33852 8942 33908
rect 2930 33740 2940 33796
rect 2996 33740 3388 33796
rect 14130 33740 14140 33796
rect 14196 33740 26012 33796
rect 26068 33740 26572 33796
rect 26628 33740 26638 33796
rect 200 33684 800 33712
rect 200 33628 1932 33684
rect 1988 33628 1998 33684
rect 2370 33628 2380 33684
rect 2436 33628 3164 33684
rect 3220 33628 3230 33684
rect 200 33600 800 33628
rect 3332 33572 3388 33740
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 8418 33628 8428 33684
rect 8484 33628 11676 33684
rect 11732 33628 11742 33684
rect 14018 33628 14028 33684
rect 14084 33628 14812 33684
rect 14868 33628 14878 33684
rect 27122 33628 27132 33684
rect 27188 33628 28924 33684
rect 28980 33628 28990 33684
rect 29362 33628 29372 33684
rect 29428 33628 30604 33684
rect 30660 33628 31612 33684
rect 31668 33628 31678 33684
rect 46274 33628 46284 33684
rect 46340 33628 52332 33684
rect 52388 33628 52398 33684
rect 31052 33572 31108 33628
rect 3332 33516 9436 33572
rect 9492 33516 9502 33572
rect 13346 33516 13356 33572
rect 13412 33516 30268 33572
rect 30324 33516 30334 33572
rect 31042 33516 31052 33572
rect 31108 33516 31118 33572
rect 38612 33516 43708 33572
rect 43764 33516 43774 33572
rect 38612 33460 38668 33516
rect 1922 33404 1932 33460
rect 1988 33404 3276 33460
rect 3332 33404 4060 33460
rect 4116 33404 4620 33460
rect 4676 33404 4956 33460
rect 5012 33404 5022 33460
rect 11106 33404 11116 33460
rect 11172 33404 38668 33460
rect 43026 33404 43036 33460
rect 43092 33404 44492 33460
rect 44548 33404 44558 33460
rect 3602 33292 3612 33348
rect 3668 33292 12908 33348
rect 12964 33292 13804 33348
rect 13860 33292 13870 33348
rect 14914 33292 14924 33348
rect 14980 33292 16604 33348
rect 16660 33292 16772 33348
rect 16930 33292 16940 33348
rect 16996 33292 17612 33348
rect 17668 33292 17678 33348
rect 30790 33292 30828 33348
rect 30884 33292 30894 33348
rect 33394 33292 33404 33348
rect 33460 33292 36316 33348
rect 36372 33292 37436 33348
rect 37492 33292 37502 33348
rect 37650 33292 37660 33348
rect 37716 33292 39452 33348
rect 39508 33292 41020 33348
rect 41076 33292 41468 33348
rect 41524 33292 41534 33348
rect 5852 33236 5908 33292
rect 16716 33236 16772 33292
rect 3266 33180 3276 33236
rect 3332 33180 3500 33236
rect 3556 33180 3566 33236
rect 5842 33180 5852 33236
rect 5908 33180 5918 33236
rect 6738 33180 6748 33236
rect 6804 33180 7420 33236
rect 7476 33180 7486 33236
rect 16034 33180 16044 33236
rect 16100 33180 16156 33236
rect 16212 33180 16222 33236
rect 16716 33180 17388 33236
rect 17444 33180 17454 33236
rect 21634 33180 21644 33236
rect 21700 33180 22764 33236
rect 22820 33180 22830 33236
rect 31154 33180 31164 33236
rect 31220 33180 31724 33236
rect 31780 33180 31790 33236
rect 41122 33180 41132 33236
rect 41188 33180 46620 33236
rect 46676 33180 47516 33236
rect 47572 33180 47582 33236
rect 8754 33068 8764 33124
rect 8820 33068 12236 33124
rect 12292 33068 12796 33124
rect 12852 33068 12862 33124
rect 14018 33068 14028 33124
rect 14084 33068 23548 33124
rect 23604 33068 24108 33124
rect 24164 33068 24892 33124
rect 24948 33068 24958 33124
rect 27794 33068 27804 33124
rect 27860 33068 32396 33124
rect 32452 33068 33740 33124
rect 33796 33068 34076 33124
rect 34132 33068 34142 33124
rect 2482 32956 2492 33012
rect 2548 32956 3052 33012
rect 3108 32956 3118 33012
rect 7634 32956 7644 33012
rect 7700 32956 15260 33012
rect 15316 32956 15326 33012
rect 15922 32956 15932 33012
rect 15988 32956 16268 33012
rect 16324 32956 16492 33012
rect 16548 32956 16558 33012
rect 30706 32956 30716 33012
rect 30772 32956 31388 33012
rect 31444 32956 32284 33012
rect 32340 32956 32350 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 6066 32844 6076 32900
rect 6132 32844 19292 32900
rect 19348 32844 19358 32900
rect 22978 32844 22988 32900
rect 23044 32844 46732 32900
rect 46788 32844 46798 32900
rect 5618 32732 5628 32788
rect 5684 32732 6412 32788
rect 6468 32732 6478 32788
rect 7186 32732 7196 32788
rect 7252 32732 9548 32788
rect 9604 32732 9614 32788
rect 11638 32732 11676 32788
rect 11732 32732 11742 32788
rect 12786 32732 12796 32788
rect 12852 32732 14140 32788
rect 14196 32732 14206 32788
rect 15138 32732 15148 32788
rect 15204 32732 15932 32788
rect 15988 32732 15998 32788
rect 16818 32732 16828 32788
rect 16884 32732 18172 32788
rect 18228 32732 18956 32788
rect 19012 32732 19022 32788
rect 22054 32732 22092 32788
rect 22148 32732 22876 32788
rect 22932 32732 22942 32788
rect 23100 32732 56588 32788
rect 56644 32732 56654 32788
rect 5628 32676 5684 32732
rect 3266 32620 3276 32676
rect 3332 32620 3612 32676
rect 3668 32620 3678 32676
rect 4284 32620 5684 32676
rect 6412 32676 6468 32732
rect 23100 32676 23156 32732
rect 6412 32620 7980 32676
rect 8036 32620 8046 32676
rect 17266 32620 17276 32676
rect 17332 32620 23156 32676
rect 26002 32620 26012 32676
rect 26068 32620 27804 32676
rect 27860 32620 27870 32676
rect 30370 32620 30380 32676
rect 30436 32620 30940 32676
rect 30996 32620 31006 32676
rect 37538 32620 37548 32676
rect 37604 32620 37996 32676
rect 38052 32620 38062 32676
rect 51650 32620 51660 32676
rect 51716 32620 52668 32676
rect 52724 32620 52734 32676
rect 4284 32564 4340 32620
rect 2930 32508 2940 32564
rect 2996 32508 3276 32564
rect 3332 32508 3948 32564
rect 4004 32508 4014 32564
rect 4274 32508 4284 32564
rect 4340 32508 4350 32564
rect 5394 32508 5404 32564
rect 5460 32508 5964 32564
rect 6020 32508 8988 32564
rect 9044 32508 9996 32564
rect 10052 32508 10062 32564
rect 19506 32508 19516 32564
rect 19572 32508 22652 32564
rect 22708 32508 22718 32564
rect 25666 32508 25676 32564
rect 25732 32508 26460 32564
rect 26516 32508 28476 32564
rect 28532 32508 28542 32564
rect 31602 32508 31612 32564
rect 31668 32508 33516 32564
rect 33572 32508 33582 32564
rect 47506 32508 47516 32564
rect 47572 32508 53900 32564
rect 53956 32508 53966 32564
rect 3378 32396 3388 32452
rect 3444 32396 3612 32452
rect 3668 32396 3678 32452
rect 8530 32396 8540 32452
rect 8596 32396 8764 32452
rect 8820 32396 8830 32452
rect 11890 32396 11900 32452
rect 11956 32396 12572 32452
rect 12628 32396 12638 32452
rect 15250 32396 15260 32452
rect 15316 32396 15708 32452
rect 15764 32396 16604 32452
rect 16660 32396 17612 32452
rect 17668 32396 17678 32452
rect 26852 32396 46172 32452
rect 46228 32396 48076 32452
rect 48132 32396 51100 32452
rect 51156 32396 51996 32452
rect 52052 32396 57372 32452
rect 57428 32396 58380 32452
rect 58436 32396 58446 32452
rect 26852 32340 26908 32396
rect 10322 32284 10332 32340
rect 10388 32284 20188 32340
rect 20244 32284 20860 32340
rect 20916 32284 20926 32340
rect 24994 32284 25004 32340
rect 25060 32284 26908 32340
rect 28242 32284 28252 32340
rect 28308 32284 28924 32340
rect 28980 32284 30380 32340
rect 30436 32284 30446 32340
rect 33394 32284 33404 32340
rect 33460 32284 41132 32340
rect 41188 32284 41198 32340
rect 5618 32172 5628 32228
rect 5684 32172 6412 32228
rect 6468 32172 8652 32228
rect 8708 32172 9884 32228
rect 9940 32172 9950 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 17378 32060 17388 32116
rect 17444 32060 29148 32116
rect 29204 32060 29214 32116
rect 46386 32060 46396 32116
rect 46452 32060 54236 32116
rect 54292 32060 54302 32116
rect 3332 31948 5180 32004
rect 5236 31948 5246 32004
rect 11106 31948 11116 32004
rect 11172 31948 11900 32004
rect 11956 31948 11966 32004
rect 12114 31948 12124 32004
rect 12180 31948 12190 32004
rect 32946 31948 32956 32004
rect 33012 31948 33852 32004
rect 33908 31948 33918 32004
rect 40572 31948 49756 32004
rect 49812 31948 49822 32004
rect 53890 31948 53900 32004
rect 53956 31948 54684 32004
rect 54740 31948 55020 32004
rect 55076 31948 55356 32004
rect 55412 31948 55422 32004
rect 3332 31892 3388 31948
rect 12124 31892 12180 31948
rect 3042 31836 3052 31892
rect 3108 31836 3388 31892
rect 8754 31836 8764 31892
rect 8820 31836 9996 31892
rect 10052 31836 10220 31892
rect 10276 31836 10668 31892
rect 10724 31836 10734 31892
rect 11666 31836 11676 31892
rect 11732 31836 13860 31892
rect 14242 31836 14252 31892
rect 14308 31836 14924 31892
rect 14980 31836 15148 31892
rect 20262 31836 20300 31892
rect 20356 31836 20366 31892
rect 21970 31836 21980 31892
rect 22036 31836 22540 31892
rect 22596 31836 22606 31892
rect 25890 31836 25900 31892
rect 25956 31836 28140 31892
rect 28196 31836 28206 31892
rect 28578 31836 28588 31892
rect 28644 31836 29260 31892
rect 29316 31836 29484 31892
rect 29540 31836 29550 31892
rect 36418 31836 36428 31892
rect 36484 31836 40348 31892
rect 40404 31836 40414 31892
rect 13804 31780 13860 31836
rect 15092 31780 15148 31836
rect 10098 31724 10108 31780
rect 10164 31724 13580 31780
rect 13636 31724 13646 31780
rect 13804 31724 14476 31780
rect 14532 31724 14542 31780
rect 15092 31724 16940 31780
rect 16996 31724 17006 31780
rect 19842 31724 19852 31780
rect 19908 31724 22428 31780
rect 22484 31724 23660 31780
rect 23716 31724 23726 31780
rect 26852 31724 33628 31780
rect 33684 31724 33694 31780
rect 26852 31668 26908 31724
rect 2706 31612 2716 31668
rect 2772 31612 3612 31668
rect 3668 31612 3678 31668
rect 4946 31612 4956 31668
rect 5012 31612 5964 31668
rect 6020 31612 6030 31668
rect 7410 31612 7420 31668
rect 7476 31612 9884 31668
rect 9940 31612 10556 31668
rect 10612 31612 10622 31668
rect 12338 31612 12348 31668
rect 12404 31612 14140 31668
rect 14196 31612 14206 31668
rect 15922 31612 15932 31668
rect 15988 31612 26908 31668
rect 27010 31612 27020 31668
rect 27076 31612 27692 31668
rect 27748 31612 27758 31668
rect 30258 31612 30268 31668
rect 30324 31612 38444 31668
rect 38500 31612 38668 31668
rect 38724 31612 38734 31668
rect 40572 31556 40628 31948
rect 53554 31836 53564 31892
rect 53620 31836 56700 31892
rect 56756 31836 56766 31892
rect 51538 31724 51548 31780
rect 51604 31724 52444 31780
rect 52500 31724 52510 31780
rect 8754 31500 8764 31556
rect 8820 31500 9772 31556
rect 9828 31500 10780 31556
rect 10836 31500 10846 31556
rect 11442 31500 11452 31556
rect 11508 31500 13020 31556
rect 13076 31500 13086 31556
rect 22866 31500 22876 31556
rect 22932 31500 24108 31556
rect 24164 31500 24174 31556
rect 27570 31500 27580 31556
rect 27636 31500 28364 31556
rect 28420 31500 28430 31556
rect 40114 31500 40124 31556
rect 40180 31500 40628 31556
rect 43586 31500 43596 31556
rect 43652 31500 46396 31556
rect 46452 31500 46462 31556
rect 47506 31500 47516 31556
rect 47572 31500 47852 31556
rect 47908 31500 48636 31556
rect 48692 31500 49084 31556
rect 49140 31500 50204 31556
rect 50260 31500 50270 31556
rect 56354 31500 56364 31556
rect 56420 31500 57148 31556
rect 57204 31500 57708 31556
rect 57764 31500 57774 31556
rect 4946 31388 4956 31444
rect 5012 31388 6636 31444
rect 6692 31388 7868 31444
rect 7924 31388 8540 31444
rect 8596 31388 9548 31444
rect 9604 31388 9614 31444
rect 12236 31388 19516 31444
rect 19572 31388 19582 31444
rect 22540 31388 40572 31444
rect 40628 31388 41468 31444
rect 41524 31388 41534 31444
rect 12236 31332 12292 31388
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 22540 31332 22596 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 1922 31276 1932 31332
rect 1988 31276 2268 31332
rect 2324 31276 8092 31332
rect 8148 31276 8158 31332
rect 8642 31276 8652 31332
rect 8708 31276 12292 31332
rect 13010 31276 13020 31332
rect 13076 31276 16884 31332
rect 22530 31276 22540 31332
rect 22596 31276 22606 31332
rect 36754 31276 36764 31332
rect 36820 31276 37884 31332
rect 37940 31276 37950 31332
rect 38612 31276 42252 31332
rect 42308 31276 42318 31332
rect 16828 31220 16884 31276
rect 2034 31164 2044 31220
rect 2100 31164 2828 31220
rect 2884 31164 3164 31220
rect 3220 31164 3230 31220
rect 14130 31164 14140 31220
rect 14196 31164 14812 31220
rect 14868 31164 15484 31220
rect 15540 31164 15550 31220
rect 16828 31164 22316 31220
rect 22372 31164 22382 31220
rect 22530 31164 22540 31220
rect 22596 31164 22652 31220
rect 22708 31164 23772 31220
rect 23828 31164 23838 31220
rect 32162 31164 32172 31220
rect 32228 31164 33180 31220
rect 33236 31164 33246 31220
rect 2370 31052 2380 31108
rect 2436 31052 2940 31108
rect 2996 31052 3006 31108
rect 14578 31052 14588 31108
rect 14644 31052 15260 31108
rect 15316 31052 15326 31108
rect 30482 31052 30492 31108
rect 30548 31052 31724 31108
rect 31780 31052 32060 31108
rect 32116 31052 32126 31108
rect 36194 31052 36204 31108
rect 36260 31052 37436 31108
rect 37492 31052 37502 31108
rect 38612 30996 38668 31276
rect 46050 31164 46060 31220
rect 46116 31164 50652 31220
rect 50708 31164 50718 31220
rect 49494 31052 49532 31108
rect 49588 31052 49598 31108
rect 2482 30940 2492 30996
rect 2548 30940 2884 30996
rect 5058 30940 5068 30996
rect 5124 30940 5516 30996
rect 5572 30940 5582 30996
rect 9090 30940 9100 30996
rect 9156 30940 10332 30996
rect 10388 30940 10556 30996
rect 10612 30940 10622 30996
rect 13570 30940 13580 30996
rect 13636 30940 14028 30996
rect 14084 30940 16380 30996
rect 16436 30940 16446 30996
rect 26852 30940 38668 30996
rect 44482 30940 44492 30996
rect 44548 30940 45724 30996
rect 45780 30940 46060 30996
rect 46116 30940 46126 30996
rect 46498 30940 46508 30996
rect 46564 30940 48076 30996
rect 48132 30940 48142 30996
rect 50306 30940 50316 30996
rect 50372 30940 50428 30996
rect 50484 30940 50494 30996
rect 2828 30884 2884 30940
rect 2818 30828 2828 30884
rect 2884 30828 2894 30884
rect 6738 30828 6748 30884
rect 6804 30828 7644 30884
rect 7700 30828 11116 30884
rect 11172 30828 12012 30884
rect 12068 30828 12078 30884
rect 15026 30828 15036 30884
rect 15092 30828 15260 30884
rect 15316 30828 16044 30884
rect 16100 30828 20524 30884
rect 20580 30828 20590 30884
rect 9986 30716 9996 30772
rect 10052 30716 10668 30772
rect 10724 30716 10734 30772
rect 21970 30716 21980 30772
rect 22036 30716 24556 30772
rect 24612 30716 24622 30772
rect 26852 30660 26908 30940
rect 27458 30828 27468 30884
rect 27524 30828 31612 30884
rect 31668 30828 31678 30884
rect 33170 30828 33180 30884
rect 33236 30828 40460 30884
rect 40516 30828 40526 30884
rect 42242 30828 42252 30884
rect 42308 30828 45388 30884
rect 45444 30828 46844 30884
rect 46900 30828 47180 30884
rect 47236 30828 47246 30884
rect 52098 30828 52108 30884
rect 52164 30828 52892 30884
rect 52948 30828 53340 30884
rect 53396 30828 53788 30884
rect 53844 30828 53854 30884
rect 55234 30828 55244 30884
rect 55300 30828 55692 30884
rect 55748 30828 57820 30884
rect 57876 30828 58268 30884
rect 58324 30828 58334 30884
rect 43810 30716 43820 30772
rect 43876 30716 52332 30772
rect 52388 30716 52398 30772
rect 9202 30604 9212 30660
rect 9268 30604 26908 30660
rect 40898 30604 40908 30660
rect 40964 30604 56700 30660
rect 56756 30604 57036 30660
rect 57092 30604 57102 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 12786 30492 12796 30548
rect 12852 30492 32060 30548
rect 32116 30492 32126 30548
rect 50642 30492 50652 30548
rect 50708 30492 51436 30548
rect 51492 30492 51502 30548
rect 14690 30380 14700 30436
rect 14756 30380 15148 30436
rect 15204 30380 15214 30436
rect 16930 30380 16940 30436
rect 16996 30380 17724 30436
rect 17780 30380 18284 30436
rect 18340 30380 19180 30436
rect 19236 30380 19246 30436
rect 37650 30380 37660 30436
rect 37716 30380 38108 30436
rect 38164 30380 38174 30436
rect 46162 30380 46172 30436
rect 46228 30380 54572 30436
rect 54628 30380 54638 30436
rect 15670 30268 15708 30324
rect 15764 30268 16828 30324
rect 16884 30268 16894 30324
rect 20514 30268 20524 30324
rect 20580 30268 21980 30324
rect 22036 30268 22764 30324
rect 22820 30268 22830 30324
rect 31938 30268 31948 30324
rect 32004 30268 33740 30324
rect 33796 30268 33806 30324
rect 35298 30268 35308 30324
rect 35364 30268 36204 30324
rect 36260 30268 36270 30324
rect 38668 30268 51436 30324
rect 51492 30268 51502 30324
rect 53106 30268 53116 30324
rect 53172 30268 53788 30324
rect 53844 30268 54236 30324
rect 54292 30268 54460 30324
rect 54516 30268 55356 30324
rect 55412 30268 55422 30324
rect 1922 30156 1932 30212
rect 1988 30156 3724 30212
rect 3780 30156 3790 30212
rect 4162 30156 4172 30212
rect 4228 30156 7308 30212
rect 7364 30156 8316 30212
rect 8372 30156 10892 30212
rect 10948 30156 11452 30212
rect 11508 30156 11900 30212
rect 11956 30156 11966 30212
rect 14914 30156 14924 30212
rect 14980 30156 15596 30212
rect 15652 30156 15662 30212
rect 16370 30156 16380 30212
rect 16436 30156 16940 30212
rect 16996 30156 18396 30212
rect 18452 30156 18462 30212
rect 38668 30100 38724 30268
rect 42354 30156 42364 30212
rect 42420 30156 43932 30212
rect 43988 30156 46620 30212
rect 46676 30156 46686 30212
rect 49746 30156 49756 30212
rect 49812 30156 50988 30212
rect 51044 30156 51324 30212
rect 51380 30156 51390 30212
rect 5842 30044 5852 30100
rect 5908 30044 6412 30100
rect 6468 30044 6636 30100
rect 6692 30044 6702 30100
rect 7970 30044 7980 30100
rect 8036 30044 8652 30100
rect 8708 30044 9100 30100
rect 9156 30044 9166 30100
rect 9426 30044 9436 30100
rect 9492 30044 11564 30100
rect 11620 30044 12908 30100
rect 12964 30044 12974 30100
rect 29698 30044 29708 30100
rect 29764 30044 30268 30100
rect 30324 30044 30334 30100
rect 30706 30044 30716 30100
rect 30772 30044 38724 30100
rect 41682 30044 41692 30100
rect 41748 30044 42476 30100
rect 42532 30044 43820 30100
rect 43876 30044 43886 30100
rect 44146 30044 44156 30100
rect 44212 30044 45388 30100
rect 45444 30044 49308 30100
rect 49364 30044 49374 30100
rect 49634 30044 49644 30100
rect 49700 30044 50204 30100
rect 50260 30044 50270 30100
rect 2706 29932 2716 29988
rect 2772 29932 3276 29988
rect 3332 29932 5068 29988
rect 5124 29932 5134 29988
rect 9650 29932 9660 29988
rect 9716 29932 10556 29988
rect 10612 29932 11116 29988
rect 11172 29932 12348 29988
rect 12404 29932 12414 29988
rect 18386 29932 18396 29988
rect 18452 29932 22428 29988
rect 22484 29932 22652 29988
rect 22708 29932 22876 29988
rect 22932 29932 23324 29988
rect 23380 29932 23390 29988
rect 24882 29932 24892 29988
rect 24948 29932 26236 29988
rect 26292 29932 26572 29988
rect 26628 29932 27356 29988
rect 27412 29932 27422 29988
rect 29026 29932 29036 29988
rect 29092 29932 31276 29988
rect 31332 29932 31836 29988
rect 31892 29932 31902 29988
rect 7522 29820 7532 29876
rect 7588 29820 8204 29876
rect 8260 29820 17948 29876
rect 18004 29820 18014 29876
rect 22306 29820 22316 29876
rect 22372 29820 24220 29876
rect 24276 29820 24286 29876
rect 27234 29820 27244 29876
rect 27300 29820 34524 29876
rect 34580 29820 35084 29876
rect 35140 29820 35980 29876
rect 36036 29820 36652 29876
rect 36708 29820 36718 29876
rect 38612 29820 38724 30044
rect 46246 29932 46284 29988
rect 46340 29932 46350 29988
rect 47618 29932 47628 29988
rect 47684 29932 48524 29988
rect 48580 29932 50876 29988
rect 50932 29932 54908 29988
rect 54964 29932 55468 29988
rect 55524 29932 55534 29988
rect 51202 29820 51212 29876
rect 51268 29820 51772 29876
rect 51828 29820 51838 29876
rect 54562 29820 54572 29876
rect 54628 29820 55244 29876
rect 55300 29820 55310 29876
rect 56354 29820 56364 29876
rect 56420 29820 56924 29876
rect 56980 29820 56990 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 4274 29708 4284 29764
rect 4340 29708 5628 29764
rect 5684 29708 15820 29764
rect 15876 29708 15886 29764
rect 21074 29708 21084 29764
rect 21140 29708 21532 29764
rect 21588 29708 22428 29764
rect 22484 29708 22494 29764
rect 29586 29708 29596 29764
rect 29652 29708 30828 29764
rect 30884 29708 35532 29764
rect 35588 29708 35598 29764
rect 36418 29708 36428 29764
rect 36484 29708 37436 29764
rect 37492 29708 42028 29764
rect 42084 29708 42094 29764
rect 43698 29708 43708 29764
rect 43764 29708 44044 29764
rect 44100 29708 44716 29764
rect 44772 29708 49924 29764
rect 43708 29652 43764 29708
rect 49868 29652 49924 29708
rect 1698 29596 1708 29652
rect 1764 29596 3276 29652
rect 3332 29596 3612 29652
rect 3668 29596 3678 29652
rect 4834 29596 4844 29652
rect 4900 29596 7196 29652
rect 7252 29596 7262 29652
rect 7634 29596 7644 29652
rect 7700 29596 9548 29652
rect 9604 29596 9614 29652
rect 18946 29596 18956 29652
rect 19012 29596 19964 29652
rect 20020 29596 27132 29652
rect 27188 29596 27198 29652
rect 27346 29596 27356 29652
rect 27412 29596 28476 29652
rect 28532 29596 28542 29652
rect 30034 29596 30044 29652
rect 30100 29596 30716 29652
rect 30772 29596 30782 29652
rect 41346 29596 41356 29652
rect 41412 29596 41916 29652
rect 41972 29596 42364 29652
rect 42420 29596 42430 29652
rect 43250 29596 43260 29652
rect 43316 29596 43764 29652
rect 44370 29596 44380 29652
rect 44436 29596 45948 29652
rect 46004 29596 46508 29652
rect 46564 29596 47404 29652
rect 47460 29596 47470 29652
rect 48738 29596 48748 29652
rect 48804 29596 49644 29652
rect 49700 29596 49710 29652
rect 49868 29596 50428 29652
rect 50484 29596 51044 29652
rect 51202 29596 51212 29652
rect 51268 29596 53452 29652
rect 53508 29596 53518 29652
rect 50988 29540 51044 29596
rect 5170 29484 5180 29540
rect 5236 29484 6076 29540
rect 6132 29484 6142 29540
rect 9090 29484 9100 29540
rect 9156 29484 9660 29540
rect 9716 29484 9726 29540
rect 14018 29484 14028 29540
rect 14084 29484 16268 29540
rect 16324 29484 16334 29540
rect 19618 29484 19628 29540
rect 19684 29484 20412 29540
rect 20468 29484 21420 29540
rect 21476 29484 25564 29540
rect 25620 29484 26460 29540
rect 26516 29484 28812 29540
rect 28868 29484 28878 29540
rect 36530 29484 36540 29540
rect 36596 29484 37884 29540
rect 37940 29484 38332 29540
rect 38388 29484 38398 29540
rect 38658 29484 38668 29540
rect 38724 29484 39116 29540
rect 39172 29484 40684 29540
rect 40740 29484 41580 29540
rect 41636 29484 41646 29540
rect 44818 29484 44828 29540
rect 44884 29484 47292 29540
rect 47348 29484 47358 29540
rect 50194 29484 50204 29540
rect 50260 29484 50932 29540
rect 50988 29484 51100 29540
rect 51156 29484 51884 29540
rect 51940 29484 51950 29540
rect 54338 29484 54348 29540
rect 54404 29484 55580 29540
rect 55636 29484 56588 29540
rect 56644 29484 57372 29540
rect 57428 29484 57438 29540
rect 1586 29372 1596 29428
rect 1652 29372 3724 29428
rect 3780 29372 3790 29428
rect 10434 29372 10444 29428
rect 10500 29372 11452 29428
rect 11508 29372 12460 29428
rect 12516 29372 12526 29428
rect 14802 29372 14812 29428
rect 14868 29372 15596 29428
rect 15652 29372 15662 29428
rect 27906 29372 27916 29428
rect 27972 29372 32844 29428
rect 32900 29372 33516 29428
rect 33572 29372 33964 29428
rect 34020 29372 34030 29428
rect 35410 29372 35420 29428
rect 35476 29372 36428 29428
rect 36484 29372 36494 29428
rect 36642 29372 36652 29428
rect 36708 29372 37324 29428
rect 37380 29372 37772 29428
rect 37828 29372 37838 29428
rect 38668 29316 38724 29484
rect 45836 29316 45892 29484
rect 50876 29428 50932 29484
rect 46610 29372 46620 29428
rect 46676 29372 47964 29428
rect 48020 29372 50316 29428
rect 50372 29372 50382 29428
rect 50876 29372 52556 29428
rect 52612 29372 52622 29428
rect 52770 29372 52780 29428
rect 52836 29372 53564 29428
rect 53620 29372 54908 29428
rect 54964 29372 54974 29428
rect 2034 29260 2044 29316
rect 2100 29260 2156 29316
rect 2212 29260 2222 29316
rect 11666 29260 11676 29316
rect 11732 29260 14924 29316
rect 14980 29260 14990 29316
rect 33516 29260 38724 29316
rect 45826 29260 45836 29316
rect 45892 29260 45902 29316
rect 46050 29260 46060 29316
rect 46116 29260 47180 29316
rect 47236 29260 48188 29316
rect 48244 29260 48972 29316
rect 49028 29260 51548 29316
rect 51604 29260 51614 29316
rect 51762 29260 51772 29316
rect 51828 29260 52668 29316
rect 52724 29260 53004 29316
rect 53060 29260 56364 29316
rect 56420 29260 56430 29316
rect 12338 29148 12348 29204
rect 12404 29148 22316 29204
rect 22372 29148 22382 29204
rect 23314 29148 23324 29204
rect 23380 29148 23996 29204
rect 24052 29148 29820 29204
rect 29876 29148 30492 29204
rect 30548 29148 30558 29204
rect 33516 29092 33572 29260
rect 38210 29148 38220 29204
rect 38276 29148 47068 29204
rect 47124 29148 47134 29204
rect 49746 29148 49756 29204
rect 49812 29148 50428 29204
rect 50484 29148 50494 29204
rect 51426 29148 51436 29204
rect 51492 29148 52108 29204
rect 52164 29148 52174 29204
rect 17154 29036 17164 29092
rect 17220 29036 17612 29092
rect 17668 29036 29596 29092
rect 29652 29036 29662 29092
rect 33506 29036 33516 29092
rect 33572 29036 33582 29092
rect 51314 29036 51324 29092
rect 51380 29036 51996 29092
rect 52052 29036 52062 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 59200 28980 59800 29008
rect 13346 28924 13356 28980
rect 13412 28924 14700 28980
rect 14756 28924 16044 28980
rect 16100 28924 23548 28980
rect 23604 28924 26460 28980
rect 26516 28924 27020 28980
rect 27076 28924 27086 28980
rect 30258 28924 30268 28980
rect 30324 28924 30828 28980
rect 30884 28924 30894 28980
rect 45938 28924 45948 28980
rect 46004 28924 46956 28980
rect 47012 28924 47022 28980
rect 56018 28924 56028 28980
rect 56084 28924 59800 28980
rect 59200 28896 59800 28924
rect 12450 28812 12460 28868
rect 12516 28812 31276 28868
rect 31332 28812 31342 28868
rect 34626 28812 34636 28868
rect 34692 28812 35756 28868
rect 35812 28812 38668 28868
rect 40898 28812 40908 28868
rect 40964 28812 41580 28868
rect 41636 28812 41748 28868
rect 42690 28812 42700 28868
rect 42756 28812 46620 28868
rect 46676 28812 46686 28868
rect 47730 28812 47740 28868
rect 47796 28812 48524 28868
rect 48580 28812 51212 28868
rect 51268 28812 51278 28868
rect 38612 28756 38668 28812
rect 41692 28756 41748 28812
rect 2594 28700 2604 28756
rect 2660 28700 5180 28756
rect 5236 28700 5246 28756
rect 22418 28700 22428 28756
rect 22484 28700 23996 28756
rect 24052 28700 24332 28756
rect 24388 28700 25900 28756
rect 25956 28700 25966 28756
rect 30594 28700 30604 28756
rect 30660 28700 31724 28756
rect 31780 28700 31790 28756
rect 35074 28700 35084 28756
rect 35140 28700 35868 28756
rect 35924 28700 36092 28756
rect 36148 28700 36158 28756
rect 38612 28700 38780 28756
rect 38836 28700 38846 28756
rect 40338 28700 40348 28756
rect 40404 28700 41468 28756
rect 41524 28700 41534 28756
rect 41692 28700 48412 28756
rect 48468 28700 49756 28756
rect 49812 28700 49822 28756
rect 50418 28700 50428 28756
rect 50484 28700 56140 28756
rect 56196 28700 56206 28756
rect 2156 28588 3276 28644
rect 3332 28588 3948 28644
rect 4004 28588 4508 28644
rect 4564 28588 4574 28644
rect 14466 28588 14476 28644
rect 14532 28588 15372 28644
rect 15428 28588 15438 28644
rect 17612 28588 18508 28644
rect 18564 28588 18574 28644
rect 30034 28588 30044 28644
rect 30100 28588 30660 28644
rect 30930 28588 30940 28644
rect 30996 28588 32284 28644
rect 32340 28588 32732 28644
rect 32788 28588 33404 28644
rect 33460 28588 33470 28644
rect 35634 28588 35644 28644
rect 35700 28588 37548 28644
rect 37604 28588 38220 28644
rect 38276 28588 38286 28644
rect 40786 28588 40796 28644
rect 40852 28588 41356 28644
rect 41412 28588 41422 28644
rect 43652 28588 46172 28644
rect 46228 28588 46238 28644
rect 51874 28588 51884 28644
rect 51940 28588 52108 28644
rect 52164 28588 54684 28644
rect 54740 28588 54750 28644
rect 55010 28588 55020 28644
rect 55076 28588 56700 28644
rect 56756 28588 57596 28644
rect 57652 28588 58044 28644
rect 58100 28588 58110 28644
rect 2156 28420 2212 28588
rect 17612 28532 17668 28588
rect 30604 28532 30660 28588
rect 43652 28532 43708 28588
rect 2930 28476 2940 28532
rect 2996 28476 3388 28532
rect 13682 28476 13692 28532
rect 13748 28476 17052 28532
rect 17108 28476 17118 28532
rect 17602 28476 17612 28532
rect 17668 28476 17678 28532
rect 30594 28476 30604 28532
rect 30660 28476 30670 28532
rect 32162 28476 32172 28532
rect 32228 28476 35084 28532
rect 35140 28476 35150 28532
rect 43474 28476 43484 28532
rect 43540 28476 43708 28532
rect 48178 28476 48188 28532
rect 48244 28476 49308 28532
rect 49364 28476 49374 28532
rect 50642 28476 50652 28532
rect 50708 28476 51660 28532
rect 51716 28476 52220 28532
rect 52276 28476 53452 28532
rect 53508 28476 53518 28532
rect 56466 28476 56476 28532
rect 56532 28476 57260 28532
rect 57316 28476 57326 28532
rect 3332 28420 3388 28476
rect 2146 28364 2156 28420
rect 2212 28364 2222 28420
rect 3332 28364 21868 28420
rect 21924 28364 21934 28420
rect 32050 28364 32060 28420
rect 32116 28364 32508 28420
rect 32564 28364 33628 28420
rect 33684 28364 33694 28420
rect 34962 28364 34972 28420
rect 35028 28364 37436 28420
rect 37492 28364 37502 28420
rect 42578 28364 42588 28420
rect 42644 28364 42924 28420
rect 42980 28364 43820 28420
rect 43876 28364 43886 28420
rect 54002 28364 54012 28420
rect 54068 28364 56588 28420
rect 56644 28364 57820 28420
rect 57876 28364 57886 28420
rect 9650 28252 9660 28308
rect 9716 28252 17612 28308
rect 17668 28252 17678 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 1250 28140 1260 28196
rect 1316 28140 16940 28196
rect 16996 28140 17948 28196
rect 18004 28140 18014 28196
rect 37762 28140 37772 28196
rect 37828 28140 49644 28196
rect 49700 28140 49710 28196
rect 49644 28084 49700 28140
rect 2370 28028 2380 28084
rect 2436 28028 3052 28084
rect 3108 28028 3500 28084
rect 3556 28028 5516 28084
rect 5572 28028 10332 28084
rect 10388 28028 10398 28084
rect 14242 28028 14252 28084
rect 14308 28028 15484 28084
rect 15540 28028 15550 28084
rect 25106 28028 25116 28084
rect 25172 28028 25676 28084
rect 25732 28028 25742 28084
rect 47058 28028 47068 28084
rect 47124 28028 48636 28084
rect 48692 28028 48702 28084
rect 49644 28028 50876 28084
rect 50932 28028 50942 28084
rect 51202 28028 51212 28084
rect 51268 28028 51772 28084
rect 51828 28028 53900 28084
rect 53956 28028 53966 28084
rect 15092 27916 16268 27972
rect 16324 27916 16334 27972
rect 28130 27916 28140 27972
rect 28196 27916 30268 27972
rect 30324 27916 30334 27972
rect 33730 27916 33740 27972
rect 33796 27916 34076 27972
rect 34132 27916 38444 27972
rect 38500 27916 38510 27972
rect 38612 27916 41580 27972
rect 41636 27916 41646 27972
rect 43026 27916 43036 27972
rect 43092 27916 43372 27972
rect 43428 27916 44492 27972
rect 44548 27916 44558 27972
rect 44706 27916 44716 27972
rect 44772 27916 45612 27972
rect 45668 27916 47964 27972
rect 48020 27916 48030 27972
rect 48850 27916 48860 27972
rect 48916 27916 53676 27972
rect 53732 27916 53742 27972
rect 54562 27916 54572 27972
rect 54628 27916 55468 27972
rect 55524 27916 57372 27972
rect 57428 27916 57438 27972
rect 15092 27860 15148 27916
rect 38612 27860 38668 27916
rect 11330 27804 11340 27860
rect 11396 27804 14588 27860
rect 14644 27804 15148 27860
rect 18274 27804 18284 27860
rect 18340 27804 18844 27860
rect 18900 27804 18910 27860
rect 27682 27804 27692 27860
rect 27748 27804 29372 27860
rect 29428 27804 29438 27860
rect 35970 27804 35980 27860
rect 36036 27804 38668 27860
rect 40002 27804 40012 27860
rect 40068 27804 41132 27860
rect 41188 27804 41198 27860
rect 41906 27804 41916 27860
rect 41972 27804 43148 27860
rect 43204 27804 43214 27860
rect 46946 27804 46956 27860
rect 47012 27804 47628 27860
rect 47684 27804 48300 27860
rect 48356 27804 48524 27860
rect 48580 27804 48590 27860
rect 48860 27804 56364 27860
rect 56420 27804 56430 27860
rect 33954 27692 33964 27748
rect 34020 27692 35196 27748
rect 35252 27692 36540 27748
rect 36596 27692 36606 27748
rect 42690 27692 42700 27748
rect 42756 27692 42924 27748
rect 42980 27692 42990 27748
rect 43810 27692 43820 27748
rect 43876 27692 46844 27748
rect 46900 27692 47180 27748
rect 47236 27692 48636 27748
rect 48692 27692 48702 27748
rect 200 27636 800 27664
rect 48860 27636 48916 27804
rect 49522 27692 49532 27748
rect 49588 27692 52332 27748
rect 52388 27692 52398 27748
rect 53004 27692 53452 27748
rect 53508 27692 54236 27748
rect 54292 27692 57820 27748
rect 57876 27692 57886 27748
rect 53004 27636 53060 27692
rect 200 27580 1932 27636
rect 1988 27580 1998 27636
rect 17938 27580 17948 27636
rect 18004 27580 19180 27636
rect 19236 27580 21644 27636
rect 21700 27580 21710 27636
rect 24770 27580 24780 27636
rect 24836 27580 26012 27636
rect 26068 27580 26078 27636
rect 34066 27580 34076 27636
rect 34132 27580 34748 27636
rect 34804 27580 35756 27636
rect 35812 27580 35822 27636
rect 37538 27580 37548 27636
rect 37604 27580 37772 27636
rect 37828 27580 37838 27636
rect 42802 27580 42812 27636
rect 42868 27580 43596 27636
rect 43652 27580 43662 27636
rect 46946 27580 46956 27636
rect 47012 27580 47068 27636
rect 47124 27580 47628 27636
rect 47684 27580 47694 27636
rect 48626 27580 48636 27636
rect 48692 27580 48916 27636
rect 50306 27580 50316 27636
rect 50372 27580 53004 27636
rect 53060 27580 53070 27636
rect 53890 27580 53900 27636
rect 53956 27580 55804 27636
rect 55860 27580 55870 27636
rect 200 27552 800 27580
rect 8194 27468 8204 27524
rect 8260 27468 31948 27524
rect 32004 27468 32014 27524
rect 36754 27468 36764 27524
rect 36820 27468 42924 27524
rect 42980 27468 42990 27524
rect 44482 27468 44492 27524
rect 44548 27468 45612 27524
rect 45668 27468 46620 27524
rect 46676 27468 47516 27524
rect 47572 27468 54236 27524
rect 54292 27468 54302 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 11330 27356 11340 27412
rect 11396 27356 13468 27412
rect 13524 27356 13534 27412
rect 15138 27356 15148 27412
rect 15204 27356 15820 27412
rect 15876 27356 30380 27412
rect 30436 27356 31164 27412
rect 31220 27356 31230 27412
rect 37090 27356 37100 27412
rect 37156 27356 37884 27412
rect 37940 27356 38668 27412
rect 41906 27356 41916 27412
rect 41972 27356 42588 27412
rect 42644 27356 42654 27412
rect 43586 27356 43596 27412
rect 43652 27356 48412 27412
rect 48468 27356 48636 27412
rect 48692 27356 48702 27412
rect 49298 27356 49308 27412
rect 49364 27356 49644 27412
rect 49700 27356 54684 27412
rect 54740 27356 54750 27412
rect 38612 27300 38668 27356
rect 3042 27244 3052 27300
rect 3108 27244 29204 27300
rect 29362 27244 29372 27300
rect 29428 27244 30492 27300
rect 30548 27244 31388 27300
rect 31444 27244 31454 27300
rect 35746 27244 35756 27300
rect 35812 27244 38444 27300
rect 38500 27244 38510 27300
rect 38612 27244 38892 27300
rect 38948 27244 38958 27300
rect 50866 27244 50876 27300
rect 50932 27244 56252 27300
rect 56308 27244 56318 27300
rect 17714 27132 17724 27188
rect 17780 27132 18508 27188
rect 18564 27132 18574 27188
rect 27570 27132 27580 27188
rect 27636 27132 28252 27188
rect 28308 27132 28588 27188
rect 28644 27132 28654 27188
rect 29148 27076 29204 27244
rect 31154 27132 31164 27188
rect 31220 27132 35644 27188
rect 35700 27132 35980 27188
rect 36036 27132 36046 27188
rect 38210 27132 38220 27188
rect 38276 27132 39676 27188
rect 39732 27132 43820 27188
rect 43876 27132 43886 27188
rect 48178 27132 48188 27188
rect 48244 27132 51884 27188
rect 51940 27132 51950 27188
rect 26674 27020 26684 27076
rect 26740 27020 27468 27076
rect 27524 27020 27534 27076
rect 28018 27020 28028 27076
rect 28084 27020 28094 27076
rect 29148 27020 33292 27076
rect 33348 27020 33358 27076
rect 34850 27020 34860 27076
rect 34916 27020 37996 27076
rect 38052 27020 38062 27076
rect 38434 27020 38444 27076
rect 38500 27020 40572 27076
rect 40628 27020 40638 27076
rect 41122 27020 41132 27076
rect 41188 27020 41580 27076
rect 41636 27020 41646 27076
rect 47954 27020 47964 27076
rect 48020 27020 49084 27076
rect 49140 27020 51212 27076
rect 51268 27020 51278 27076
rect 52658 27020 52668 27076
rect 52724 27020 53228 27076
rect 53284 27020 53788 27076
rect 53844 27020 54348 27076
rect 54404 27020 54414 27076
rect 28028 26964 28084 27020
rect 13010 26908 13020 26964
rect 13076 26908 13804 26964
rect 13860 26908 13870 26964
rect 16258 26908 16268 26964
rect 16324 26908 17164 26964
rect 17220 26908 18060 26964
rect 18116 26908 20300 26964
rect 20356 26908 20366 26964
rect 20514 26908 20524 26964
rect 20580 26908 21980 26964
rect 22036 26908 23772 26964
rect 23828 26908 24556 26964
rect 24612 26908 24622 26964
rect 26338 26908 26348 26964
rect 26404 26908 27244 26964
rect 27300 26908 28084 26964
rect 30604 26908 30828 26964
rect 30884 26908 30894 26964
rect 34626 26908 34636 26964
rect 34692 26908 34972 26964
rect 35028 26908 36988 26964
rect 37044 26908 37492 26964
rect 37650 26908 37660 26964
rect 37716 26908 38108 26964
rect 38164 26908 38668 26964
rect 38724 26908 38734 26964
rect 41346 26908 41356 26964
rect 41412 26908 42364 26964
rect 42420 26908 42430 26964
rect 42588 26908 42924 26964
rect 42980 26908 42990 26964
rect 43250 26908 43260 26964
rect 43316 26908 44492 26964
rect 44548 26908 45276 26964
rect 45332 26908 45342 26964
rect 46386 26908 46396 26964
rect 46452 26908 47740 26964
rect 47796 26908 48748 26964
rect 48804 26908 48814 26964
rect 49186 26908 49196 26964
rect 49252 26908 49308 26964
rect 49364 26908 49374 26964
rect 50306 26908 50316 26964
rect 50372 26908 50428 26964
rect 50484 26908 50494 26964
rect 30594 26852 30604 26908
rect 30660 26852 30670 26908
rect 37436 26852 37492 26908
rect 42588 26852 42644 26908
rect 24434 26796 24444 26852
rect 24500 26796 24892 26852
rect 24948 26796 25676 26852
rect 25732 26796 25742 26852
rect 32162 26796 32172 26852
rect 32228 26796 32844 26852
rect 32900 26796 32910 26852
rect 35634 26796 35644 26852
rect 35700 26796 36316 26852
rect 36372 26796 36382 26852
rect 37436 26796 38892 26852
rect 38948 26796 38958 26852
rect 39218 26796 39228 26852
rect 39284 26796 40124 26852
rect 40180 26796 40190 26852
rect 42578 26796 42588 26852
rect 42644 26796 42654 26852
rect 44146 26796 44156 26852
rect 44212 26796 45836 26852
rect 45892 26796 48076 26852
rect 48132 26796 48142 26852
rect 56802 26796 56812 26852
rect 56868 26796 57372 26852
rect 57428 26796 57438 26852
rect 42018 26684 42028 26740
rect 42084 26684 42364 26740
rect 42420 26684 42430 26740
rect 44482 26684 44492 26740
rect 44548 26684 46508 26740
rect 46564 26684 46574 26740
rect 48850 26684 48860 26740
rect 48916 26684 49196 26740
rect 49252 26684 49262 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 24994 26572 25004 26628
rect 25060 26572 25564 26628
rect 25620 26572 25630 26628
rect 34514 26572 34524 26628
rect 34580 26572 36932 26628
rect 53554 26572 53564 26628
rect 53620 26572 55356 26628
rect 55412 26572 57708 26628
rect 57764 26572 57774 26628
rect 36876 26516 36932 26572
rect 7522 26460 7532 26516
rect 7588 26460 28700 26516
rect 28756 26460 28766 26516
rect 35410 26460 35420 26516
rect 35476 26460 35868 26516
rect 35924 26460 35934 26516
rect 36866 26460 36876 26516
rect 36932 26460 44828 26516
rect 44884 26460 49532 26516
rect 49588 26460 49598 26516
rect 53666 26460 53676 26516
rect 53732 26460 53900 26516
rect 53956 26460 53966 26516
rect 19170 26348 19180 26404
rect 19236 26348 32060 26404
rect 32116 26348 35980 26404
rect 36036 26348 36764 26404
rect 36820 26348 36830 26404
rect 37986 26348 37996 26404
rect 38052 26348 39788 26404
rect 39844 26348 39854 26404
rect 43138 26348 43148 26404
rect 43204 26348 47404 26404
rect 47460 26348 51324 26404
rect 51380 26348 51390 26404
rect 51762 26348 51772 26404
rect 51828 26348 52556 26404
rect 52612 26348 52622 26404
rect 53442 26348 53452 26404
rect 53508 26348 54012 26404
rect 54068 26348 54908 26404
rect 54964 26348 57372 26404
rect 57428 26348 57438 26404
rect 18386 26236 18396 26292
rect 18452 26236 18956 26292
rect 19012 26236 19022 26292
rect 19842 26236 19852 26292
rect 19908 26236 20412 26292
rect 20468 26236 20478 26292
rect 28466 26236 28476 26292
rect 28532 26236 29932 26292
rect 29988 26236 29998 26292
rect 32498 26236 32508 26292
rect 32564 26236 33180 26292
rect 33236 26236 33246 26292
rect 35634 26236 35644 26292
rect 35700 26236 38220 26292
rect 38276 26236 39340 26292
rect 39396 26236 43820 26292
rect 43876 26236 47068 26292
rect 47124 26236 52668 26292
rect 52724 26236 52734 26292
rect 56242 26236 56252 26292
rect 56308 26236 56812 26292
rect 56868 26236 56878 26292
rect 19618 26124 19628 26180
rect 19684 26124 20860 26180
rect 20916 26124 21756 26180
rect 21812 26124 21822 26180
rect 33506 26124 33516 26180
rect 33572 26124 35420 26180
rect 35476 26124 35486 26180
rect 40562 26124 40572 26180
rect 40628 26124 41356 26180
rect 41412 26124 41468 26180
rect 41524 26124 42140 26180
rect 42196 26124 42206 26180
rect 45826 26124 45836 26180
rect 45892 26124 48748 26180
rect 48804 26124 49868 26180
rect 49924 26124 50204 26180
rect 50260 26124 50270 26180
rect 50978 26124 50988 26180
rect 51044 26124 53452 26180
rect 53508 26124 53518 26180
rect 18162 26012 18172 26068
rect 18228 26012 31276 26068
rect 31332 26012 31342 26068
rect 35522 26012 35532 26068
rect 35588 26012 36428 26068
rect 36484 26012 36494 26068
rect 37762 26012 37772 26068
rect 37828 26012 38444 26068
rect 38500 26012 39116 26068
rect 39172 26012 39182 26068
rect 44146 26012 44156 26068
rect 44212 26012 44268 26068
rect 44324 26012 44334 26068
rect 46162 26012 46172 26068
rect 46228 26012 46844 26068
rect 46900 26012 48300 26068
rect 48356 26012 49420 26068
rect 49476 26012 49486 26068
rect 51762 26012 51772 26068
rect 51828 26012 52332 26068
rect 52388 26012 53676 26068
rect 53732 26012 53742 26068
rect 46172 25956 46228 26012
rect 6178 25900 6188 25956
rect 6244 25900 28364 25956
rect 28420 25900 28430 25956
rect 37090 25900 37100 25956
rect 37156 25900 38668 25956
rect 38882 25900 38892 25956
rect 38948 25900 40124 25956
rect 40180 25900 41804 25956
rect 41860 25900 46228 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 38612 25844 38668 25900
rect 13346 25788 13356 25844
rect 13412 25788 32284 25844
rect 32340 25788 32350 25844
rect 32722 25788 32732 25844
rect 32788 25788 33292 25844
rect 33348 25788 33358 25844
rect 36530 25788 36540 25844
rect 36596 25788 38332 25844
rect 38388 25788 38398 25844
rect 38612 25788 39004 25844
rect 39060 25788 39070 25844
rect 39218 25788 39228 25844
rect 39284 25788 41132 25844
rect 41188 25788 41198 25844
rect 48626 25788 48636 25844
rect 48692 25788 51324 25844
rect 51380 25788 51390 25844
rect 51538 25788 51548 25844
rect 51604 25788 52892 25844
rect 52948 25788 52958 25844
rect 11106 25676 11116 25732
rect 11172 25676 18172 25732
rect 18228 25676 18238 25732
rect 20962 25676 20972 25732
rect 21028 25676 21868 25732
rect 21924 25676 21934 25732
rect 32610 25676 32620 25732
rect 32676 25676 33852 25732
rect 33908 25676 33918 25732
rect 35074 25676 35084 25732
rect 35140 25676 35868 25732
rect 35924 25676 35934 25732
rect 36978 25676 36988 25732
rect 37044 25676 37940 25732
rect 38098 25676 38108 25732
rect 38164 25676 40348 25732
rect 40404 25676 40414 25732
rect 48738 25676 48748 25732
rect 48804 25676 52668 25732
rect 52724 25676 56028 25732
rect 56084 25676 56094 25732
rect 11442 25564 11452 25620
rect 11508 25564 32956 25620
rect 33012 25564 33022 25620
rect 35634 25564 35644 25620
rect 35700 25564 37100 25620
rect 37156 25564 37166 25620
rect 37884 25508 37940 25676
rect 38658 25564 38668 25620
rect 38724 25564 43148 25620
rect 43204 25564 43708 25620
rect 43764 25564 43774 25620
rect 48626 25564 48636 25620
rect 48692 25564 52332 25620
rect 52388 25564 55244 25620
rect 55300 25564 55310 25620
rect 31490 25452 31500 25508
rect 31556 25452 33964 25508
rect 34020 25452 34030 25508
rect 35410 25452 35420 25508
rect 35476 25452 35868 25508
rect 35924 25452 36876 25508
rect 36932 25452 37660 25508
rect 37716 25452 37726 25508
rect 37884 25452 39116 25508
rect 39172 25452 39182 25508
rect 39330 25452 39340 25508
rect 39396 25452 40684 25508
rect 40740 25452 40750 25508
rect 43250 25452 43260 25508
rect 43316 25452 44156 25508
rect 44212 25452 44716 25508
rect 44772 25452 44782 25508
rect 45490 25452 45500 25508
rect 45556 25452 45612 25508
rect 45668 25452 45678 25508
rect 47730 25452 47740 25508
rect 47796 25452 49308 25508
rect 49364 25452 49374 25508
rect 49522 25452 49532 25508
rect 49588 25452 51548 25508
rect 51604 25452 51614 25508
rect 51772 25452 55132 25508
rect 55188 25452 55198 25508
rect 55682 25452 55692 25508
rect 55748 25452 56476 25508
rect 56532 25452 56542 25508
rect 51772 25396 51828 25452
rect 31826 25340 31836 25396
rect 31892 25340 32396 25396
rect 32452 25340 32462 25396
rect 32722 25340 32732 25396
rect 32788 25340 33516 25396
rect 33572 25340 33582 25396
rect 34290 25340 34300 25396
rect 34356 25340 37884 25396
rect 37940 25340 37950 25396
rect 38322 25340 38332 25396
rect 38388 25340 40908 25396
rect 40964 25340 40974 25396
rect 41122 25340 41132 25396
rect 41188 25340 43372 25396
rect 43428 25340 43438 25396
rect 43820 25340 47404 25396
rect 47460 25340 47470 25396
rect 47618 25340 47628 25396
rect 47684 25340 48636 25396
rect 48692 25340 48702 25396
rect 48860 25340 50876 25396
rect 50932 25340 50942 25396
rect 51762 25340 51772 25396
rect 51828 25340 51838 25396
rect 52098 25340 52108 25396
rect 52164 25340 54236 25396
rect 54292 25340 54302 25396
rect 32732 25284 32788 25340
rect 20402 25228 20412 25284
rect 20468 25228 21532 25284
rect 21588 25228 21598 25284
rect 27794 25228 27804 25284
rect 27860 25228 28140 25284
rect 28196 25228 28588 25284
rect 28644 25228 32788 25284
rect 35186 25228 35196 25284
rect 35252 25228 36316 25284
rect 36372 25228 36382 25284
rect 36754 25228 36764 25284
rect 36820 25228 38556 25284
rect 38612 25228 38622 25284
rect 38780 25228 39340 25284
rect 39396 25228 39406 25284
rect 39554 25228 39564 25284
rect 39620 25228 39630 25284
rect 40114 25228 40124 25284
rect 40180 25228 42252 25284
rect 42308 25228 42318 25284
rect 38780 25172 38836 25228
rect 3266 25116 3276 25172
rect 3332 25116 19684 25172
rect 24098 25116 24108 25172
rect 24164 25116 24668 25172
rect 24724 25116 24734 25172
rect 29698 25116 29708 25172
rect 29764 25116 30268 25172
rect 30324 25116 34524 25172
rect 34580 25116 34590 25172
rect 38322 25116 38332 25172
rect 38388 25116 38836 25172
rect 39564 25172 39620 25228
rect 39564 25116 40348 25172
rect 40404 25116 40414 25172
rect 5506 25004 5516 25060
rect 5572 25004 18956 25060
rect 19012 25004 19022 25060
rect 19628 24948 19684 25116
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 20188 25004 30828 25060
rect 30884 25004 30894 25060
rect 33730 25004 33740 25060
rect 33796 25004 37772 25060
rect 37828 25004 37838 25060
rect 20188 24948 20244 25004
rect 43820 24948 43876 25340
rect 48860 25284 48916 25340
rect 51772 25284 51828 25340
rect 56140 25284 56196 25452
rect 45490 25228 45500 25284
rect 45556 25228 46732 25284
rect 46788 25228 46798 25284
rect 46946 25228 46956 25284
rect 47012 25228 48188 25284
rect 48244 25228 48412 25284
rect 48468 25228 48916 25284
rect 49410 25228 49420 25284
rect 49476 25228 50092 25284
rect 50148 25228 50158 25284
rect 50372 25228 51828 25284
rect 52322 25228 52332 25284
rect 52388 25228 52668 25284
rect 52724 25228 52734 25284
rect 56130 25228 56140 25284
rect 56196 25228 56206 25284
rect 50372 25172 50428 25228
rect 2930 24892 2940 24948
rect 2996 24892 8428 24948
rect 19628 24892 20244 24948
rect 21410 24892 21420 24948
rect 21476 24892 22540 24948
rect 22596 24892 22606 24948
rect 25890 24892 25900 24948
rect 25956 24892 26460 24948
rect 26516 24892 27020 24948
rect 27076 24892 27580 24948
rect 27636 24892 27646 24948
rect 29810 24892 29820 24948
rect 29876 24892 30044 24948
rect 30100 24892 30604 24948
rect 30660 24892 43876 24948
rect 43932 25116 44044 25172
rect 44100 25116 44110 25172
rect 48066 25116 48076 25172
rect 48132 25116 48636 25172
rect 48692 25116 50428 25172
rect 52546 25116 52556 25172
rect 52612 25116 54460 25172
rect 54516 25116 54526 25172
rect 55346 25116 55356 25172
rect 55412 25116 55692 25172
rect 55748 25116 55758 25172
rect 55906 25116 55916 25172
rect 55972 25116 57820 25172
rect 57876 25116 58044 25172
rect 58100 25116 58110 25172
rect 8372 24724 8428 24892
rect 21420 24836 21476 24892
rect 43932 24836 43988 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 52770 25004 52780 25060
rect 52836 25004 56028 25060
rect 56084 25004 56094 25060
rect 51650 24892 51660 24948
rect 51716 24892 51996 24948
rect 52052 24892 52062 24948
rect 14690 24780 14700 24836
rect 14756 24780 15260 24836
rect 15316 24780 18844 24836
rect 18900 24780 21476 24836
rect 24658 24780 24668 24836
rect 24724 24780 26908 24836
rect 26964 24780 26974 24836
rect 27794 24780 27804 24836
rect 27860 24780 36204 24836
rect 36260 24780 36270 24836
rect 36754 24780 36764 24836
rect 36820 24780 37324 24836
rect 37380 24780 38668 24836
rect 38724 24780 38734 24836
rect 40562 24780 40572 24836
rect 40628 24780 42420 24836
rect 42578 24780 42588 24836
rect 42644 24780 43988 24836
rect 44156 24780 45948 24836
rect 46004 24780 46956 24836
rect 47012 24780 47022 24836
rect 47170 24780 47180 24836
rect 47236 24780 47852 24836
rect 47908 24780 49980 24836
rect 50036 24780 50046 24836
rect 54114 24780 54124 24836
rect 54180 24780 54796 24836
rect 54852 24780 54862 24836
rect 42364 24724 42420 24780
rect 44156 24724 44212 24780
rect 8372 24668 21196 24724
rect 21252 24668 21262 24724
rect 25666 24668 25676 24724
rect 25732 24668 27916 24724
rect 27972 24668 27982 24724
rect 32722 24668 32732 24724
rect 32788 24668 33628 24724
rect 33684 24668 33694 24724
rect 35970 24668 35980 24724
rect 36036 24668 36046 24724
rect 42364 24668 44212 24724
rect 44370 24668 44380 24724
rect 44436 24668 47292 24724
rect 47348 24668 47358 24724
rect 35980 24612 36036 24668
rect 49980 24612 50036 24780
rect 50306 24668 50316 24724
rect 50372 24668 52108 24724
rect 52164 24668 52174 24724
rect 18274 24556 18284 24612
rect 18340 24556 20636 24612
rect 20692 24556 20702 24612
rect 24882 24556 24892 24612
rect 24948 24556 25788 24612
rect 25844 24556 25854 24612
rect 26852 24556 32732 24612
rect 32788 24556 32798 24612
rect 32946 24556 32956 24612
rect 33012 24556 33404 24612
rect 33460 24556 34076 24612
rect 34132 24556 35924 24612
rect 35980 24556 36764 24612
rect 36820 24556 36830 24612
rect 41430 24556 41468 24612
rect 41524 24556 41534 24612
rect 43922 24556 43932 24612
rect 43988 24556 44604 24612
rect 44660 24556 44670 24612
rect 45378 24556 45388 24612
rect 45444 24556 45948 24612
rect 46004 24556 46014 24612
rect 47618 24556 47628 24612
rect 47684 24556 48748 24612
rect 48804 24556 48814 24612
rect 49980 24556 53228 24612
rect 53284 24556 54908 24612
rect 54964 24556 54974 24612
rect 56130 24556 56140 24612
rect 56196 24556 59388 24612
rect 59444 24556 59454 24612
rect 26852 24500 26908 24556
rect 35868 24500 35924 24556
rect 15092 24444 26908 24500
rect 28466 24444 28476 24500
rect 28532 24444 29708 24500
rect 29764 24444 29774 24500
rect 34290 24444 34300 24500
rect 34356 24444 34972 24500
rect 35028 24444 35420 24500
rect 35476 24444 35486 24500
rect 35868 24444 36316 24500
rect 36372 24444 36382 24500
rect 36530 24444 36540 24500
rect 36596 24444 45724 24500
rect 45780 24444 47740 24500
rect 47796 24444 47806 24500
rect 49634 24444 49644 24500
rect 49700 24444 50204 24500
rect 50260 24444 50270 24500
rect 51734 24444 51772 24500
rect 51828 24444 51838 24500
rect 55458 24444 55468 24500
rect 55524 24444 55804 24500
rect 55860 24444 57036 24500
rect 57092 24444 57372 24500
rect 57428 24444 57438 24500
rect 5058 24332 5068 24388
rect 5124 24332 14364 24388
rect 14420 24332 14430 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 15092 24276 15148 24444
rect 20962 24332 20972 24388
rect 21028 24332 25116 24388
rect 25172 24332 25182 24388
rect 26002 24332 26012 24388
rect 26068 24332 27804 24388
rect 27860 24332 27870 24388
rect 34150 24332 34188 24388
rect 34244 24332 34254 24388
rect 35970 24332 35980 24388
rect 36036 24332 36540 24388
rect 36596 24332 36606 24388
rect 46498 24332 46508 24388
rect 46564 24332 55916 24388
rect 55972 24332 55982 24388
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 11666 24220 11676 24276
rect 11732 24220 15148 24276
rect 22530 24220 22540 24276
rect 22596 24220 22764 24276
rect 22820 24220 23212 24276
rect 23268 24220 23278 24276
rect 44146 24220 44156 24276
rect 44212 24220 45108 24276
rect 45266 24220 45276 24276
rect 45332 24220 47516 24276
rect 47572 24220 52780 24276
rect 52836 24220 52846 24276
rect 45052 24164 45108 24220
rect 9986 24108 9996 24164
rect 10052 24108 25228 24164
rect 25284 24108 25294 24164
rect 33954 24108 33964 24164
rect 34020 24108 34524 24164
rect 34580 24108 44044 24164
rect 44100 24108 44110 24164
rect 45052 24108 45388 24164
rect 45444 24108 48524 24164
rect 48580 24108 48590 24164
rect 48738 24108 48748 24164
rect 48804 24108 49756 24164
rect 49812 24108 49822 24164
rect 55122 24108 55132 24164
rect 55188 24108 56924 24164
rect 56980 24108 57596 24164
rect 57652 24108 57662 24164
rect 21298 23996 21308 24052
rect 21364 23996 24332 24052
rect 24388 23996 26124 24052
rect 26180 23996 26190 24052
rect 32162 23996 32172 24052
rect 32228 23996 39788 24052
rect 39844 23996 39854 24052
rect 41458 23996 41468 24052
rect 41524 23996 46620 24052
rect 46676 23996 47964 24052
rect 48020 23996 49084 24052
rect 49140 23996 49150 24052
rect 49858 23996 49868 24052
rect 49924 23996 50316 24052
rect 50372 23996 50382 24052
rect 50754 23996 50764 24052
rect 50820 23996 51660 24052
rect 51716 23996 57820 24052
rect 57876 23996 57886 24052
rect 17490 23884 17500 23940
rect 17556 23884 18284 23940
rect 18340 23884 18350 23940
rect 22988 23828 23044 23996
rect 34738 23884 34748 23940
rect 34804 23884 34972 23940
rect 35028 23884 35038 23940
rect 36502 23884 36540 23940
rect 36596 23884 36606 23940
rect 42354 23884 42364 23940
rect 42420 23884 43708 23940
rect 43764 23884 43774 23940
rect 46946 23884 46956 23940
rect 47012 23884 50428 23940
rect 50978 23884 50988 23940
rect 51044 23884 52668 23940
rect 52724 23884 52734 23940
rect 52994 23884 53004 23940
rect 53060 23884 53452 23940
rect 53508 23884 53518 23940
rect 50372 23828 50428 23884
rect 22978 23772 22988 23828
rect 23044 23772 23054 23828
rect 33954 23772 33964 23828
rect 34020 23772 35980 23828
rect 36036 23772 36046 23828
rect 36306 23772 36316 23828
rect 36372 23772 37436 23828
rect 37492 23772 37502 23828
rect 44482 23772 44492 23828
rect 44548 23772 45724 23828
rect 45780 23772 45948 23828
rect 46004 23772 46014 23828
rect 47170 23772 47180 23828
rect 47236 23772 47964 23828
rect 48020 23772 48030 23828
rect 50372 23772 51772 23828
rect 51828 23772 51838 23828
rect 53666 23772 53676 23828
rect 53732 23772 54012 23828
rect 54068 23772 54078 23828
rect 21970 23660 21980 23716
rect 22036 23660 23100 23716
rect 23156 23660 24108 23716
rect 24164 23660 24174 23716
rect 28914 23660 28924 23716
rect 28980 23660 30044 23716
rect 30100 23660 31052 23716
rect 31108 23660 31836 23716
rect 31892 23660 34860 23716
rect 34916 23660 36540 23716
rect 36596 23660 36606 23716
rect 41010 23660 41020 23716
rect 41076 23660 41804 23716
rect 41860 23660 41870 23716
rect 41990 23660 42028 23716
rect 42084 23660 42094 23716
rect 42914 23660 42924 23716
rect 42980 23660 45388 23716
rect 45444 23660 45454 23716
rect 45602 23660 45612 23716
rect 45668 23660 46620 23716
rect 46676 23660 46686 23716
rect 47282 23660 47292 23716
rect 47348 23660 50428 23716
rect 50484 23660 51044 23716
rect 51874 23660 51884 23716
rect 51940 23660 52556 23716
rect 52612 23660 53004 23716
rect 53060 23660 53070 23716
rect 53862 23660 53900 23716
rect 53956 23660 53966 23716
rect 21746 23548 21756 23604
rect 21812 23548 24668 23604
rect 24724 23548 26236 23604
rect 26292 23548 27132 23604
rect 27188 23548 27198 23604
rect 30818 23548 30828 23604
rect 30884 23548 31612 23604
rect 31668 23548 31678 23604
rect 34150 23548 34188 23604
rect 34244 23548 34254 23604
rect 35410 23548 35420 23604
rect 35476 23548 36652 23604
rect 36708 23548 36718 23604
rect 37426 23548 37436 23604
rect 37492 23548 40236 23604
rect 40292 23548 43708 23604
rect 43764 23548 43774 23604
rect 43922 23548 43932 23604
rect 43988 23548 44380 23604
rect 44436 23548 47124 23604
rect 47954 23548 47964 23604
rect 48020 23548 50484 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 47068 23492 47124 23548
rect 4946 23436 4956 23492
rect 5012 23436 14308 23492
rect 15362 23436 15372 23492
rect 15428 23436 17948 23492
rect 18004 23436 19404 23492
rect 19460 23436 19470 23492
rect 20290 23436 20300 23492
rect 20356 23436 21308 23492
rect 21364 23436 21374 23492
rect 25330 23436 25340 23492
rect 25396 23436 26124 23492
rect 26180 23436 26190 23492
rect 26852 23436 35532 23492
rect 35588 23436 35598 23492
rect 38658 23436 38668 23492
rect 38724 23436 39676 23492
rect 39732 23436 41468 23492
rect 41524 23436 44268 23492
rect 44324 23436 45836 23492
rect 45892 23436 46284 23492
rect 46340 23436 46508 23492
rect 46564 23436 46574 23492
rect 46732 23436 46844 23492
rect 46900 23436 46910 23492
rect 47068 23436 48300 23492
rect 48356 23436 48366 23492
rect 48962 23436 48972 23492
rect 49028 23436 49532 23492
rect 49588 23436 49598 23492
rect 14252 23380 14308 23436
rect 26852 23380 26908 23436
rect 46732 23380 46788 23436
rect 50428 23380 50484 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 50988 23380 51044 23660
rect 59200 23604 59800 23632
rect 52658 23548 52668 23604
rect 52724 23548 53564 23604
rect 53620 23548 54012 23604
rect 54068 23548 54078 23604
rect 56018 23548 56028 23604
rect 56084 23548 59800 23604
rect 59200 23520 59800 23548
rect 8306 23324 8316 23380
rect 8372 23268 8428 23380
rect 14252 23324 26908 23380
rect 27122 23324 27132 23380
rect 27188 23324 28028 23380
rect 28084 23324 28094 23380
rect 28924 23324 33964 23380
rect 34020 23324 34030 23380
rect 40450 23324 40460 23380
rect 40516 23324 41356 23380
rect 41412 23324 41422 23380
rect 41916 23324 43820 23380
rect 43876 23324 44604 23380
rect 44660 23324 46788 23380
rect 46946 23324 46956 23380
rect 47012 23324 47740 23380
rect 47796 23324 47806 23380
rect 49158 23324 49196 23380
rect 49252 23324 49262 23380
rect 50418 23324 50428 23380
rect 50484 23324 50494 23380
rect 50642 23324 50652 23380
rect 50708 23324 51044 23380
rect 51874 23324 51884 23380
rect 51940 23324 52220 23380
rect 52276 23324 52286 23380
rect 53890 23324 53900 23380
rect 53956 23324 55020 23380
rect 55076 23324 55086 23380
rect 55234 23324 55244 23380
rect 55300 23324 55310 23380
rect 55570 23324 55580 23380
rect 55636 23324 56140 23380
rect 56196 23324 56206 23380
rect 56466 23324 56476 23380
rect 56532 23324 56924 23380
rect 56980 23324 57484 23380
rect 57540 23324 57550 23380
rect 28924 23268 28980 23324
rect 41916 23268 41972 23324
rect 8372 23212 28980 23268
rect 29138 23212 29148 23268
rect 29204 23212 29820 23268
rect 29876 23212 29886 23268
rect 31714 23212 31724 23268
rect 31780 23212 33068 23268
rect 33124 23212 33134 23268
rect 36754 23212 36764 23268
rect 36820 23212 41972 23268
rect 42130 23212 42140 23268
rect 42196 23212 45500 23268
rect 45556 23212 45566 23268
rect 45826 23212 45836 23268
rect 45892 23212 46396 23268
rect 46452 23212 46462 23268
rect 47012 23156 47068 23324
rect 55244 23268 55300 23324
rect 47170 23212 47180 23268
rect 47236 23212 50204 23268
rect 50260 23212 50270 23268
rect 52098 23212 52108 23268
rect 52164 23212 53788 23268
rect 53844 23212 53854 23268
rect 54796 23212 55300 23268
rect 25666 23100 25676 23156
rect 25732 23100 26012 23156
rect 26068 23100 27244 23156
rect 27300 23100 27310 23156
rect 35858 23100 35868 23156
rect 35924 23100 36316 23156
rect 36372 23100 36540 23156
rect 36596 23100 40348 23156
rect 40404 23100 42700 23156
rect 42756 23100 42766 23156
rect 43586 23100 43596 23156
rect 43652 23100 46172 23156
rect 46228 23100 47068 23156
rect 48962 23100 48972 23156
rect 49028 23100 50988 23156
rect 51044 23100 51054 23156
rect 51650 23100 51660 23156
rect 51716 23100 53676 23156
rect 53732 23100 53742 23156
rect 54796 23044 54852 23212
rect 33730 22988 33740 23044
rect 33796 22988 34636 23044
rect 34692 22988 35756 23044
rect 35812 22988 35822 23044
rect 40786 22988 40796 23044
rect 40852 22988 41132 23044
rect 41188 22988 41198 23044
rect 42466 22988 42476 23044
rect 42532 22988 43036 23044
rect 43092 22988 45052 23044
rect 45108 22988 45118 23044
rect 45462 22988 45500 23044
rect 45556 22988 45566 23044
rect 46162 22988 46172 23044
rect 46228 22988 48188 23044
rect 48244 22988 48254 23044
rect 49046 22988 49084 23044
rect 49140 22988 49150 23044
rect 49858 22988 49868 23044
rect 49924 22988 50092 23044
rect 50148 22988 50158 23044
rect 50530 22988 50540 23044
rect 50596 22988 51548 23044
rect 51604 22988 51614 23044
rect 51874 22988 51884 23044
rect 51940 22988 54852 23044
rect 55010 22988 55020 23044
rect 55076 22988 55132 23044
rect 55188 22988 55198 23044
rect 12002 22876 12012 22932
rect 12068 22876 30716 22932
rect 30772 22876 30782 22932
rect 32162 22876 32172 22932
rect 32228 22876 38668 22932
rect 38742 22876 38780 22932
rect 38836 22876 38846 22932
rect 44146 22876 44156 22932
rect 44212 22876 45612 22932
rect 45668 22876 45678 22932
rect 46386 22876 46396 22932
rect 46452 22876 46956 22932
rect 47012 22876 47022 22932
rect 38612 22820 38668 22876
rect 48188 22820 48244 22988
rect 48738 22876 48748 22932
rect 48804 22876 48860 22932
rect 48916 22876 48926 22932
rect 49186 22876 49196 22932
rect 49252 22876 49532 22932
rect 49588 22876 49756 22932
rect 49812 22876 55356 22932
rect 55412 22876 55422 22932
rect 58146 22876 58156 22932
rect 58212 22876 58604 22932
rect 58660 22876 58670 22932
rect 31714 22764 31724 22820
rect 31780 22764 33404 22820
rect 33460 22764 33470 22820
rect 38612 22764 42252 22820
rect 42308 22764 42812 22820
rect 42868 22764 42878 22820
rect 46834 22764 46844 22820
rect 46900 22764 47180 22820
rect 47236 22764 47246 22820
rect 48188 22764 51884 22820
rect 51940 22764 51950 22820
rect 53106 22764 53116 22820
rect 53172 22764 53452 22820
rect 53508 22764 55692 22820
rect 55748 22764 55758 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 10098 22652 10108 22708
rect 10164 22652 29596 22708
rect 29652 22652 29662 22708
rect 31602 22652 31612 22708
rect 31668 22652 34748 22708
rect 34804 22652 34814 22708
rect 36082 22652 36092 22708
rect 36148 22652 36428 22708
rect 36484 22652 37548 22708
rect 37604 22652 37614 22708
rect 37762 22652 37772 22708
rect 37828 22652 42028 22708
rect 42084 22652 42094 22708
rect 43698 22652 43708 22708
rect 43764 22652 47516 22708
rect 47572 22652 51996 22708
rect 52052 22652 53900 22708
rect 53956 22652 53966 22708
rect 30370 22540 30380 22596
rect 30436 22540 34412 22596
rect 34468 22540 34478 22596
rect 35074 22540 35084 22596
rect 35140 22540 35756 22596
rect 35812 22540 42588 22596
rect 42644 22540 43596 22596
rect 43652 22540 43662 22596
rect 44482 22540 44492 22596
rect 44548 22540 49196 22596
rect 49252 22540 49262 22596
rect 49522 22540 49532 22596
rect 49588 22540 52556 22596
rect 52612 22540 52622 22596
rect 54002 22540 54012 22596
rect 54068 22540 55244 22596
rect 55300 22540 55310 22596
rect 23202 22428 23212 22484
rect 23268 22428 23772 22484
rect 23828 22428 25116 22484
rect 25172 22428 25182 22484
rect 33170 22428 33180 22484
rect 33236 22428 37996 22484
rect 38052 22428 38062 22484
rect 40002 22428 40012 22484
rect 40068 22428 40572 22484
rect 40628 22428 40638 22484
rect 47506 22428 47516 22484
rect 47572 22428 49868 22484
rect 49924 22428 54684 22484
rect 54740 22428 54750 22484
rect 28914 22316 28924 22372
rect 28980 22316 29260 22372
rect 29316 22316 29708 22372
rect 29764 22316 32172 22372
rect 32228 22316 32238 22372
rect 33506 22316 33516 22372
rect 33572 22316 35420 22372
rect 35476 22316 35486 22372
rect 38546 22316 38556 22372
rect 38612 22316 38892 22372
rect 38948 22316 38958 22372
rect 40674 22316 40684 22372
rect 40740 22316 41356 22372
rect 41412 22316 42588 22372
rect 42644 22316 43148 22372
rect 43204 22316 44156 22372
rect 44212 22316 44222 22372
rect 46050 22316 46060 22372
rect 46116 22316 46732 22372
rect 46788 22316 46798 22372
rect 48850 22316 48860 22372
rect 48916 22316 49420 22372
rect 49476 22316 49486 22372
rect 52546 22316 52556 22372
rect 52612 22316 53004 22372
rect 53060 22316 55804 22372
rect 55860 22316 55870 22372
rect 56690 22316 56700 22372
rect 56756 22316 57820 22372
rect 57876 22316 57886 22372
rect 200 22260 800 22288
rect 200 22204 1932 22260
rect 1988 22204 1998 22260
rect 17826 22204 17836 22260
rect 17892 22204 18732 22260
rect 18788 22204 18798 22260
rect 33282 22204 33292 22260
rect 33348 22204 34076 22260
rect 34132 22204 34142 22260
rect 34402 22204 34412 22260
rect 34468 22204 39228 22260
rect 39284 22204 40236 22260
rect 40292 22204 40908 22260
rect 40964 22204 40974 22260
rect 41122 22204 41132 22260
rect 41188 22204 43596 22260
rect 43652 22204 43662 22260
rect 45042 22204 45052 22260
rect 45108 22204 45388 22260
rect 45444 22204 45454 22260
rect 46946 22204 46956 22260
rect 47012 22204 48188 22260
rect 48244 22204 53676 22260
rect 53732 22204 53742 22260
rect 54786 22204 54796 22260
rect 54852 22204 56812 22260
rect 56868 22204 56878 22260
rect 200 22176 800 22204
rect 33516 22148 33572 22204
rect 29474 22092 29484 22148
rect 29540 22092 29932 22148
rect 29988 22092 30156 22148
rect 30212 22092 31388 22148
rect 31444 22092 31454 22148
rect 33506 22092 33516 22148
rect 33572 22092 33582 22148
rect 35252 22092 35756 22148
rect 35812 22092 35822 22148
rect 37986 22092 37996 22148
rect 38052 22092 38668 22148
rect 38724 22092 38734 22148
rect 39330 22092 39340 22148
rect 39396 22092 39900 22148
rect 39956 22092 39966 22148
rect 40114 22092 40124 22148
rect 40180 22092 43036 22148
rect 43092 22092 43102 22148
rect 43922 22092 43932 22148
rect 43988 22092 45948 22148
rect 46004 22092 46014 22148
rect 47394 22092 47404 22148
rect 47460 22092 48300 22148
rect 48356 22092 49532 22148
rect 49588 22092 49598 22148
rect 49970 22092 49980 22148
rect 50036 22092 50204 22148
rect 50260 22092 50270 22148
rect 50372 22092 51548 22148
rect 51604 22092 51614 22148
rect 53330 22092 53340 22148
rect 53396 22092 53676 22148
rect 53732 22092 55132 22148
rect 55188 22092 55198 22148
rect 55346 22092 55356 22148
rect 55412 22092 55580 22148
rect 55636 22092 55646 22148
rect 35252 22036 35308 22092
rect 30706 21980 30716 22036
rect 30772 21980 30782 22036
rect 31714 21980 31724 22036
rect 31780 21980 35308 22036
rect 35756 21980 40460 22036
rect 40516 21980 40526 22036
rect 41234 21980 41244 22036
rect 41300 21980 41468 22036
rect 41524 21980 44156 22036
rect 44212 21980 44492 22036
rect 44548 21980 44558 22036
rect 44706 21980 44716 22036
rect 44772 21980 49756 22036
rect 49812 21980 49822 22036
rect 50306 21980 50316 22036
rect 50372 21980 50428 22092
rect 51762 21980 51772 22036
rect 51828 21980 52108 22036
rect 52164 21980 52174 22036
rect 53442 21980 53452 22036
rect 53508 21980 53788 22036
rect 53844 21980 53854 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 30716 21924 30772 21980
rect 35756 21924 35812 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 29810 21868 29820 21924
rect 29876 21868 30156 21924
rect 30212 21868 35812 21924
rect 47012 21868 50148 21924
rect 50978 21868 50988 21924
rect 51044 21868 51324 21924
rect 51380 21868 51390 21924
rect 52658 21868 52668 21924
rect 52724 21868 54236 21924
rect 54292 21868 55132 21924
rect 55188 21868 57708 21924
rect 57764 21868 57774 21924
rect 47012 21812 47068 21868
rect 50092 21812 50148 21868
rect 13122 21756 13132 21812
rect 13188 21756 32228 21812
rect 33730 21756 33740 21812
rect 33796 21756 35980 21812
rect 36036 21756 38780 21812
rect 38836 21756 38948 21812
rect 39442 21756 39452 21812
rect 39508 21756 40236 21812
rect 40292 21756 40302 21812
rect 41906 21756 41916 21812
rect 41972 21756 41982 21812
rect 44034 21756 44044 21812
rect 44100 21756 44380 21812
rect 44436 21756 44446 21812
rect 45490 21756 45500 21812
rect 45556 21756 46732 21812
rect 46788 21756 47068 21812
rect 48066 21756 48076 21812
rect 48132 21756 48300 21812
rect 48356 21756 48366 21812
rect 48962 21756 48972 21812
rect 49028 21756 49420 21812
rect 49476 21756 49486 21812
rect 49634 21756 49644 21812
rect 49700 21756 49756 21812
rect 49812 21756 49822 21812
rect 50092 21756 50652 21812
rect 50708 21756 50718 21812
rect 51202 21756 51212 21812
rect 51268 21756 54516 21812
rect 32172 21700 32228 21756
rect 38892 21700 38948 21756
rect 41916 21700 41972 21756
rect 22642 21644 22652 21700
rect 22708 21644 23100 21700
rect 23156 21644 23324 21700
rect 23380 21644 24780 21700
rect 24836 21644 30044 21700
rect 30100 21644 30110 21700
rect 30930 21644 30940 21700
rect 30996 21644 31948 21700
rect 32004 21644 32014 21700
rect 32172 21644 34524 21700
rect 34580 21644 34590 21700
rect 37090 21644 37100 21700
rect 37156 21644 38668 21700
rect 38724 21644 38734 21700
rect 38892 21644 41972 21700
rect 42354 21644 42364 21700
rect 42420 21644 43932 21700
rect 43988 21644 43998 21700
rect 45378 21644 45388 21700
rect 45444 21644 45948 21700
rect 46004 21644 46014 21700
rect 46162 21644 46172 21700
rect 46228 21644 50316 21700
rect 50372 21644 50382 21700
rect 51426 21644 51436 21700
rect 51492 21644 51660 21700
rect 51716 21644 52108 21700
rect 52164 21644 52174 21700
rect 53218 21644 53228 21700
rect 53284 21644 54236 21700
rect 54292 21644 54302 21700
rect 39452 21588 39508 21644
rect 54460 21588 54516 21756
rect 55010 21644 55020 21700
rect 55076 21644 55244 21700
rect 55300 21644 56476 21700
rect 56532 21644 56542 21700
rect 9426 21532 9436 21588
rect 9492 21532 21196 21588
rect 21252 21532 21262 21588
rect 22418 21532 22428 21588
rect 22484 21532 22988 21588
rect 23044 21532 23054 21588
rect 38098 21532 38108 21588
rect 38164 21532 39284 21588
rect 39442 21532 39452 21588
rect 39508 21532 39518 21588
rect 40450 21532 40460 21588
rect 40516 21532 44492 21588
rect 44548 21532 44558 21588
rect 45042 21532 45052 21588
rect 45108 21532 45612 21588
rect 45668 21532 45678 21588
rect 46946 21532 46956 21588
rect 47012 21532 48748 21588
rect 48804 21532 48814 21588
rect 49186 21532 49196 21588
rect 49252 21532 49532 21588
rect 49588 21532 49598 21588
rect 50082 21532 50092 21588
rect 50148 21532 50988 21588
rect 51044 21532 51100 21588
rect 51156 21532 51166 21588
rect 51874 21532 51884 21588
rect 51940 21532 54124 21588
rect 54180 21532 54190 21588
rect 54460 21532 55748 21588
rect 39228 21476 39284 21532
rect 55692 21476 55748 21532
rect 21746 21420 21756 21476
rect 21812 21420 22316 21476
rect 22372 21420 22382 21476
rect 22530 21420 22540 21476
rect 22596 21420 23436 21476
rect 23492 21420 23502 21476
rect 39228 21420 39564 21476
rect 39620 21420 39630 21476
rect 41010 21420 41020 21476
rect 41076 21420 42476 21476
rect 42532 21420 42542 21476
rect 43138 21420 43148 21476
rect 43204 21420 45164 21476
rect 45220 21420 48860 21476
rect 48916 21420 48926 21476
rect 50306 21420 50316 21476
rect 50372 21420 51212 21476
rect 51268 21420 51278 21476
rect 51426 21420 51436 21476
rect 51492 21420 51548 21476
rect 51604 21420 52668 21476
rect 52724 21420 52734 21476
rect 53190 21420 53228 21476
rect 53284 21420 53294 21476
rect 55682 21420 55692 21476
rect 55748 21420 55758 21476
rect 42476 21364 42532 21420
rect 33618 21308 33628 21364
rect 33684 21308 33964 21364
rect 34020 21308 36428 21364
rect 36484 21308 36494 21364
rect 40898 21308 40908 21364
rect 40964 21308 41916 21364
rect 41972 21308 41982 21364
rect 42476 21308 43036 21364
rect 43092 21308 43102 21364
rect 47012 21308 47964 21364
rect 48020 21308 50932 21364
rect 51090 21308 51100 21364
rect 51156 21308 52668 21364
rect 52724 21308 56364 21364
rect 56420 21308 56430 21364
rect 47012 21252 47068 21308
rect 50876 21252 50932 21308
rect 30594 21196 30604 21252
rect 30660 21196 32620 21252
rect 32676 21196 33180 21252
rect 33236 21196 33246 21252
rect 35532 21196 47068 21252
rect 48290 21196 48300 21252
rect 48356 21196 48748 21252
rect 48804 21196 50820 21252
rect 50876 21196 53228 21252
rect 53284 21196 53294 21252
rect 57474 21196 57484 21252
rect 57540 21196 57550 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 31052 20916 31108 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 35532 21028 35588 21196
rect 50764 21140 50820 21196
rect 57484 21140 57540 21196
rect 38770 21084 38780 21140
rect 38836 21084 41356 21140
rect 41412 21084 41422 21140
rect 41804 21084 45388 21140
rect 45444 21084 46844 21140
rect 46900 21084 46910 21140
rect 49970 21084 49980 21140
rect 50036 21084 50316 21140
rect 50372 21084 50382 21140
rect 50530 21084 50540 21140
rect 50596 21084 50708 21140
rect 50764 21084 51884 21140
rect 51940 21084 51950 21140
rect 57250 21084 57260 21140
rect 57316 21084 57540 21140
rect 41804 21028 41860 21084
rect 50652 21028 50708 21084
rect 31276 20972 32172 21028
rect 32228 20972 32620 21028
rect 32676 20972 32844 21028
rect 32900 20972 35588 21028
rect 36642 20972 36652 21028
rect 36708 20972 41020 21028
rect 41076 20972 41086 21028
rect 41234 20972 41244 21028
rect 41300 20972 41860 21028
rect 42018 20972 42028 21028
rect 42084 20972 44716 21028
rect 44772 20972 46900 21028
rect 48626 20972 48636 21028
rect 48692 20972 49532 21028
rect 49588 20972 49598 21028
rect 49746 20972 49756 21028
rect 49812 20972 50596 21028
rect 50652 20972 50988 21028
rect 51044 20972 51054 21028
rect 53788 20972 55020 21028
rect 55076 20972 56028 21028
rect 56084 20972 56094 21028
rect 31276 20916 31332 20972
rect 46844 20916 46900 20972
rect 50540 20916 50596 20972
rect 53788 20916 53844 20972
rect 6626 20860 6636 20916
rect 6692 20860 26908 20916
rect 31042 20860 31052 20916
rect 31108 20860 31118 20916
rect 31266 20860 31276 20916
rect 31332 20860 31342 20916
rect 35522 20860 35532 20916
rect 35588 20860 43596 20916
rect 43652 20860 43662 20916
rect 44482 20860 44492 20916
rect 44548 20860 46788 20916
rect 46844 20860 50316 20916
rect 50372 20860 50382 20916
rect 50540 20860 53844 20916
rect 54002 20860 54012 20916
rect 54068 20860 54348 20916
rect 54404 20860 54414 20916
rect 26852 20692 26908 20860
rect 46732 20804 46788 20860
rect 29922 20748 29932 20804
rect 29988 20748 30716 20804
rect 30772 20748 30782 20804
rect 38658 20748 38668 20804
rect 38724 20748 39340 20804
rect 39396 20748 39406 20804
rect 42354 20748 42364 20804
rect 42420 20748 43484 20804
rect 43540 20748 43820 20804
rect 43876 20748 43886 20804
rect 46246 20748 46284 20804
rect 46340 20748 46350 20804
rect 46722 20748 46732 20804
rect 46788 20748 49196 20804
rect 49252 20748 49262 20804
rect 49410 20748 49420 20804
rect 49476 20748 54124 20804
rect 54180 20748 54190 20804
rect 24994 20636 25004 20692
rect 25060 20636 25564 20692
rect 25620 20636 26124 20692
rect 26180 20636 26460 20692
rect 26516 20636 26684 20692
rect 26740 20636 26750 20692
rect 26852 20636 35644 20692
rect 35700 20636 35710 20692
rect 36194 20636 36204 20692
rect 36260 20636 36988 20692
rect 37044 20636 37054 20692
rect 38434 20636 38444 20692
rect 38500 20636 43708 20692
rect 43764 20636 43774 20692
rect 44034 20636 44044 20692
rect 44100 20636 47068 20692
rect 47124 20636 47134 20692
rect 48626 20636 48636 20692
rect 48692 20636 50148 20692
rect 50278 20636 50316 20692
rect 50372 20636 50382 20692
rect 50652 20636 54572 20692
rect 54628 20636 54638 20692
rect 50092 20580 50148 20636
rect 50652 20580 50708 20636
rect 2706 20524 2716 20580
rect 2772 20524 3276 20580
rect 3332 20524 16604 20580
rect 16660 20524 16670 20580
rect 23426 20524 23436 20580
rect 23492 20524 23996 20580
rect 24052 20524 24444 20580
rect 24500 20524 24510 20580
rect 26002 20524 26012 20580
rect 26068 20524 27244 20580
rect 27300 20524 27916 20580
rect 27972 20524 27982 20580
rect 31154 20524 31164 20580
rect 31220 20524 31836 20580
rect 31892 20524 31902 20580
rect 38444 20524 40348 20580
rect 40404 20524 40414 20580
rect 42130 20524 42140 20580
rect 42196 20524 44156 20580
rect 44212 20524 44222 20580
rect 48738 20524 48748 20580
rect 48804 20524 49084 20580
rect 49140 20524 49150 20580
rect 50082 20524 50092 20580
rect 50148 20524 50708 20580
rect 50866 20524 50876 20580
rect 50932 20524 52108 20580
rect 52164 20524 52174 20580
rect 52994 20524 53004 20580
rect 53060 20524 53452 20580
rect 53508 20524 53518 20580
rect 55542 20524 55580 20580
rect 55636 20524 55646 20580
rect 38444 20468 38500 20524
rect 24098 20412 24108 20468
rect 24164 20412 24780 20468
rect 24836 20412 28252 20468
rect 28308 20412 28318 20468
rect 34626 20412 34636 20468
rect 34692 20412 36652 20468
rect 36708 20412 36718 20468
rect 38434 20412 38444 20468
rect 38500 20412 38510 20468
rect 43026 20412 43036 20468
rect 43092 20412 46788 20468
rect 48822 20412 48860 20468
rect 48916 20412 48926 20468
rect 49634 20412 49644 20468
rect 49700 20412 50428 20468
rect 50978 20412 50988 20468
rect 51044 20412 51772 20468
rect 51828 20412 52220 20468
rect 52276 20412 52286 20468
rect 54114 20412 54124 20468
rect 54180 20412 54684 20468
rect 54740 20412 54750 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 46732 20356 46788 20412
rect 30034 20300 30044 20356
rect 30100 20300 34300 20356
rect 34356 20300 34366 20356
rect 34514 20300 34524 20356
rect 34580 20300 35868 20356
rect 35924 20300 35934 20356
rect 39414 20300 39452 20356
rect 39508 20300 39518 20356
rect 40898 20300 40908 20356
rect 40964 20300 42476 20356
rect 42532 20300 42542 20356
rect 43698 20300 43708 20356
rect 43764 20300 44156 20356
rect 44212 20300 44380 20356
rect 44436 20300 44446 20356
rect 46722 20300 46732 20356
rect 46788 20300 46798 20356
rect 50372 20244 50428 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 50988 20300 53452 20356
rect 53508 20300 56588 20356
rect 56644 20300 56654 20356
rect 50988 20244 51044 20300
rect 27122 20188 27132 20244
rect 27188 20188 27198 20244
rect 33954 20188 33964 20244
rect 34020 20188 34972 20244
rect 35028 20188 35038 20244
rect 35410 20188 35420 20244
rect 35476 20188 35756 20244
rect 35812 20188 36204 20244
rect 36260 20188 36270 20244
rect 37314 20188 37324 20244
rect 37380 20188 37772 20244
rect 37828 20188 39900 20244
rect 39956 20188 39966 20244
rect 42242 20188 42252 20244
rect 42308 20188 45500 20244
rect 45556 20188 45566 20244
rect 48626 20188 48636 20244
rect 48692 20188 48702 20244
rect 50372 20188 51044 20244
rect 52770 20188 52780 20244
rect 52836 20188 53340 20244
rect 53396 20188 53406 20244
rect 54338 20188 54348 20244
rect 54404 20188 55916 20244
rect 55972 20188 57484 20244
rect 57540 20188 57550 20244
rect 27132 20132 27188 20188
rect 48636 20132 48692 20188
rect 24322 20076 24332 20132
rect 24388 20076 25564 20132
rect 25620 20076 25900 20132
rect 25956 20076 25966 20132
rect 27132 20076 28140 20132
rect 28196 20076 28206 20132
rect 28690 20076 28700 20132
rect 28756 20076 29932 20132
rect 29988 20076 35532 20132
rect 35588 20076 35598 20132
rect 37202 20076 37212 20132
rect 37268 20076 39004 20132
rect 39060 20076 39070 20132
rect 39554 20076 39564 20132
rect 39620 20076 40348 20132
rect 40404 20076 47516 20132
rect 47572 20076 48692 20132
rect 50754 20076 50764 20132
rect 50820 20076 51100 20132
rect 51156 20076 51324 20132
rect 51380 20076 51390 20132
rect 52098 20076 52108 20132
rect 52164 20076 53676 20132
rect 53732 20076 53742 20132
rect 27132 20020 27188 20076
rect 26674 19964 26684 20020
rect 26740 19964 27188 20020
rect 28354 19964 28364 20020
rect 28420 19964 30716 20020
rect 30772 19964 30782 20020
rect 30940 19964 37884 20020
rect 37940 19964 37950 20020
rect 38098 19964 38108 20020
rect 38164 19964 42252 20020
rect 42308 19964 42318 20020
rect 43698 19964 43708 20020
rect 43764 19964 45500 20020
rect 45556 19964 46396 20020
rect 46452 19964 46462 20020
rect 46610 19964 46620 20020
rect 46676 19964 48188 20020
rect 48244 19964 48254 20020
rect 48514 19964 48524 20020
rect 48580 19964 48636 20020
rect 48692 19964 48702 20020
rect 51202 19964 51212 20020
rect 51268 19964 51548 20020
rect 51604 19964 51614 20020
rect 52882 19964 52892 20020
rect 52948 19964 53788 20020
rect 53844 19964 54460 20020
rect 54516 19964 54526 20020
rect 54786 19964 54796 20020
rect 54852 19964 55132 20020
rect 55188 19964 55244 20020
rect 55300 19964 55310 20020
rect 30940 19908 30996 19964
rect 22194 19852 22204 19908
rect 22260 19852 23548 19908
rect 23604 19852 28700 19908
rect 28756 19852 28766 19908
rect 29810 19852 29820 19908
rect 29876 19852 30996 19908
rect 33506 19852 33516 19908
rect 33572 19852 35196 19908
rect 35252 19852 35262 19908
rect 36082 19852 36092 19908
rect 36148 19852 43820 19908
rect 43876 19852 43886 19908
rect 44230 19852 44268 19908
rect 44324 19852 44334 19908
rect 45602 19852 45612 19908
rect 45668 19852 46172 19908
rect 46228 19852 46238 19908
rect 48962 19852 48972 19908
rect 49028 19852 49084 19908
rect 49140 19852 49150 19908
rect 51314 19852 51324 19908
rect 51380 19852 51884 19908
rect 51940 19852 51950 19908
rect 26852 19740 28028 19796
rect 28084 19740 35588 19796
rect 37090 19740 37100 19796
rect 37156 19740 37884 19796
rect 37940 19740 39452 19796
rect 39508 19740 39518 19796
rect 39890 19740 39900 19796
rect 39956 19740 40684 19796
rect 40740 19740 40750 19796
rect 41122 19740 41132 19796
rect 41188 19740 41468 19796
rect 41524 19740 41534 19796
rect 45602 19740 45612 19796
rect 45668 19740 48412 19796
rect 48468 19740 48478 19796
rect 48850 19740 48860 19796
rect 48916 19740 49868 19796
rect 49924 19740 57932 19796
rect 57988 19740 57998 19796
rect 26852 19684 26908 19740
rect 26562 19628 26572 19684
rect 26628 19628 26908 19684
rect 27682 19628 27692 19684
rect 27748 19628 30380 19684
rect 30436 19628 30446 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 35532 19572 35588 19740
rect 41468 19684 41524 19740
rect 41468 19628 46284 19684
rect 46340 19628 46508 19684
rect 46564 19628 46574 19684
rect 47058 19628 47068 19684
rect 47124 19628 50540 19684
rect 50596 19628 51772 19684
rect 51828 19628 56028 19684
rect 56084 19628 56094 19684
rect 34178 19516 34188 19572
rect 34244 19516 34300 19572
rect 34356 19516 34366 19572
rect 35532 19516 38108 19572
rect 38164 19516 38174 19572
rect 38770 19516 38780 19572
rect 38836 19516 39228 19572
rect 39284 19516 40684 19572
rect 40740 19516 40750 19572
rect 42354 19516 42364 19572
rect 42420 19516 44828 19572
rect 44884 19516 45052 19572
rect 45108 19516 45118 19572
rect 45266 19516 45276 19572
rect 45332 19516 45370 19572
rect 47058 19516 47068 19572
rect 47124 19516 48076 19572
rect 48132 19516 48142 19572
rect 48514 19516 48524 19572
rect 48580 19516 49196 19572
rect 49252 19516 52892 19572
rect 52948 19516 52958 19572
rect 53330 19516 53340 19572
rect 53396 19516 55356 19572
rect 55412 19516 55422 19572
rect 48076 19460 48132 19516
rect 34290 19404 34300 19460
rect 34356 19404 34972 19460
rect 35028 19404 36316 19460
rect 36372 19404 36382 19460
rect 38612 19404 39340 19460
rect 39396 19404 39406 19460
rect 40786 19404 40796 19460
rect 40852 19404 47292 19460
rect 47348 19404 47358 19460
rect 48076 19404 49980 19460
rect 50036 19404 50540 19460
rect 50596 19404 50606 19460
rect 50866 19404 50876 19460
rect 50932 19404 50988 19460
rect 51044 19404 51054 19460
rect 51202 19404 51212 19460
rect 51268 19404 51324 19460
rect 51380 19404 51390 19460
rect 51650 19404 51660 19460
rect 51716 19404 51996 19460
rect 52052 19404 52062 19460
rect 55458 19404 55468 19460
rect 55524 19404 55580 19460
rect 55636 19404 55646 19460
rect 38612 19348 38668 19404
rect 24434 19292 24444 19348
rect 24500 19292 26572 19348
rect 26628 19292 26638 19348
rect 31042 19292 31052 19348
rect 31108 19292 31836 19348
rect 31892 19292 32396 19348
rect 32452 19292 32462 19348
rect 32722 19292 32732 19348
rect 32788 19292 38668 19348
rect 39218 19292 39228 19348
rect 39284 19292 40012 19348
rect 40068 19292 42028 19348
rect 42084 19292 42094 19348
rect 42802 19292 42812 19348
rect 42868 19292 45164 19348
rect 45220 19292 45230 19348
rect 46386 19292 46396 19348
rect 46452 19292 49420 19348
rect 49476 19292 49486 19348
rect 49858 19292 49868 19348
rect 49924 19292 51996 19348
rect 52052 19292 52062 19348
rect 55318 19292 55356 19348
rect 55412 19292 57260 19348
rect 57316 19292 57326 19348
rect 31266 19180 31276 19236
rect 31332 19180 31948 19236
rect 32004 19180 32014 19236
rect 33618 19180 33628 19236
rect 33684 19180 34076 19236
rect 34132 19180 34860 19236
rect 34916 19180 34926 19236
rect 38322 19180 38332 19236
rect 38388 19180 38892 19236
rect 38948 19180 39676 19236
rect 39732 19180 39742 19236
rect 43250 19180 43260 19236
rect 43316 19180 43708 19236
rect 43764 19180 43774 19236
rect 44370 19180 44380 19236
rect 44436 19180 44940 19236
rect 44996 19180 45006 19236
rect 45266 19180 45276 19236
rect 45332 19180 46172 19236
rect 46228 19180 50260 19236
rect 50978 19180 50988 19236
rect 51044 19180 51212 19236
rect 51268 19180 51772 19236
rect 51828 19180 51838 19236
rect 55458 19180 55468 19236
rect 55524 19180 56140 19236
rect 56196 19180 56206 19236
rect 50204 19124 50260 19180
rect 20850 19068 20860 19124
rect 20916 19068 21644 19124
rect 21700 19068 21710 19124
rect 30146 19068 30156 19124
rect 30212 19068 30604 19124
rect 30660 19068 30828 19124
rect 30884 19068 31388 19124
rect 31444 19068 33516 19124
rect 33572 19068 33582 19124
rect 34738 19068 34748 19124
rect 34804 19068 36540 19124
rect 36596 19068 38668 19124
rect 39106 19068 39116 19124
rect 39172 19068 40012 19124
rect 40068 19068 43596 19124
rect 43652 19068 43662 19124
rect 45910 19068 45948 19124
rect 46004 19068 46014 19124
rect 47618 19068 47628 19124
rect 47684 19068 48188 19124
rect 48244 19068 49980 19124
rect 50036 19068 50046 19124
rect 50204 19068 51100 19124
rect 51156 19068 51166 19124
rect 51510 19068 51548 19124
rect 51604 19068 51614 19124
rect 54338 19068 54348 19124
rect 54404 19068 54908 19124
rect 54964 19068 55132 19124
rect 55188 19068 55198 19124
rect 38612 19012 38668 19068
rect 18946 18956 18956 19012
rect 19012 18956 22092 19012
rect 22148 18956 22158 19012
rect 28690 18956 28700 19012
rect 28756 18956 31724 19012
rect 31780 18956 31790 19012
rect 35522 18956 35532 19012
rect 35588 18956 37996 19012
rect 38052 18956 38062 19012
rect 38612 18956 39004 19012
rect 39060 18956 41580 19012
rect 41636 18956 41646 19012
rect 42252 18956 48972 19012
rect 49028 18956 49038 19012
rect 49186 18956 49196 19012
rect 49252 18956 51828 19012
rect 51986 18956 51996 19012
rect 52052 18956 54012 19012
rect 54068 18956 54078 19012
rect 42252 18900 42308 18956
rect 51772 18900 51828 18956
rect 21298 18844 21308 18900
rect 21364 18844 26460 18900
rect 26516 18844 26526 18900
rect 39554 18844 39564 18900
rect 39620 18844 42308 18900
rect 44146 18844 44156 18900
rect 44212 18844 45724 18900
rect 45780 18844 49476 18900
rect 51772 18844 51996 18900
rect 52052 18844 53900 18900
rect 53956 18844 54796 18900
rect 54852 18844 54862 18900
rect 55234 18844 55244 18900
rect 55300 18844 55356 18900
rect 55412 18844 55422 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 26562 18732 26572 18788
rect 26628 18732 28476 18788
rect 28532 18732 28542 18788
rect 36866 18732 36876 18788
rect 36932 18732 42140 18788
rect 42196 18732 42812 18788
rect 42868 18732 42878 18788
rect 43586 18732 43596 18788
rect 43652 18732 45612 18788
rect 45668 18732 45678 18788
rect 48178 18732 48188 18788
rect 48244 18732 49196 18788
rect 49252 18732 49262 18788
rect 26898 18620 26908 18676
rect 26964 18620 27244 18676
rect 27300 18620 27580 18676
rect 27636 18620 29820 18676
rect 29876 18620 29886 18676
rect 33394 18620 33404 18676
rect 33460 18620 40068 18676
rect 40786 18620 40796 18676
rect 40852 18620 40862 18676
rect 42214 18620 42252 18676
rect 42308 18620 42318 18676
rect 43138 18620 43148 18676
rect 43204 18620 43932 18676
rect 43988 18620 43998 18676
rect 48374 18620 48412 18676
rect 48468 18620 48478 18676
rect 23202 18508 23212 18564
rect 23268 18508 24220 18564
rect 24276 18508 24286 18564
rect 26450 18508 26460 18564
rect 26516 18508 27692 18564
rect 27748 18508 27758 18564
rect 31602 18508 31612 18564
rect 31668 18508 33068 18564
rect 33124 18508 34020 18564
rect 34850 18508 34860 18564
rect 34916 18508 35308 18564
rect 35364 18508 35374 18564
rect 36082 18508 36092 18564
rect 36148 18508 37100 18564
rect 37156 18508 37884 18564
rect 37940 18508 37950 18564
rect 38210 18508 38220 18564
rect 38276 18508 38556 18564
rect 38612 18508 39004 18564
rect 39060 18508 39070 18564
rect 16594 18396 16604 18452
rect 16660 18396 18172 18452
rect 18228 18396 18238 18452
rect 21186 18396 21196 18452
rect 21252 18396 22204 18452
rect 22260 18396 22652 18452
rect 22708 18396 22718 18452
rect 26114 18396 26124 18452
rect 26180 18396 27804 18452
rect 27860 18396 29260 18452
rect 29316 18396 29326 18452
rect 31938 18396 31948 18452
rect 32004 18396 32620 18452
rect 32676 18396 32686 18452
rect 33964 18340 34020 18508
rect 40012 18452 40068 18620
rect 40796 18452 40852 18620
rect 49420 18564 49476 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 50978 18732 50988 18788
rect 51044 18732 53900 18788
rect 53956 18732 54348 18788
rect 54404 18732 58268 18788
rect 58324 18732 58334 18788
rect 49970 18620 49980 18676
rect 50036 18620 51660 18676
rect 51716 18620 51726 18676
rect 54450 18620 54460 18676
rect 54516 18620 55692 18676
rect 55748 18620 57540 18676
rect 57484 18564 57540 18620
rect 42130 18508 42140 18564
rect 42196 18508 44044 18564
rect 44100 18508 44110 18564
rect 44370 18508 44380 18564
rect 44436 18508 44828 18564
rect 44884 18508 45276 18564
rect 45332 18508 45342 18564
rect 48290 18508 48300 18564
rect 48356 18508 48636 18564
rect 48692 18508 48702 18564
rect 48962 18508 48972 18564
rect 49028 18508 49252 18564
rect 49420 18508 50988 18564
rect 51044 18508 51054 18564
rect 52658 18508 52668 18564
rect 52724 18508 54460 18564
rect 54516 18508 56252 18564
rect 56308 18508 56318 18564
rect 57474 18508 57484 18564
rect 57540 18508 58828 18564
rect 58884 18508 58894 18564
rect 49196 18452 49252 18508
rect 35074 18396 35084 18452
rect 35140 18396 35756 18452
rect 35812 18396 35822 18452
rect 36306 18396 36316 18452
rect 36372 18396 36540 18452
rect 36596 18396 36606 18452
rect 37538 18396 37548 18452
rect 37604 18396 38108 18452
rect 38164 18396 38174 18452
rect 40002 18396 40012 18452
rect 40068 18396 40078 18452
rect 40338 18396 40348 18452
rect 40404 18396 41804 18452
rect 41860 18396 41870 18452
rect 43810 18396 43820 18452
rect 43876 18396 44268 18452
rect 44324 18396 44492 18452
rect 44548 18396 44558 18452
rect 45826 18396 45836 18452
rect 45892 18396 46620 18452
rect 46676 18396 48972 18452
rect 49028 18396 49038 18452
rect 49196 18396 49644 18452
rect 49700 18396 49710 18452
rect 50754 18396 50764 18452
rect 50820 18396 50988 18452
rect 51044 18396 51054 18452
rect 51314 18396 51324 18452
rect 51380 18396 51884 18452
rect 51940 18396 52780 18452
rect 52836 18396 52846 18452
rect 53638 18396 53676 18452
rect 53732 18396 53742 18452
rect 53890 18396 53900 18452
rect 53956 18396 53994 18452
rect 54450 18396 54460 18452
rect 54516 18396 55468 18452
rect 55524 18396 56476 18452
rect 56532 18396 56542 18452
rect 45836 18340 45892 18396
rect 22754 18284 22764 18340
rect 22820 18284 24332 18340
rect 24388 18284 24398 18340
rect 28018 18284 28028 18340
rect 28084 18284 28812 18340
rect 28868 18284 28878 18340
rect 31826 18284 31836 18340
rect 31892 18284 32396 18340
rect 32452 18284 32462 18340
rect 33926 18284 33964 18340
rect 34020 18284 34030 18340
rect 35970 18284 35980 18340
rect 36036 18284 37436 18340
rect 37492 18284 37996 18340
rect 38052 18284 38062 18340
rect 38882 18284 38892 18340
rect 38948 18284 39228 18340
rect 39284 18284 39900 18340
rect 39956 18284 39966 18340
rect 42242 18284 42252 18340
rect 42308 18284 42700 18340
rect 42756 18284 42766 18340
rect 44706 18284 44716 18340
rect 44772 18284 45892 18340
rect 46722 18284 46732 18340
rect 46788 18284 48860 18340
rect 48916 18284 53340 18340
rect 53396 18284 53406 18340
rect 54674 18284 54684 18340
rect 54740 18284 56588 18340
rect 56644 18284 57148 18340
rect 57204 18284 57708 18340
rect 57764 18284 57774 18340
rect 58034 18284 58044 18340
rect 58100 18284 58492 18340
rect 58548 18284 58558 18340
rect 59200 18228 59800 18256
rect 24546 18172 24556 18228
rect 24612 18172 25788 18228
rect 25844 18172 25854 18228
rect 29586 18172 29596 18228
rect 29652 18172 37212 18228
rect 37268 18172 37278 18228
rect 39106 18172 39116 18228
rect 39172 18172 39452 18228
rect 39508 18172 39518 18228
rect 41906 18172 41916 18228
rect 41972 18172 42252 18228
rect 42308 18172 42318 18228
rect 42466 18172 42476 18228
rect 42532 18172 43708 18228
rect 43764 18172 43774 18228
rect 45714 18172 45724 18228
rect 45780 18172 46172 18228
rect 46228 18172 46238 18228
rect 48290 18172 48300 18228
rect 48356 18172 48524 18228
rect 48580 18172 48590 18228
rect 49746 18172 49756 18228
rect 49812 18172 49980 18228
rect 50036 18172 55580 18228
rect 55636 18172 55646 18228
rect 55906 18172 55916 18228
rect 55972 18172 59800 18228
rect 59200 18144 59800 18172
rect 25890 18060 25900 18116
rect 25956 18060 30492 18116
rect 30548 18060 30558 18116
rect 40226 18060 40236 18116
rect 40292 18060 42812 18116
rect 42868 18060 44156 18116
rect 44212 18060 44222 18116
rect 50978 18060 50988 18116
rect 51044 18060 51324 18116
rect 51380 18060 52108 18116
rect 52164 18060 52444 18116
rect 52500 18060 52510 18116
rect 52770 18060 52780 18116
rect 52836 18060 58044 18116
rect 58100 18060 58110 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 35532 17948 36988 18004
rect 37044 17948 37054 18004
rect 37426 17948 37436 18004
rect 37492 17948 41132 18004
rect 41188 17948 41198 18004
rect 49634 17948 49644 18004
rect 49700 17948 51324 18004
rect 51380 17948 52332 18004
rect 52388 17948 52556 18004
rect 52612 17948 52622 18004
rect 53218 17948 53228 18004
rect 53284 17948 54124 18004
rect 54180 17948 54190 18004
rect 35532 17892 35588 17948
rect 16706 17836 16716 17892
rect 16772 17836 17500 17892
rect 17556 17836 17566 17892
rect 22866 17836 22876 17892
rect 22932 17836 26124 17892
rect 26180 17836 26190 17892
rect 30818 17836 30828 17892
rect 30884 17836 31164 17892
rect 31220 17836 32508 17892
rect 32564 17836 32956 17892
rect 33012 17836 34748 17892
rect 34804 17836 35588 17892
rect 35970 17836 35980 17892
rect 36036 17836 36046 17892
rect 38770 17836 38780 17892
rect 38836 17836 39004 17892
rect 39060 17836 39070 17892
rect 39890 17836 39900 17892
rect 39956 17836 41244 17892
rect 41300 17836 41310 17892
rect 44370 17836 44380 17892
rect 44436 17836 48860 17892
rect 48916 17836 50932 17892
rect 15138 17724 15148 17780
rect 15204 17724 16268 17780
rect 16324 17724 16334 17780
rect 19842 17724 19852 17780
rect 19908 17724 20524 17780
rect 20580 17724 23212 17780
rect 23268 17724 23278 17780
rect 24322 17724 24332 17780
rect 24388 17724 24892 17780
rect 24948 17724 24958 17780
rect 27570 17724 27580 17780
rect 27636 17724 31500 17780
rect 31556 17724 31566 17780
rect 35980 17668 36036 17836
rect 39900 17668 39956 17836
rect 50876 17780 50932 17836
rect 46050 17724 46060 17780
rect 46116 17724 50428 17780
rect 50866 17724 50876 17780
rect 50932 17724 51268 17780
rect 51762 17724 51772 17780
rect 51828 17724 56028 17780
rect 56084 17724 56094 17780
rect 50372 17668 50428 17724
rect 51212 17668 51268 17724
rect 15922 17612 15932 17668
rect 15988 17612 16828 17668
rect 16884 17612 17836 17668
rect 17892 17612 17902 17668
rect 20290 17612 20300 17668
rect 20356 17612 21420 17668
rect 21476 17612 22652 17668
rect 22708 17612 22718 17668
rect 23874 17612 23884 17668
rect 23940 17612 25900 17668
rect 25956 17612 25966 17668
rect 26786 17612 26796 17668
rect 26852 17612 27524 17668
rect 32386 17612 32396 17668
rect 32452 17612 34412 17668
rect 34468 17612 36036 17668
rect 39218 17612 39228 17668
rect 39284 17612 39956 17668
rect 42242 17612 42252 17668
rect 42308 17612 42812 17668
rect 42868 17612 42878 17668
rect 46162 17612 46172 17668
rect 46228 17612 46620 17668
rect 46676 17612 47404 17668
rect 47460 17612 47470 17668
rect 49532 17612 49644 17668
rect 49700 17612 49710 17668
rect 50372 17612 50596 17668
rect 51202 17612 51212 17668
rect 51268 17612 51278 17668
rect 53442 17612 53452 17668
rect 53508 17612 54236 17668
rect 54292 17612 54302 17668
rect 54786 17612 54796 17668
rect 54852 17612 54908 17668
rect 54964 17612 55132 17668
rect 55188 17612 55198 17668
rect 22652 17556 22708 17612
rect 27468 17556 27524 17612
rect 49532 17556 49588 17612
rect 18610 17500 18620 17556
rect 18676 17500 20188 17556
rect 20244 17500 20254 17556
rect 22652 17500 24668 17556
rect 24724 17500 24734 17556
rect 27458 17500 27468 17556
rect 27524 17500 28252 17556
rect 28308 17500 28318 17556
rect 28466 17500 28476 17556
rect 28532 17500 29484 17556
rect 29540 17500 29550 17556
rect 29698 17500 29708 17556
rect 29764 17500 29932 17556
rect 29988 17500 30380 17556
rect 30436 17500 30446 17556
rect 33730 17500 33740 17556
rect 33796 17500 36988 17556
rect 37044 17500 37054 17556
rect 37650 17500 37660 17556
rect 37716 17500 40460 17556
rect 40516 17500 40526 17556
rect 44370 17500 44380 17556
rect 44436 17500 44828 17556
rect 44884 17500 44894 17556
rect 45154 17500 45164 17556
rect 45220 17500 49588 17556
rect 49718 17500 49756 17556
rect 49812 17500 49822 17556
rect 50540 17444 50596 17612
rect 50978 17500 50988 17556
rect 51044 17500 56700 17556
rect 56756 17500 57036 17556
rect 57092 17500 57102 17556
rect 16258 17388 16268 17444
rect 16324 17388 16940 17444
rect 16996 17388 17612 17444
rect 17668 17388 18508 17444
rect 18564 17388 18574 17444
rect 22082 17388 22092 17444
rect 22148 17388 23996 17444
rect 24052 17388 24062 17444
rect 26674 17388 26684 17444
rect 26740 17388 27580 17444
rect 27636 17388 27646 17444
rect 28802 17388 28812 17444
rect 28868 17388 33628 17444
rect 33684 17388 33694 17444
rect 33842 17388 33852 17444
rect 33908 17388 34524 17444
rect 34580 17388 34590 17444
rect 36082 17388 36092 17444
rect 36148 17388 38668 17444
rect 38724 17388 38734 17444
rect 41234 17388 41244 17444
rect 41300 17388 50316 17444
rect 50372 17388 50382 17444
rect 50540 17388 51884 17444
rect 51940 17388 51950 17444
rect 53330 17388 53340 17444
rect 53396 17388 54236 17444
rect 54292 17388 56476 17444
rect 56532 17388 56542 17444
rect 26114 17276 26124 17332
rect 26180 17276 26908 17332
rect 26964 17276 28028 17332
rect 28084 17276 28094 17332
rect 30818 17276 30828 17332
rect 30884 17276 31948 17332
rect 32004 17276 32014 17332
rect 33282 17276 33292 17332
rect 33348 17276 35084 17332
rect 35140 17276 35150 17332
rect 35970 17276 35980 17332
rect 36036 17276 36316 17332
rect 36372 17276 36382 17332
rect 36978 17276 36988 17332
rect 37044 17276 37660 17332
rect 37716 17276 37726 17332
rect 42914 17276 42924 17332
rect 42980 17276 43148 17332
rect 43204 17276 43214 17332
rect 43922 17276 43932 17332
rect 43988 17276 44268 17332
rect 44324 17276 46060 17332
rect 46116 17276 46126 17332
rect 47506 17276 47516 17332
rect 47572 17276 48300 17332
rect 48356 17276 48366 17332
rect 51762 17276 51772 17332
rect 51828 17276 51884 17332
rect 51940 17276 51950 17332
rect 53218 17276 53228 17332
rect 53284 17276 54908 17332
rect 54964 17276 54974 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 24882 17164 24892 17220
rect 24948 17164 25564 17220
rect 25620 17164 25630 17220
rect 31154 17164 31164 17220
rect 31220 17164 34524 17220
rect 34580 17164 34590 17220
rect 34748 17164 37772 17220
rect 37828 17164 38108 17220
rect 38164 17164 38174 17220
rect 39890 17164 39900 17220
rect 39956 17164 40684 17220
rect 40740 17164 40750 17220
rect 42578 17164 42588 17220
rect 42644 17164 43372 17220
rect 43428 17164 45444 17220
rect 47506 17164 47516 17220
rect 47572 17164 48748 17220
rect 48804 17164 48814 17220
rect 48962 17164 48972 17220
rect 49028 17164 50428 17220
rect 51958 17164 51996 17220
rect 52052 17164 52062 17220
rect 34748 17108 34804 17164
rect 45388 17108 45444 17164
rect 50372 17108 50428 17164
rect 2706 17052 2716 17108
rect 2772 17052 3276 17108
rect 3332 17052 7532 17108
rect 7588 17052 7598 17108
rect 17826 17052 17836 17108
rect 17892 17052 22988 17108
rect 23044 17052 23054 17108
rect 25330 17052 25340 17108
rect 25396 17052 25900 17108
rect 25956 17052 26460 17108
rect 26516 17052 26526 17108
rect 31266 17052 31276 17108
rect 31332 17052 31612 17108
rect 31668 17052 32396 17108
rect 32452 17052 32462 17108
rect 33394 17052 33404 17108
rect 33460 17052 34748 17108
rect 34804 17052 34814 17108
rect 34962 17052 34972 17108
rect 35028 17052 35308 17108
rect 35364 17052 36484 17108
rect 36754 17052 36764 17108
rect 36820 17052 37548 17108
rect 37604 17052 37614 17108
rect 37986 17052 37996 17108
rect 38052 17052 41580 17108
rect 41636 17052 41646 17108
rect 41906 17052 41916 17108
rect 41972 17052 43596 17108
rect 43652 17052 43662 17108
rect 45378 17052 45388 17108
rect 45444 17052 45612 17108
rect 45668 17052 45678 17108
rect 45826 17052 45836 17108
rect 45892 17052 49420 17108
rect 49476 17052 49486 17108
rect 50372 17052 52332 17108
rect 52388 17052 52668 17108
rect 52724 17052 53004 17108
rect 53060 17052 53070 17108
rect 53778 17052 53788 17108
rect 53844 17052 53854 17108
rect 54002 17052 54012 17108
rect 54068 17052 55468 17108
rect 55524 17052 55534 17108
rect 36428 16996 36484 17052
rect 53788 16996 53844 17052
rect 23202 16940 23212 16996
rect 23268 16940 23660 16996
rect 23716 16940 24220 16996
rect 24276 16940 26236 16996
rect 26292 16940 26302 16996
rect 32610 16940 32620 16996
rect 32676 16940 36204 16996
rect 36260 16940 36270 16996
rect 36428 16940 37436 16996
rect 37492 16940 37502 16996
rect 38210 16940 38220 16996
rect 38276 16940 38780 16996
rect 38836 16940 39676 16996
rect 39732 16940 39742 16996
rect 40674 16940 40684 16996
rect 40740 16940 42588 16996
rect 42644 16940 42654 16996
rect 44706 16940 44716 16996
rect 44772 16940 47852 16996
rect 47908 16940 47918 16996
rect 53442 16940 53452 16996
rect 53508 16940 58716 16996
rect 58772 16940 58782 16996
rect 200 16884 800 16912
rect 200 16828 1932 16884
rect 1988 16828 1998 16884
rect 18386 16828 18396 16884
rect 18452 16828 19628 16884
rect 19684 16828 19964 16884
rect 20020 16828 20030 16884
rect 20178 16828 20188 16884
rect 20244 16828 21308 16884
rect 21364 16828 21868 16884
rect 21924 16828 21934 16884
rect 22978 16828 22988 16884
rect 23044 16828 25788 16884
rect 25844 16828 25854 16884
rect 28690 16828 28700 16884
rect 28756 16828 29484 16884
rect 29540 16828 30828 16884
rect 30884 16828 30894 16884
rect 32050 16828 32060 16884
rect 32116 16828 33180 16884
rect 33236 16828 33246 16884
rect 33618 16828 33628 16884
rect 33684 16828 33694 16884
rect 34514 16828 34524 16884
rect 34580 16828 34972 16884
rect 35028 16828 35532 16884
rect 35588 16828 35980 16884
rect 36036 16828 36046 16884
rect 36306 16828 36316 16884
rect 36372 16828 36540 16884
rect 36596 16828 36606 16884
rect 36754 16828 36764 16884
rect 36820 16828 39452 16884
rect 39508 16828 39518 16884
rect 40124 16828 41468 16884
rect 41524 16828 41534 16884
rect 42690 16828 42700 16884
rect 42756 16828 43708 16884
rect 43764 16828 43774 16884
rect 45714 16828 45724 16884
rect 45780 16828 46060 16884
rect 46116 16828 46126 16884
rect 47964 16828 55132 16884
rect 55188 16828 55198 16884
rect 56354 16828 56364 16884
rect 56420 16828 56430 16884
rect 56690 16828 56700 16884
rect 56756 16828 57708 16884
rect 57764 16828 58940 16884
rect 58996 16828 59006 16884
rect 200 16800 800 16828
rect 33628 16772 33684 16828
rect 40124 16772 40180 16828
rect 47964 16772 48020 16828
rect 33628 16716 35644 16772
rect 35700 16716 38780 16772
rect 38836 16716 40180 16772
rect 45490 16716 45500 16772
rect 45556 16716 47404 16772
rect 47460 16716 47964 16772
rect 48020 16716 48030 16772
rect 48290 16716 48300 16772
rect 48356 16716 48748 16772
rect 48804 16716 49980 16772
rect 50036 16716 50046 16772
rect 50754 16716 50764 16772
rect 50820 16716 51772 16772
rect 51828 16716 51838 16772
rect 54786 16716 54796 16772
rect 54852 16716 55356 16772
rect 55412 16716 55422 16772
rect 56364 16660 56420 16828
rect 24658 16604 24668 16660
rect 24724 16604 25452 16660
rect 25508 16604 25676 16660
rect 25732 16604 25742 16660
rect 32498 16604 32508 16660
rect 32564 16604 34860 16660
rect 34916 16604 35868 16660
rect 35924 16604 35934 16660
rect 36530 16604 36540 16660
rect 36596 16604 37212 16660
rect 37268 16604 37436 16660
rect 37492 16604 37502 16660
rect 42802 16604 42812 16660
rect 42868 16604 47516 16660
rect 47572 16604 47582 16660
rect 48178 16604 48188 16660
rect 48244 16604 49532 16660
rect 49588 16604 55692 16660
rect 55748 16604 55758 16660
rect 56364 16604 56700 16660
rect 56756 16604 56766 16660
rect 34262 16492 34300 16548
rect 34356 16492 34366 16548
rect 36978 16492 36988 16548
rect 37044 16492 45500 16548
rect 45556 16492 46172 16548
rect 46228 16492 46238 16548
rect 46946 16492 46956 16548
rect 47012 16492 52220 16548
rect 52276 16492 52286 16548
rect 55804 16492 56028 16548
rect 56084 16492 56812 16548
rect 56868 16492 57148 16548
rect 57204 16492 57214 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 42924 16380 44660 16436
rect 42924 16324 42980 16380
rect 44604 16324 44660 16380
rect 46956 16380 49588 16436
rect 49746 16380 49756 16436
rect 49812 16380 55580 16436
rect 55636 16380 55646 16436
rect 46956 16324 47012 16380
rect 49532 16324 49588 16380
rect 14802 16268 14812 16324
rect 14868 16268 15820 16324
rect 15876 16268 16044 16324
rect 16100 16268 16110 16324
rect 36194 16268 36204 16324
rect 36260 16268 36428 16324
rect 36484 16268 36494 16324
rect 42886 16268 42924 16324
rect 42980 16268 42990 16324
rect 43250 16268 43260 16324
rect 43316 16268 44156 16324
rect 44212 16268 44222 16324
rect 44604 16268 47012 16324
rect 47142 16268 47180 16324
rect 47236 16268 47246 16324
rect 48290 16268 48300 16324
rect 48356 16268 48412 16324
rect 48468 16268 48478 16324
rect 49532 16268 50092 16324
rect 50148 16268 50158 16324
rect 50530 16268 50540 16324
rect 50596 16268 51436 16324
rect 51492 16268 51502 16324
rect 51986 16268 51996 16324
rect 52052 16268 52220 16324
rect 52276 16268 52286 16324
rect 53218 16268 53228 16324
rect 53284 16268 54460 16324
rect 54516 16268 54526 16324
rect 55804 16212 55860 16492
rect 19170 16156 19180 16212
rect 19236 16156 19964 16212
rect 20020 16156 21532 16212
rect 21588 16156 21598 16212
rect 23202 16156 23212 16212
rect 23268 16156 24892 16212
rect 24948 16156 36652 16212
rect 36708 16156 36718 16212
rect 42130 16156 42140 16212
rect 42196 16156 43596 16212
rect 43652 16156 43662 16212
rect 46050 16156 46060 16212
rect 46116 16156 49532 16212
rect 49588 16156 49598 16212
rect 50194 16156 50204 16212
rect 50260 16156 55860 16212
rect 16034 16044 16044 16100
rect 16100 16044 17164 16100
rect 17220 16044 17230 16100
rect 23538 16044 23548 16100
rect 23604 16044 24108 16100
rect 24164 16044 24174 16100
rect 31938 16044 31948 16100
rect 32004 16044 33796 16100
rect 37762 16044 37772 16100
rect 37828 16044 38668 16100
rect 38724 16044 38734 16100
rect 39106 16044 39116 16100
rect 39172 16044 39340 16100
rect 39396 16044 39406 16100
rect 41906 16044 41916 16100
rect 41972 16044 43484 16100
rect 43540 16044 45836 16100
rect 45892 16044 45902 16100
rect 46162 16044 46172 16100
rect 46228 16044 48300 16100
rect 48356 16044 48366 16100
rect 48524 16044 49868 16100
rect 49924 16044 49980 16100
rect 50036 16044 50046 16100
rect 51090 16044 51100 16100
rect 51156 16044 51772 16100
rect 51828 16044 51838 16100
rect 54114 16044 54124 16100
rect 54180 16044 56700 16100
rect 56756 16044 56766 16100
rect 33740 15988 33796 16044
rect 41916 15988 41972 16044
rect 48524 15988 48580 16044
rect 14690 15932 14700 15988
rect 14756 15932 16380 15988
rect 16436 15932 16446 15988
rect 28354 15932 28364 15988
rect 28420 15932 29148 15988
rect 29204 15932 29214 15988
rect 33730 15932 33740 15988
rect 33796 15932 34524 15988
rect 34580 15932 34590 15988
rect 36642 15932 36652 15988
rect 36708 15932 37884 15988
rect 37940 15932 41972 15988
rect 44146 15932 44156 15988
rect 44212 15932 45276 15988
rect 45332 15932 47068 15988
rect 47124 15932 47134 15988
rect 48402 15932 48412 15988
rect 48468 15932 48524 15988
rect 48580 15932 48590 15988
rect 49718 15932 49756 15988
rect 49812 15932 49822 15988
rect 50194 15932 50204 15988
rect 50260 15932 51100 15988
rect 51156 15932 51166 15988
rect 53974 15932 54012 15988
rect 54068 15932 54078 15988
rect 55682 15932 55692 15988
rect 55748 15932 56364 15988
rect 56420 15932 56430 15988
rect 56802 15932 56812 15988
rect 56868 15932 57372 15988
rect 57428 15932 57438 15988
rect 56812 15876 56868 15932
rect 14802 15820 14812 15876
rect 14868 15820 17052 15876
rect 17108 15820 17118 15876
rect 18946 15820 18956 15876
rect 19012 15820 20468 15876
rect 32722 15820 32732 15876
rect 32788 15820 35196 15876
rect 35252 15820 35262 15876
rect 36754 15820 36764 15876
rect 36820 15820 41468 15876
rect 41524 15820 41534 15876
rect 42466 15820 42476 15876
rect 42532 15820 42812 15876
rect 42868 15820 42878 15876
rect 46386 15820 46396 15876
rect 46452 15820 46956 15876
rect 47012 15820 47022 15876
rect 47842 15820 47852 15876
rect 47908 15820 51548 15876
rect 51604 15820 51614 15876
rect 53330 15820 53340 15876
rect 53396 15820 55020 15876
rect 55076 15820 55804 15876
rect 55860 15820 55870 15876
rect 55990 15820 56028 15876
rect 56084 15820 56094 15876
rect 56242 15820 56252 15876
rect 56308 15820 56868 15876
rect 20412 15764 20468 15820
rect 16370 15708 16380 15764
rect 16436 15708 18844 15764
rect 18900 15708 18910 15764
rect 20402 15708 20412 15764
rect 20468 15708 21980 15764
rect 22036 15708 37212 15764
rect 37268 15708 37278 15764
rect 40226 15708 40236 15764
rect 40292 15708 42364 15764
rect 42420 15708 50204 15764
rect 50260 15708 50270 15764
rect 51314 15708 51324 15764
rect 51380 15708 51660 15764
rect 51716 15708 51726 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 24098 15596 24108 15652
rect 24164 15596 27132 15652
rect 27188 15596 27198 15652
rect 28466 15596 28476 15652
rect 28532 15596 30044 15652
rect 30100 15596 30110 15652
rect 30370 15596 30380 15652
rect 30436 15596 33740 15652
rect 33796 15596 33806 15652
rect 36866 15596 36876 15652
rect 36932 15596 38220 15652
rect 38276 15596 38286 15652
rect 39106 15596 39116 15652
rect 39172 15596 40236 15652
rect 40292 15596 40348 15652
rect 40404 15596 40414 15652
rect 42018 15596 42028 15652
rect 42084 15596 43260 15652
rect 43316 15596 43326 15652
rect 43670 15596 43708 15652
rect 43764 15596 43774 15652
rect 44258 15596 44268 15652
rect 44324 15596 45052 15652
rect 45108 15596 45118 15652
rect 46946 15596 46956 15652
rect 47012 15596 47404 15652
rect 47460 15596 48076 15652
rect 48132 15596 48142 15652
rect 48738 15596 48748 15652
rect 48804 15596 48860 15652
rect 48916 15596 48926 15652
rect 49074 15596 49084 15652
rect 49140 15596 49644 15652
rect 49700 15596 49710 15652
rect 51538 15596 51548 15652
rect 51604 15596 55020 15652
rect 55076 15596 57260 15652
rect 57316 15596 57326 15652
rect 16146 15484 16156 15540
rect 16212 15484 16828 15540
rect 16884 15484 17612 15540
rect 17668 15484 23772 15540
rect 23828 15484 23838 15540
rect 27458 15484 27468 15540
rect 27524 15484 27916 15540
rect 27972 15484 27982 15540
rect 28242 15484 28252 15540
rect 28308 15484 28700 15540
rect 28756 15484 28766 15540
rect 29586 15484 29596 15540
rect 29652 15484 32620 15540
rect 32676 15484 32686 15540
rect 35970 15484 35980 15540
rect 36036 15484 37100 15540
rect 37156 15484 37166 15540
rect 38098 15484 38108 15540
rect 38164 15484 50596 15540
rect 50540 15428 50596 15484
rect 52668 15484 53676 15540
rect 53732 15484 54572 15540
rect 54628 15484 54638 15540
rect 52668 15428 52724 15484
rect 27122 15372 27132 15428
rect 27188 15372 36708 15428
rect 39554 15372 39564 15428
rect 39620 15372 42476 15428
rect 42532 15372 42542 15428
rect 42774 15372 42812 15428
rect 42868 15372 42878 15428
rect 43586 15372 43596 15428
rect 43652 15372 44604 15428
rect 44660 15372 44670 15428
rect 47506 15372 47516 15428
rect 47572 15372 48412 15428
rect 48468 15372 48636 15428
rect 48692 15372 50428 15428
rect 50540 15372 52668 15428
rect 52724 15372 52734 15428
rect 54422 15372 54460 15428
rect 54516 15372 54526 15428
rect 56662 15372 56700 15428
rect 56756 15372 56766 15428
rect 27906 15260 27916 15316
rect 27972 15260 28364 15316
rect 28420 15260 28430 15316
rect 29138 15260 29148 15316
rect 29204 15260 30380 15316
rect 30436 15260 30446 15316
rect 30604 15260 31948 15316
rect 32004 15260 32014 15316
rect 30604 15204 30660 15260
rect 36652 15204 36708 15372
rect 50372 15316 50428 15372
rect 38210 15260 38220 15316
rect 38276 15260 42980 15316
rect 43698 15260 43708 15316
rect 43764 15260 46172 15316
rect 46228 15260 46238 15316
rect 47170 15260 47180 15316
rect 47236 15260 47246 15316
rect 50372 15260 51548 15316
rect 51604 15260 51614 15316
rect 51762 15260 51772 15316
rect 51828 15260 52556 15316
rect 52612 15260 52622 15316
rect 53218 15260 53228 15316
rect 53284 15260 54236 15316
rect 54292 15260 54302 15316
rect 55794 15260 55804 15316
rect 55860 15260 56364 15316
rect 56420 15260 57484 15316
rect 57540 15260 57550 15316
rect 42924 15204 42980 15260
rect 47180 15204 47236 15260
rect 24434 15148 24444 15204
rect 24500 15148 30660 15204
rect 31826 15148 31836 15204
rect 31892 15148 32284 15204
rect 32340 15148 32844 15204
rect 32900 15148 33292 15204
rect 33348 15148 33358 15204
rect 36642 15148 36652 15204
rect 36708 15148 36718 15204
rect 37090 15148 37100 15204
rect 37156 15148 42476 15204
rect 42532 15148 42700 15204
rect 42756 15148 42766 15204
rect 42924 15148 44268 15204
rect 44324 15148 44334 15204
rect 47180 15148 47404 15204
rect 47460 15148 47470 15204
rect 51426 15148 51436 15204
rect 51492 15148 51502 15204
rect 52770 15148 52780 15204
rect 52836 15148 53340 15204
rect 53396 15148 53452 15204
rect 53508 15148 53676 15204
rect 53732 15148 53742 15204
rect 55654 15148 55692 15204
rect 55748 15148 55758 15204
rect 51436 15092 51492 15148
rect 52098 15092 52108 15148
rect 52164 15092 52174 15148
rect 20514 15036 20524 15092
rect 20580 15036 25676 15092
rect 25732 15036 25742 15092
rect 28802 15036 28812 15092
rect 28868 15036 29596 15092
rect 29652 15036 29662 15092
rect 35186 15036 35196 15092
rect 35252 15036 36876 15092
rect 36932 15036 36942 15092
rect 40674 15036 40684 15092
rect 40740 15036 41468 15092
rect 41524 15036 41534 15092
rect 42466 15036 42476 15092
rect 42532 15036 45724 15092
rect 45780 15036 47740 15092
rect 47796 15036 47806 15092
rect 50194 15036 50204 15092
rect 50260 15036 51492 15092
rect 52108 15036 53172 15092
rect 54114 15036 54124 15092
rect 54180 15036 54796 15092
rect 54852 15036 54862 15092
rect 53116 14980 53172 15036
rect 25554 14924 25564 14980
rect 25620 14924 26236 14980
rect 26292 14924 26302 14980
rect 40114 14924 40124 14980
rect 40180 14924 40190 14980
rect 41570 14924 41580 14980
rect 41636 14924 41916 14980
rect 41972 14924 41982 14980
rect 43474 14924 43484 14980
rect 43540 14924 43820 14980
rect 43876 14924 43886 14980
rect 44034 14924 44044 14980
rect 44100 14924 44604 14980
rect 44660 14924 44670 14980
rect 48962 14924 48972 14980
rect 49028 14924 50316 14980
rect 50372 14924 52108 14980
rect 52164 14924 52174 14980
rect 52322 14924 52332 14980
rect 52388 14924 52398 14980
rect 53106 14924 53116 14980
rect 53172 14924 53182 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 30930 14812 30940 14868
rect 30996 14812 33180 14868
rect 33236 14812 33246 14868
rect 14242 14700 14252 14756
rect 14308 14700 14924 14756
rect 14980 14700 16156 14756
rect 16212 14700 16222 14756
rect 18946 14700 18956 14756
rect 19012 14700 20524 14756
rect 20580 14700 20590 14756
rect 40124 14644 40180 14924
rect 41916 14868 41972 14924
rect 52332 14868 52388 14924
rect 41916 14812 50988 14868
rect 51044 14812 51054 14868
rect 52332 14812 53788 14868
rect 53844 14812 53854 14868
rect 41682 14700 41692 14756
rect 41748 14700 41916 14756
rect 41972 14700 41982 14756
rect 43250 14700 43260 14756
rect 43316 14700 45948 14756
rect 46004 14700 47964 14756
rect 48020 14700 48030 14756
rect 48850 14700 48860 14756
rect 48916 14700 51324 14756
rect 51380 14700 51390 14756
rect 52294 14700 52332 14756
rect 52388 14700 52398 14756
rect 20290 14588 20300 14644
rect 20356 14588 21532 14644
rect 21588 14588 21598 14644
rect 28242 14588 28252 14644
rect 28308 14588 28700 14644
rect 28756 14588 28766 14644
rect 32050 14588 32060 14644
rect 32116 14588 32732 14644
rect 32788 14588 39900 14644
rect 39956 14588 39966 14644
rect 40124 14588 41580 14644
rect 41636 14588 48972 14644
rect 49028 14588 49038 14644
rect 50166 14588 50204 14644
rect 50260 14588 50270 14644
rect 50372 14588 51436 14644
rect 51492 14588 58044 14644
rect 58100 14588 58110 14644
rect 50372 14532 50428 14588
rect 14466 14476 14476 14532
rect 14532 14476 17108 14532
rect 20626 14476 20636 14532
rect 20692 14476 22316 14532
rect 22372 14476 22382 14532
rect 22642 14476 22652 14532
rect 22708 14476 24220 14532
rect 24276 14476 24286 14532
rect 25778 14476 25788 14532
rect 25844 14476 26796 14532
rect 26852 14476 26862 14532
rect 27346 14476 27356 14532
rect 27412 14476 29484 14532
rect 29540 14476 29550 14532
rect 31938 14476 31948 14532
rect 32004 14476 35308 14532
rect 35364 14476 35374 14532
rect 35532 14476 38668 14532
rect 39190 14476 39228 14532
rect 39284 14476 39294 14532
rect 40786 14476 40796 14532
rect 40852 14476 41692 14532
rect 41748 14476 41758 14532
rect 43110 14476 43148 14532
rect 43204 14476 43214 14532
rect 44818 14476 44828 14532
rect 44884 14476 49364 14532
rect 50082 14476 50092 14532
rect 50148 14476 50428 14532
rect 50530 14476 50540 14532
rect 50596 14476 51212 14532
rect 51268 14476 51548 14532
rect 51604 14476 51614 14532
rect 54674 14476 54684 14532
rect 54740 14476 55020 14532
rect 55076 14476 55086 14532
rect 17052 14420 17108 14476
rect 35532 14420 35588 14476
rect 13794 14364 13804 14420
rect 13860 14364 14700 14420
rect 14756 14364 15932 14420
rect 15988 14364 16660 14420
rect 17042 14364 17052 14420
rect 17108 14364 20188 14420
rect 24098 14364 24108 14420
rect 24164 14364 31052 14420
rect 31108 14364 31118 14420
rect 31276 14364 35588 14420
rect 35746 14364 35756 14420
rect 35812 14364 38444 14420
rect 38500 14364 38510 14420
rect 16604 14308 16660 14364
rect 20132 14308 20188 14364
rect 31276 14308 31332 14364
rect 6962 14252 6972 14308
rect 7028 14252 13020 14308
rect 13076 14252 13086 14308
rect 14914 14252 14924 14308
rect 14980 14252 16044 14308
rect 16100 14252 16110 14308
rect 16594 14252 16604 14308
rect 16660 14252 17948 14308
rect 18004 14252 18014 14308
rect 20132 14252 26124 14308
rect 26180 14252 26190 14308
rect 26674 14252 26684 14308
rect 26740 14252 27468 14308
rect 27524 14252 29820 14308
rect 29876 14252 30268 14308
rect 30324 14252 30492 14308
rect 30548 14252 31332 14308
rect 32722 14252 32732 14308
rect 32788 14252 33292 14308
rect 33348 14252 33358 14308
rect 33954 14252 33964 14308
rect 34020 14252 36316 14308
rect 36372 14252 36988 14308
rect 37044 14252 37548 14308
rect 37604 14252 37614 14308
rect 38612 14196 38668 14476
rect 49308 14420 49364 14476
rect 40674 14364 40684 14420
rect 40740 14364 44268 14420
rect 44324 14364 45500 14420
rect 45556 14364 45566 14420
rect 45714 14364 45724 14420
rect 45780 14364 45790 14420
rect 47058 14364 47068 14420
rect 47124 14364 47740 14420
rect 47796 14364 47806 14420
rect 49298 14364 49308 14420
rect 49364 14364 51996 14420
rect 52052 14364 52062 14420
rect 52882 14364 52892 14420
rect 52948 14364 54124 14420
rect 54180 14364 54190 14420
rect 55122 14364 55132 14420
rect 55188 14364 56140 14420
rect 56196 14364 57148 14420
rect 57204 14364 57214 14420
rect 38882 14252 38892 14308
rect 38948 14252 39564 14308
rect 39620 14252 39630 14308
rect 41346 14252 41356 14308
rect 41412 14252 45388 14308
rect 45444 14252 45454 14308
rect 45724 14196 45780 14364
rect 46162 14252 46172 14308
rect 46228 14252 46732 14308
rect 46788 14252 46798 14308
rect 47170 14252 47180 14308
rect 47236 14252 48188 14308
rect 48244 14252 52556 14308
rect 52612 14252 53228 14308
rect 53284 14252 53294 14308
rect 53554 14252 53564 14308
rect 53620 14252 54348 14308
rect 54404 14252 54414 14308
rect 54786 14252 54796 14308
rect 54852 14252 55356 14308
rect 55412 14252 57036 14308
rect 57092 14252 57102 14308
rect 35858 14140 35868 14196
rect 35924 14140 35934 14196
rect 38612 14140 38780 14196
rect 38836 14140 38846 14196
rect 40002 14140 40012 14196
rect 40068 14140 41468 14196
rect 41524 14140 41534 14196
rect 44482 14140 44492 14196
rect 44548 14140 45164 14196
rect 45220 14140 45230 14196
rect 45490 14140 45500 14196
rect 45556 14140 45780 14196
rect 47058 14140 47068 14196
rect 47124 14140 47964 14196
rect 48020 14140 48972 14196
rect 49028 14140 49038 14196
rect 51426 14140 51436 14196
rect 51492 14140 51548 14196
rect 51604 14140 51614 14196
rect 52406 14140 52444 14196
rect 52500 14140 53340 14196
rect 53396 14140 55580 14196
rect 55636 14140 55646 14196
rect 56690 14140 56700 14196
rect 56756 14140 57484 14196
rect 57540 14140 57550 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 35868 14084 35924 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 24770 14028 24780 14084
rect 24836 14028 25340 14084
rect 25396 14028 25564 14084
rect 25620 14028 25630 14084
rect 35756 14028 42140 14084
rect 42196 14028 42206 14084
rect 42364 14028 46508 14084
rect 46564 14028 46574 14084
rect 51874 14028 51884 14084
rect 51940 14028 53564 14084
rect 53620 14028 53630 14084
rect 54450 14028 54460 14084
rect 54516 14028 55132 14084
rect 55188 14028 55468 14084
rect 55524 14028 57932 14084
rect 57988 14028 57998 14084
rect 13906 13916 13916 13972
rect 13972 13916 14476 13972
rect 14532 13916 14542 13972
rect 15362 13916 15372 13972
rect 15428 13916 16492 13972
rect 16548 13916 16558 13972
rect 22306 13916 22316 13972
rect 22372 13916 22988 13972
rect 23044 13916 23436 13972
rect 23492 13916 23502 13972
rect 24546 13916 24556 13972
rect 24612 13916 25452 13972
rect 25508 13916 26012 13972
rect 26068 13916 26078 13972
rect 26226 13916 26236 13972
rect 26292 13916 27804 13972
rect 27860 13916 27870 13972
rect 34738 13916 34748 13972
rect 34804 13916 35196 13972
rect 35252 13916 35262 13972
rect 15474 13804 15484 13860
rect 15540 13804 16716 13860
rect 16772 13804 16782 13860
rect 26852 13804 34860 13860
rect 34916 13804 34926 13860
rect 26852 13748 26908 13804
rect 35756 13748 35812 14028
rect 42364 13972 42420 14028
rect 38658 13916 38668 13972
rect 38724 13916 39004 13972
rect 39060 13916 40236 13972
rect 40292 13916 40302 13972
rect 40572 13916 41356 13972
rect 41412 13916 42420 13972
rect 42914 13916 42924 13972
rect 42980 13916 43260 13972
rect 43316 13916 43932 13972
rect 43988 13916 47404 13972
rect 47460 13916 47470 13972
rect 47730 13916 47740 13972
rect 47796 13916 50316 13972
rect 50372 13916 51100 13972
rect 51156 13916 52444 13972
rect 52500 13916 52510 13972
rect 39666 13804 39676 13860
rect 39732 13804 40348 13860
rect 40404 13804 40414 13860
rect 40572 13748 40628 13916
rect 14690 13692 14700 13748
rect 14756 13692 15036 13748
rect 15092 13692 15260 13748
rect 15316 13692 15326 13748
rect 17938 13692 17948 13748
rect 18004 13692 26908 13748
rect 27010 13692 27020 13748
rect 27076 13692 27804 13748
rect 27860 13692 27870 13748
rect 28466 13692 28476 13748
rect 28532 13692 28812 13748
rect 28868 13692 30268 13748
rect 30324 13692 30334 13748
rect 35746 13692 35756 13748
rect 35812 13692 35822 13748
rect 36530 13692 36540 13748
rect 36596 13692 38108 13748
rect 38164 13692 38174 13748
rect 39824 13692 39900 13748
rect 39956 13692 40628 13748
rect 40796 13804 41916 13860
rect 41972 13804 42812 13860
rect 42868 13804 42878 13860
rect 43708 13804 44268 13860
rect 44324 13804 44334 13860
rect 46722 13804 46732 13860
rect 46788 13804 46956 13860
rect 47012 13804 47022 13860
rect 48850 13804 48860 13860
rect 48916 13804 49980 13860
rect 50036 13804 50046 13860
rect 53442 13804 53452 13860
rect 53508 13804 55356 13860
rect 55412 13804 55422 13860
rect 55580 13804 56364 13860
rect 56420 13804 56430 13860
rect 57698 13804 57708 13860
rect 57764 13804 58044 13860
rect 58100 13804 58110 13860
rect 40796 13636 40852 13804
rect 42476 13748 42532 13804
rect 43708 13748 43764 13804
rect 55580 13748 55636 13804
rect 41010 13692 41020 13748
rect 41076 13692 41804 13748
rect 41860 13692 41870 13748
rect 42466 13692 42476 13748
rect 42532 13692 42542 13748
rect 42914 13692 42924 13748
rect 42980 13692 43484 13748
rect 43540 13692 43550 13748
rect 43698 13692 43708 13748
rect 43764 13692 43774 13748
rect 46498 13692 46508 13748
rect 46564 13692 47068 13748
rect 47124 13692 47134 13748
rect 48402 13692 48412 13748
rect 48468 13692 49420 13748
rect 49476 13692 51884 13748
rect 51940 13692 51950 13748
rect 52210 13692 52220 13748
rect 52276 13692 55636 13748
rect 56466 13692 56476 13748
rect 56532 13692 57372 13748
rect 57428 13692 57438 13748
rect 20850 13580 20860 13636
rect 20916 13580 21980 13636
rect 22036 13580 23436 13636
rect 23492 13580 23502 13636
rect 24882 13580 24892 13636
rect 24948 13580 25676 13636
rect 25732 13580 28700 13636
rect 28756 13580 29260 13636
rect 29316 13580 29326 13636
rect 35410 13580 35420 13636
rect 35476 13580 36204 13636
rect 36260 13580 36270 13636
rect 39218 13580 39228 13636
rect 39284 13580 40852 13636
rect 41458 13580 41468 13636
rect 41524 13580 42252 13636
rect 42308 13580 42318 13636
rect 42690 13580 42700 13636
rect 42756 13580 43932 13636
rect 43988 13580 46172 13636
rect 46228 13580 46238 13636
rect 47394 13580 47404 13636
rect 47460 13580 48188 13636
rect 48244 13580 48254 13636
rect 49298 13580 49308 13636
rect 49364 13580 50988 13636
rect 51044 13580 51054 13636
rect 53778 13580 53788 13636
rect 53844 13580 54236 13636
rect 54292 13580 54460 13636
rect 54516 13580 54526 13636
rect 55570 13580 55580 13636
rect 55636 13580 56588 13636
rect 56644 13580 56654 13636
rect 39676 13524 39732 13580
rect 15922 13468 15932 13524
rect 15988 13468 16828 13524
rect 16884 13468 16894 13524
rect 29698 13468 29708 13524
rect 29764 13468 31500 13524
rect 31556 13468 31566 13524
rect 39666 13468 39676 13524
rect 39732 13468 39742 13524
rect 40646 13468 40684 13524
rect 40740 13468 40750 13524
rect 41234 13468 41244 13524
rect 41300 13468 42924 13524
rect 42980 13468 42990 13524
rect 45686 13468 45724 13524
rect 45780 13468 45790 13524
rect 46722 13468 46732 13524
rect 46788 13468 47964 13524
rect 48020 13468 48300 13524
rect 48356 13468 48366 13524
rect 50418 13468 50428 13524
rect 50484 13468 50988 13524
rect 51044 13468 51054 13524
rect 51762 13468 51772 13524
rect 51828 13468 52556 13524
rect 52612 13468 54124 13524
rect 54180 13468 55020 13524
rect 55076 13468 55086 13524
rect 55570 13468 55580 13524
rect 55636 13468 55916 13524
rect 55972 13468 55982 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 16492 13300 16548 13468
rect 25666 13356 25676 13412
rect 25732 13356 26348 13412
rect 26404 13356 26414 13412
rect 31826 13356 31836 13412
rect 31892 13356 32396 13412
rect 32452 13356 32462 13412
rect 39442 13356 39452 13412
rect 39508 13356 40348 13412
rect 40404 13356 40414 13412
rect 41542 13356 41580 13412
rect 41636 13356 41646 13412
rect 52182 13356 52220 13412
rect 52276 13356 52286 13412
rect 54002 13356 54012 13412
rect 54068 13356 54796 13412
rect 54852 13356 54862 13412
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 41580 13300 41636 13356
rect 16482 13244 16492 13300
rect 16548 13244 16558 13300
rect 39218 13244 39228 13300
rect 39284 13244 41636 13300
rect 43474 13244 43484 13300
rect 43540 13244 44156 13300
rect 44212 13244 44222 13300
rect 50306 13244 50316 13300
rect 50372 13244 53900 13300
rect 53956 13244 53966 13300
rect 14354 13132 14364 13188
rect 14420 13132 15260 13188
rect 15316 13132 15326 13188
rect 36866 13132 36876 13188
rect 36932 13132 51100 13188
rect 51156 13132 51166 13188
rect 51436 13132 59388 13188
rect 59444 13132 59454 13188
rect 51436 13076 51492 13132
rect 19842 13020 19852 13076
rect 19908 13020 20860 13076
rect 20916 13020 21196 13076
rect 21252 13020 21262 13076
rect 28578 13020 28588 13076
rect 28644 13020 29596 13076
rect 29652 13020 29662 13076
rect 39414 13020 39452 13076
rect 39508 13020 39518 13076
rect 39778 13020 39788 13076
rect 39844 13020 40572 13076
rect 40628 13020 40638 13076
rect 42018 13020 42028 13076
rect 42084 13020 42924 13076
rect 42980 13020 42990 13076
rect 45938 13020 45948 13076
rect 46004 13020 46060 13076
rect 46116 13020 46126 13076
rect 51090 13020 51100 13076
rect 51156 13020 51492 13076
rect 51762 13020 51772 13076
rect 51828 13020 52668 13076
rect 52724 13020 52734 13076
rect 54870 13020 54908 13076
rect 54964 13020 54974 13076
rect 55728 13020 55804 13076
rect 55860 13020 57260 13076
rect 57316 13020 57326 13076
rect 24658 12908 24668 12964
rect 24724 12908 24892 12964
rect 24948 12908 25116 12964
rect 25172 12908 25900 12964
rect 25956 12908 25966 12964
rect 29698 12908 29708 12964
rect 29764 12908 29774 12964
rect 32946 12908 32956 12964
rect 33012 12908 33964 12964
rect 34020 12908 37996 12964
rect 38052 12908 38062 12964
rect 38434 12908 38444 12964
rect 38500 12908 39340 12964
rect 39396 12908 39406 12964
rect 42130 12908 42140 12964
rect 42196 12908 46508 12964
rect 46564 12908 46574 12964
rect 48066 12908 48076 12964
rect 48132 12908 49644 12964
rect 49700 12908 49710 12964
rect 49858 12908 49868 12964
rect 49924 12908 55020 12964
rect 55076 12908 55086 12964
rect 56802 12908 56812 12964
rect 56868 12908 57036 12964
rect 57092 12908 57102 12964
rect 29708 12852 29764 12908
rect 19954 12796 19964 12852
rect 20020 12796 20524 12852
rect 20580 12796 20590 12852
rect 28802 12796 28812 12852
rect 28868 12796 29764 12852
rect 31490 12796 31500 12852
rect 31556 12796 32620 12852
rect 32676 12796 32686 12852
rect 33170 12796 33180 12852
rect 33236 12796 33852 12852
rect 33908 12796 39116 12852
rect 39172 12796 39182 12852
rect 44118 12796 44156 12852
rect 44212 12796 44222 12852
rect 44370 12796 44380 12852
rect 44436 12796 45836 12852
rect 45892 12796 51996 12852
rect 52052 12796 52062 12852
rect 53414 12796 53452 12852
rect 53508 12796 53518 12852
rect 54226 12796 54236 12852
rect 54292 12796 54684 12852
rect 54740 12796 54908 12852
rect 54964 12796 54974 12852
rect 18498 12684 18508 12740
rect 18564 12684 19068 12740
rect 19124 12684 19134 12740
rect 28578 12684 28588 12740
rect 28644 12684 29260 12740
rect 29316 12684 29708 12740
rect 29764 12684 30940 12740
rect 30996 12684 31006 12740
rect 40338 12684 40348 12740
rect 40404 12684 41916 12740
rect 41972 12684 51884 12740
rect 51940 12684 51950 12740
rect 52546 12684 52556 12740
rect 52612 12684 53004 12740
rect 53060 12684 53070 12740
rect 53218 12684 53228 12740
rect 53284 12684 53676 12740
rect 53732 12684 53742 12740
rect 57698 12684 57708 12740
rect 57764 12684 57988 12740
rect 20514 12572 20524 12628
rect 20580 12572 21196 12628
rect 21252 12572 21868 12628
rect 21924 12572 36652 12628
rect 36708 12572 36718 12628
rect 39078 12572 39116 12628
rect 39172 12572 39182 12628
rect 44706 12572 44716 12628
rect 44772 12572 45276 12628
rect 45332 12572 45342 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 49532 12516 49588 12684
rect 57932 12628 57988 12684
rect 50978 12572 50988 12628
rect 51044 12572 51436 12628
rect 51492 12572 51502 12628
rect 51650 12572 51660 12628
rect 51716 12572 56812 12628
rect 56868 12572 56878 12628
rect 57922 12572 57932 12628
rect 57988 12572 57998 12628
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 26338 12460 26348 12516
rect 26404 12460 26572 12516
rect 26628 12460 31164 12516
rect 31220 12460 31230 12516
rect 42662 12460 42700 12516
rect 42756 12460 42766 12516
rect 45154 12460 45164 12516
rect 45220 12460 47516 12516
rect 47572 12460 47582 12516
rect 49522 12460 49532 12516
rect 49588 12460 49598 12516
rect 50988 12460 54236 12516
rect 54292 12460 54302 12516
rect 57110 12460 57148 12516
rect 57204 12460 57214 12516
rect 50988 12404 51044 12460
rect 2706 12348 2716 12404
rect 2772 12348 3724 12404
rect 3780 12348 3790 12404
rect 15474 12348 15484 12404
rect 15540 12348 15550 12404
rect 34738 12348 34748 12404
rect 34804 12348 35084 12404
rect 35140 12348 35532 12404
rect 35588 12348 35598 12404
rect 35858 12348 35868 12404
rect 35924 12348 36764 12404
rect 36820 12348 36830 12404
rect 50754 12348 50764 12404
rect 50820 12348 51044 12404
rect 51202 12348 51212 12404
rect 51268 12348 54684 12404
rect 54740 12348 54750 12404
rect 56018 12348 56028 12404
rect 56084 12348 58156 12404
rect 58212 12348 58940 12404
rect 58996 12348 59006 12404
rect 15484 12180 15540 12348
rect 36418 12236 36428 12292
rect 36484 12236 37100 12292
rect 37156 12236 37166 12292
rect 40562 12236 40572 12292
rect 40628 12236 42644 12292
rect 44482 12236 44492 12292
rect 44548 12236 46172 12292
rect 46228 12236 46238 12292
rect 47058 12236 47068 12292
rect 47124 12236 49868 12292
rect 49924 12236 49934 12292
rect 50082 12236 50092 12292
rect 50148 12236 50988 12292
rect 51044 12236 51660 12292
rect 51716 12236 51996 12292
rect 52052 12236 52062 12292
rect 42588 12180 42644 12236
rect 15484 12124 15708 12180
rect 15764 12124 21980 12180
rect 22036 12124 22046 12180
rect 30370 12124 30380 12180
rect 30436 12124 31276 12180
rect 31332 12124 31342 12180
rect 31826 12124 31836 12180
rect 31892 12124 32508 12180
rect 32564 12124 32574 12180
rect 36194 12124 36204 12180
rect 36260 12124 37212 12180
rect 37268 12124 37278 12180
rect 37874 12124 37884 12180
rect 37940 12124 38780 12180
rect 38836 12124 42364 12180
rect 42420 12124 42430 12180
rect 42588 12124 49420 12180
rect 49476 12124 49486 12180
rect 51202 12124 51212 12180
rect 51268 12124 51324 12180
rect 51380 12124 51390 12180
rect 51734 12124 51772 12180
rect 51828 12124 51838 12180
rect 2482 12012 2492 12068
rect 2548 12012 3164 12068
rect 3220 12012 14252 12068
rect 14308 12012 14318 12068
rect 18946 12012 18956 12068
rect 19012 12012 19404 12068
rect 19460 12012 20300 12068
rect 20356 12012 20366 12068
rect 29922 12012 29932 12068
rect 29988 12012 30492 12068
rect 30548 12012 30558 12068
rect 31042 12012 31052 12068
rect 31108 12012 33516 12068
rect 33572 12012 42700 12068
rect 42756 12012 42766 12068
rect 45938 12012 45948 12068
rect 46004 12012 46508 12068
rect 46564 12012 46574 12068
rect 47478 12012 47516 12068
rect 47572 12012 47582 12068
rect 48150 12012 48188 12068
rect 48244 12012 48254 12068
rect 50372 12012 50764 12068
rect 50820 12012 50830 12068
rect 51314 12012 51324 12068
rect 51380 12012 51436 12068
rect 51492 12012 52668 12068
rect 52724 12012 52734 12068
rect 45948 11956 46004 12012
rect 50372 11956 50428 12012
rect 53116 11956 53172 12348
rect 53442 12236 53452 12292
rect 53508 12236 53676 12292
rect 53732 12236 53742 12292
rect 54226 12236 54236 12292
rect 54292 12236 55356 12292
rect 55412 12236 58044 12292
rect 58100 12236 58110 12292
rect 59200 12180 59800 12208
rect 53554 12124 53564 12180
rect 53620 12124 53900 12180
rect 53956 12124 53966 12180
rect 56130 12124 56140 12180
rect 56196 12124 59800 12180
rect 59200 12096 59800 12124
rect 53414 12012 53452 12068
rect 53508 12012 53518 12068
rect 55682 12012 55692 12068
rect 55748 12012 57036 12068
rect 57092 12012 57820 12068
rect 57876 12012 57886 12068
rect 19058 11900 19068 11956
rect 19124 11900 19516 11956
rect 19572 11900 20524 11956
rect 20580 11900 27356 11956
rect 27412 11900 27422 11956
rect 30930 11900 30940 11956
rect 30996 11900 32620 11956
rect 32676 11900 33964 11956
rect 34020 11900 34188 11956
rect 34244 11900 35588 11956
rect 36082 11900 36092 11956
rect 36148 11900 37324 11956
rect 37380 11900 37390 11956
rect 40674 11900 40684 11956
rect 40740 11900 46004 11956
rect 46386 11900 46396 11956
rect 46452 11900 50428 11956
rect 50876 11900 51940 11956
rect 53106 11900 53116 11956
rect 53172 11900 53182 11956
rect 53452 11900 54908 11956
rect 54964 11900 54974 11956
rect 35532 11844 35588 11900
rect 50876 11844 50932 11900
rect 51884 11844 51940 11900
rect 53452 11844 53508 11900
rect 23202 11788 23212 11844
rect 23268 11788 23772 11844
rect 23828 11788 23838 11844
rect 32498 11788 32508 11844
rect 32564 11788 33628 11844
rect 33684 11788 33694 11844
rect 35532 11788 37548 11844
rect 37604 11788 37614 11844
rect 38546 11788 38556 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 23426 11676 23436 11732
rect 23492 11676 31836 11732
rect 31892 11676 31902 11732
rect 38612 11676 38668 11844
rect 44146 11788 44156 11844
rect 44212 11788 44222 11844
rect 44482 11788 44492 11844
rect 44548 11788 45164 11844
rect 45220 11788 45230 11844
rect 45826 11788 45836 11844
rect 45892 11788 46284 11844
rect 46340 11788 46350 11844
rect 49410 11788 49420 11844
rect 49476 11788 50932 11844
rect 51090 11788 51100 11844
rect 51156 11788 51660 11844
rect 51716 11788 51726 11844
rect 51884 11788 53508 11844
rect 53666 11788 53676 11844
rect 53732 11788 54180 11844
rect 54450 11788 54460 11844
rect 54516 11788 57708 11844
rect 57764 11788 57774 11844
rect 44156 11732 44212 11788
rect 51660 11732 51716 11788
rect 54124 11732 54180 11788
rect 38724 11676 38734 11732
rect 38882 11676 38892 11732
rect 38948 11676 44268 11732
rect 44324 11676 44334 11732
rect 45042 11676 45052 11732
rect 45108 11676 45724 11732
rect 45780 11676 46844 11732
rect 46900 11676 46910 11732
rect 51660 11676 52444 11732
rect 52500 11676 52510 11732
rect 54114 11676 54124 11732
rect 54180 11676 54190 11732
rect 26114 11564 26124 11620
rect 26180 11564 32060 11620
rect 32116 11564 32126 11620
rect 43138 11564 43148 11620
rect 43204 11564 44156 11620
rect 44212 11564 44222 11620
rect 44370 11564 44380 11620
rect 44436 11564 44940 11620
rect 44996 11564 45006 11620
rect 50306 11564 50316 11620
rect 50372 11564 51660 11620
rect 51716 11564 51726 11620
rect 51874 11564 51884 11620
rect 51940 11564 52220 11620
rect 52276 11564 52286 11620
rect 53778 11564 53788 11620
rect 53844 11564 54460 11620
rect 54516 11564 55020 11620
rect 55076 11564 57932 11620
rect 57988 11564 57998 11620
rect 44380 11508 44436 11564
rect 43250 11452 43260 11508
rect 43316 11452 44436 11508
rect 48290 11452 48300 11508
rect 48356 11452 48748 11508
rect 48804 11452 48814 11508
rect 49158 11452 49196 11508
rect 49252 11452 49262 11508
rect 49644 11452 51100 11508
rect 51156 11452 51166 11508
rect 55122 11452 55132 11508
rect 55188 11452 56476 11508
rect 56532 11452 56542 11508
rect 57362 11452 57372 11508
rect 57428 11452 58380 11508
rect 58436 11452 58446 11508
rect 49644 11396 49700 11452
rect 15138 11340 15148 11396
rect 15204 11340 15708 11396
rect 15764 11340 15774 11396
rect 19282 11340 19292 11396
rect 19348 11340 19740 11396
rect 19796 11340 19806 11396
rect 22866 11340 22876 11396
rect 22932 11340 23996 11396
rect 24052 11340 24062 11396
rect 30594 11340 30604 11396
rect 30660 11340 31052 11396
rect 31108 11340 31948 11396
rect 32004 11340 33628 11396
rect 33684 11340 44044 11396
rect 44100 11340 44110 11396
rect 47170 11340 47180 11396
rect 47236 11340 47852 11396
rect 47908 11340 47918 11396
rect 48738 11340 48748 11396
rect 48804 11340 49700 11396
rect 50194 11340 50204 11396
rect 50260 11340 50652 11396
rect 50708 11340 51548 11396
rect 51604 11340 53788 11396
rect 53844 11340 53854 11396
rect 47180 11284 47236 11340
rect 17266 11228 17276 11284
rect 17332 11228 30380 11284
rect 30436 11228 30446 11284
rect 32162 11228 32172 11284
rect 32228 11228 32396 11284
rect 32452 11228 32462 11284
rect 34850 11228 34860 11284
rect 34916 11228 35084 11284
rect 35140 11228 35980 11284
rect 36036 11228 36046 11284
rect 40786 11228 40796 11284
rect 40852 11228 41468 11284
rect 41524 11228 42196 11284
rect 42914 11228 42924 11284
rect 42980 11228 43596 11284
rect 43652 11228 43662 11284
rect 43922 11228 43932 11284
rect 43988 11228 45276 11284
rect 45332 11228 47236 11284
rect 48738 11228 48748 11284
rect 48804 11228 49980 11284
rect 50036 11228 50046 11284
rect 50306 11228 50316 11284
rect 50372 11228 50876 11284
rect 50932 11228 51212 11284
rect 51268 11228 51278 11284
rect 52882 11228 52892 11284
rect 52948 11228 53228 11284
rect 53284 11228 53294 11284
rect 30482 11116 30492 11172
rect 30548 11116 31276 11172
rect 31332 11116 31724 11172
rect 31780 11116 33180 11172
rect 33236 11116 33246 11172
rect 36530 11116 36540 11172
rect 36596 11116 41916 11172
rect 41972 11116 41982 11172
rect 42140 11060 42196 11228
rect 42690 11116 42700 11172
rect 42756 11116 45388 11172
rect 45444 11116 46844 11172
rect 46900 11116 46910 11172
rect 49606 11116 49644 11172
rect 49700 11116 49710 11172
rect 50372 11116 50764 11172
rect 50820 11116 51044 11172
rect 52546 11116 52556 11172
rect 52612 11116 53564 11172
rect 53620 11116 53900 11172
rect 53956 11116 53966 11172
rect 50372 11060 50428 11116
rect 40226 11004 40236 11060
rect 40292 11004 41692 11060
rect 41748 11004 41758 11060
rect 42018 11004 42028 11060
rect 42084 11004 42196 11060
rect 44258 11004 44268 11060
rect 44324 11004 45724 11060
rect 45780 11004 45790 11060
rect 46844 11004 50428 11060
rect 50988 11060 51044 11116
rect 50988 11004 54684 11060
rect 54740 11004 54750 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 36306 10892 36316 10948
rect 36372 10892 37100 10948
rect 37156 10892 38668 10948
rect 38724 10892 46620 10948
rect 46676 10892 46686 10948
rect 200 10836 800 10864
rect 46844 10836 46900 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 49074 10892 49084 10948
rect 49140 10892 50428 10948
rect 52770 10892 52780 10948
rect 52836 10892 56476 10948
rect 56532 10892 56542 10948
rect 50372 10836 50428 10892
rect 200 10780 1932 10836
rect 1988 10780 1998 10836
rect 2706 10780 2716 10836
rect 2772 10780 3276 10836
rect 3332 10780 10668 10836
rect 10724 10780 10734 10836
rect 14802 10780 14812 10836
rect 14868 10780 15820 10836
rect 15876 10780 15886 10836
rect 22642 10780 22652 10836
rect 22708 10780 24108 10836
rect 24164 10780 28364 10836
rect 28420 10780 28430 10836
rect 42018 10780 42028 10836
rect 42084 10780 42094 10836
rect 42354 10780 42364 10836
rect 42420 10780 46060 10836
rect 46116 10780 46900 10836
rect 49494 10780 49532 10836
rect 49588 10780 49598 10836
rect 50372 10780 54572 10836
rect 54628 10780 54638 10836
rect 57026 10780 57036 10836
rect 57092 10780 57820 10836
rect 57876 10780 57886 10836
rect 200 10752 800 10780
rect 16258 10668 16268 10724
rect 16324 10668 16828 10724
rect 16884 10668 18060 10724
rect 18116 10668 18126 10724
rect 20132 10668 23996 10724
rect 24052 10668 24062 10724
rect 26450 10668 26460 10724
rect 26516 10668 27580 10724
rect 27636 10668 27646 10724
rect 29922 10668 29932 10724
rect 29988 10668 30492 10724
rect 30548 10668 30558 10724
rect 33170 10668 33180 10724
rect 33236 10668 38668 10724
rect 38724 10668 38734 10724
rect 20132 10612 20188 10668
rect 16482 10556 16492 10612
rect 16548 10556 16940 10612
rect 16996 10556 17724 10612
rect 17780 10556 20188 10612
rect 24994 10556 25004 10612
rect 25060 10556 25900 10612
rect 25956 10556 26684 10612
rect 26740 10556 26750 10612
rect 31154 10556 31164 10612
rect 31220 10556 32060 10612
rect 32116 10556 32126 10612
rect 34178 10556 34188 10612
rect 34244 10556 34254 10612
rect 39442 10556 39452 10612
rect 39508 10556 40236 10612
rect 40292 10556 40302 10612
rect 34188 10500 34244 10556
rect 15026 10444 15036 10500
rect 15092 10444 16156 10500
rect 16212 10444 16716 10500
rect 16772 10444 16782 10500
rect 17602 10444 17612 10500
rect 17668 10444 18284 10500
rect 18340 10444 19292 10500
rect 19348 10444 19358 10500
rect 33730 10444 33740 10500
rect 33796 10444 34244 10500
rect 42028 10500 42084 10780
rect 45714 10668 45724 10724
rect 45780 10668 45948 10724
rect 46004 10668 46014 10724
rect 49970 10668 49980 10724
rect 50036 10668 51100 10724
rect 51156 10668 51166 10724
rect 52770 10668 52780 10724
rect 52836 10668 53340 10724
rect 53396 10668 53406 10724
rect 49074 10556 49084 10612
rect 49140 10556 49980 10612
rect 50036 10556 56364 10612
rect 56420 10556 56430 10612
rect 42028 10444 49756 10500
rect 49812 10444 49980 10500
rect 50036 10444 50046 10500
rect 54562 10444 54572 10500
rect 54628 10444 55020 10500
rect 55076 10444 56028 10500
rect 56084 10444 56094 10500
rect 25554 10332 25564 10388
rect 25620 10332 26236 10388
rect 26292 10332 27244 10388
rect 27300 10332 27310 10388
rect 50978 10332 50988 10388
rect 51044 10332 51268 10388
rect 51212 10276 51268 10332
rect 25218 10220 25228 10276
rect 25284 10220 25294 10276
rect 25554 10220 25564 10276
rect 25620 10220 25788 10276
rect 25844 10220 25854 10276
rect 38658 10220 38668 10276
rect 38724 10220 44492 10276
rect 44548 10220 44558 10276
rect 51212 10220 54012 10276
rect 54068 10220 54078 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 25228 10052 25284 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 25442 10108 25452 10164
rect 25508 10108 34412 10164
rect 34468 10108 34478 10164
rect 48598 10108 48636 10164
rect 48692 10108 48702 10164
rect 51062 10108 51100 10164
rect 51156 10108 51166 10164
rect 51426 10108 51436 10164
rect 51492 10108 51660 10164
rect 51716 10108 51726 10164
rect 14914 9996 14924 10052
rect 14980 9996 17500 10052
rect 17556 9996 17566 10052
rect 17826 9996 17836 10052
rect 17892 9996 18620 10052
rect 18676 9996 19068 10052
rect 19124 9996 19134 10052
rect 25228 9996 26124 10052
rect 26180 9996 26684 10052
rect 26740 9996 26750 10052
rect 33170 9996 33180 10052
rect 33236 9996 33740 10052
rect 33796 9996 33806 10052
rect 33954 9996 33964 10052
rect 34020 9996 35084 10052
rect 35140 9996 35980 10052
rect 36036 9996 36046 10052
rect 43138 9996 43148 10052
rect 43204 9996 44716 10052
rect 44772 9996 45836 10052
rect 45892 9996 45902 10052
rect 47842 9996 47852 10052
rect 47908 9996 51828 10052
rect 51986 9996 51996 10052
rect 52052 9996 55580 10052
rect 55636 9996 55646 10052
rect 57362 9996 57372 10052
rect 57428 9996 58492 10052
rect 58548 9996 58558 10052
rect 33740 9940 33796 9996
rect 51772 9940 51828 9996
rect 16034 9884 16044 9940
rect 16100 9884 18284 9940
rect 18340 9884 18350 9940
rect 21074 9884 21084 9940
rect 21140 9884 21532 9940
rect 21588 9884 21756 9940
rect 21812 9884 28028 9940
rect 28084 9884 28094 9940
rect 33740 9884 34412 9940
rect 34468 9884 34478 9940
rect 34850 9884 34860 9940
rect 34916 9884 35532 9940
rect 35588 9884 35598 9940
rect 35746 9884 35756 9940
rect 35812 9884 41916 9940
rect 41972 9884 41982 9940
rect 45154 9884 45164 9940
rect 45220 9884 46508 9940
rect 46564 9884 46574 9940
rect 50306 9884 50316 9940
rect 50372 9884 51212 9940
rect 51268 9884 51278 9940
rect 51772 9884 52108 9940
rect 52164 9884 52174 9940
rect 52322 9884 52332 9940
rect 52388 9884 52556 9940
rect 52612 9884 53788 9940
rect 53844 9884 53854 9940
rect 55206 9884 55244 9940
rect 55300 9884 57708 9940
rect 57764 9884 57774 9940
rect 14690 9772 14700 9828
rect 14756 9772 15596 9828
rect 15652 9772 15662 9828
rect 22530 9772 22540 9828
rect 22596 9772 22988 9828
rect 23044 9772 24108 9828
rect 24164 9772 25228 9828
rect 25284 9772 25294 9828
rect 25526 9772 25564 9828
rect 25620 9772 25630 9828
rect 26002 9772 26012 9828
rect 26068 9772 26460 9828
rect 26516 9772 26796 9828
rect 26852 9772 26862 9828
rect 28130 9772 28140 9828
rect 28196 9772 29484 9828
rect 29540 9772 29550 9828
rect 34738 9772 34748 9828
rect 34804 9772 36540 9828
rect 36596 9772 36764 9828
rect 36820 9772 36830 9828
rect 38546 9772 38556 9828
rect 38612 9772 39116 9828
rect 39172 9772 40012 9828
rect 40068 9772 40078 9828
rect 41458 9772 41468 9828
rect 41524 9772 41692 9828
rect 41748 9772 42812 9828
rect 42868 9772 42878 9828
rect 48178 9772 48188 9828
rect 48244 9772 53340 9828
rect 53396 9772 53406 9828
rect 54786 9772 54796 9828
rect 54852 9772 58044 9828
rect 58100 9772 58110 9828
rect 2706 9660 2716 9716
rect 2772 9660 3276 9716
rect 3332 9660 16492 9716
rect 16548 9660 16558 9716
rect 29138 9660 29148 9716
rect 29204 9660 30604 9716
rect 30660 9660 30670 9716
rect 34066 9660 34076 9716
rect 34132 9660 35868 9716
rect 35924 9660 36092 9716
rect 36148 9660 36158 9716
rect 40338 9660 40348 9716
rect 40404 9660 42476 9716
rect 42532 9660 42542 9716
rect 47058 9660 47068 9716
rect 47124 9660 48524 9716
rect 48580 9660 48590 9716
rect 50082 9660 50092 9716
rect 50148 9660 50428 9716
rect 50484 9660 51324 9716
rect 51380 9660 51390 9716
rect 52098 9660 52108 9716
rect 52164 9660 54348 9716
rect 54404 9660 57372 9716
rect 57428 9660 57438 9716
rect 25106 9548 25116 9604
rect 25172 9548 25676 9604
rect 25732 9548 27468 9604
rect 27524 9548 33068 9604
rect 33124 9548 33134 9604
rect 38658 9548 38668 9604
rect 38724 9548 39340 9604
rect 39396 9548 42980 9604
rect 47394 9548 47404 9604
rect 47460 9548 48188 9604
rect 48244 9548 48254 9604
rect 50306 9548 50316 9604
rect 50372 9548 50540 9604
rect 50596 9548 50606 9604
rect 51874 9548 51884 9604
rect 51940 9548 53004 9604
rect 53060 9548 56028 9604
rect 56084 9548 56094 9604
rect 56438 9548 56476 9604
rect 56532 9548 56542 9604
rect 22866 9436 22876 9492
rect 22932 9436 23212 9492
rect 23268 9436 23772 9492
rect 23828 9436 24892 9492
rect 24948 9436 35420 9492
rect 35476 9436 35486 9492
rect 35858 9436 35868 9492
rect 35924 9436 39900 9492
rect 39956 9436 39966 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 42924 9380 42980 9548
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 26674 9324 26684 9380
rect 26740 9324 27132 9380
rect 27188 9324 42476 9380
rect 42532 9324 42542 9380
rect 42914 9324 42924 9380
rect 42980 9324 42990 9380
rect 56018 9324 56028 9380
rect 56084 9324 58268 9380
rect 58324 9324 58334 9380
rect 32498 9212 32508 9268
rect 32564 9212 32844 9268
rect 32900 9212 33852 9268
rect 33908 9212 33918 9268
rect 34626 9212 34636 9268
rect 34692 9212 35196 9268
rect 35252 9212 35262 9268
rect 40338 9212 40348 9268
rect 40404 9212 40908 9268
rect 40964 9212 42140 9268
rect 42196 9212 42206 9268
rect 43810 9212 43820 9268
rect 43876 9212 47292 9268
rect 47348 9212 47358 9268
rect 50372 9212 54460 9268
rect 54516 9212 54526 9268
rect 55122 9212 55132 9268
rect 55188 9212 56476 9268
rect 56532 9212 56542 9268
rect 50372 9156 50428 9212
rect 13010 9100 13020 9156
rect 13076 9100 13804 9156
rect 13860 9100 13870 9156
rect 26898 9100 26908 9156
rect 26964 9100 27356 9156
rect 27412 9100 28028 9156
rect 28084 9100 28094 9156
rect 34290 9100 34300 9156
rect 34356 9100 35532 9156
rect 35588 9100 35868 9156
rect 35924 9100 36372 9156
rect 36316 9044 36372 9100
rect 36988 9100 39340 9156
rect 39396 9100 39406 9156
rect 45714 9100 45724 9156
rect 45780 9100 50428 9156
rect 50754 9100 50764 9156
rect 50820 9100 51324 9156
rect 51380 9100 51390 9156
rect 52658 9100 52668 9156
rect 52724 9100 53452 9156
rect 53508 9100 53518 9156
rect 20290 8988 20300 9044
rect 20356 8988 21084 9044
rect 21140 8988 21150 9044
rect 30146 8988 30156 9044
rect 30212 8988 32172 9044
rect 32228 8988 32238 9044
rect 33618 8988 33628 9044
rect 33684 8988 34188 9044
rect 34244 8988 34254 9044
rect 36306 8988 36316 9044
rect 36372 8988 36382 9044
rect 34402 8876 34412 8932
rect 34468 8876 36764 8932
rect 36820 8876 36830 8932
rect 36988 8820 37044 9100
rect 38210 8988 38220 9044
rect 38276 8988 39452 9044
rect 39508 8988 39518 9044
rect 46722 8988 46732 9044
rect 46788 8988 51884 9044
rect 51940 8988 51950 9044
rect 37762 8876 37772 8932
rect 37828 8876 38668 8932
rect 38724 8876 38734 8932
rect 43138 8876 43148 8932
rect 43204 8876 43820 8932
rect 43876 8876 43886 8932
rect 47506 8876 47516 8932
rect 47572 8876 47964 8932
rect 48020 8876 48030 8932
rect 53554 8876 53564 8932
rect 53620 8876 55020 8932
rect 55076 8876 55086 8932
rect 31826 8764 31836 8820
rect 31892 8764 37044 8820
rect 42914 8764 42924 8820
rect 42980 8764 43260 8820
rect 43316 8764 43326 8820
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 24434 8428 24444 8484
rect 24500 8428 25116 8484
rect 25172 8428 25182 8484
rect 29810 8428 29820 8484
rect 29876 8428 30604 8484
rect 30660 8428 30670 8484
rect 33282 8428 33292 8484
rect 33348 8428 33628 8484
rect 33684 8428 33694 8484
rect 36082 8428 36092 8484
rect 36148 8428 37772 8484
rect 37828 8428 37838 8484
rect 42018 8428 42028 8484
rect 42084 8428 42364 8484
rect 42420 8428 42924 8484
rect 42980 8428 45388 8484
rect 45444 8428 45454 8484
rect 46834 8428 46844 8484
rect 46900 8428 47292 8484
rect 47348 8428 48636 8484
rect 48692 8428 48702 8484
rect 54338 8428 54348 8484
rect 54404 8428 55468 8484
rect 55524 8428 55534 8484
rect 19730 8316 19740 8372
rect 19796 8316 20412 8372
rect 20468 8316 21980 8372
rect 22036 8316 22764 8372
rect 22820 8316 22830 8372
rect 23538 8316 23548 8372
rect 23604 8316 24220 8372
rect 24276 8316 24892 8372
rect 24948 8316 25340 8372
rect 25396 8316 25406 8372
rect 30482 8316 30492 8372
rect 30548 8316 31164 8372
rect 31220 8316 32284 8372
rect 32340 8316 32350 8372
rect 34626 8316 34636 8372
rect 34692 8316 35532 8372
rect 35588 8316 35598 8372
rect 36418 8316 36428 8372
rect 36484 8316 36988 8372
rect 37044 8316 37212 8372
rect 37268 8316 37278 8372
rect 39218 8316 39228 8372
rect 39284 8316 39676 8372
rect 39732 8316 39742 8372
rect 40786 8316 40796 8372
rect 40852 8316 42588 8372
rect 42644 8316 42654 8372
rect 47058 8316 47068 8372
rect 47124 8316 47134 8372
rect 48402 8316 48412 8372
rect 48468 8316 49532 8372
rect 49588 8316 49598 8372
rect 51986 8316 51996 8372
rect 52052 8316 53788 8372
rect 53844 8316 53854 8372
rect 57474 8316 57484 8372
rect 57540 8316 58828 8372
rect 58884 8316 58894 8372
rect 47068 8260 47124 8316
rect 17266 8204 17276 8260
rect 17332 8204 18508 8260
rect 18564 8204 19180 8260
rect 19236 8204 19246 8260
rect 20626 8204 20636 8260
rect 20692 8204 22204 8260
rect 22260 8204 22270 8260
rect 24994 8204 25004 8260
rect 25060 8204 25900 8260
rect 25956 8204 26124 8260
rect 26180 8204 26190 8260
rect 26898 8204 26908 8260
rect 26964 8204 27468 8260
rect 27524 8204 27534 8260
rect 36530 8204 36540 8260
rect 36596 8204 37548 8260
rect 37604 8204 37614 8260
rect 38994 8204 39004 8260
rect 39060 8204 39452 8260
rect 39508 8204 41132 8260
rect 41188 8204 41198 8260
rect 41906 8204 41916 8260
rect 41972 8204 42700 8260
rect 42756 8204 43484 8260
rect 43540 8204 44044 8260
rect 44100 8204 44110 8260
rect 46834 8204 46844 8260
rect 46900 8204 47180 8260
rect 47236 8204 47740 8260
rect 47796 8204 47806 8260
rect 48066 8204 48076 8260
rect 48132 8204 52444 8260
rect 52500 8204 52510 8260
rect 52994 8204 53004 8260
rect 53060 8204 53340 8260
rect 53396 8204 53406 8260
rect 53554 8204 53564 8260
rect 53620 8204 54572 8260
rect 54628 8204 54638 8260
rect 55234 8204 55244 8260
rect 55300 8204 55916 8260
rect 55972 8204 55982 8260
rect 23874 8092 23884 8148
rect 23940 8092 26796 8148
rect 26852 8092 26862 8148
rect 27346 8092 27356 8148
rect 27412 8092 27804 8148
rect 27860 8092 28476 8148
rect 28532 8092 28542 8148
rect 33058 8092 33068 8148
rect 33124 8092 34188 8148
rect 34244 8092 35196 8148
rect 35252 8092 35262 8148
rect 38434 8092 38444 8148
rect 38500 8092 38780 8148
rect 38836 8092 39900 8148
rect 39956 8092 39966 8148
rect 46722 8092 46732 8148
rect 46788 8092 47852 8148
rect 47908 8092 49420 8148
rect 49476 8092 49486 8148
rect 49746 8092 49756 8148
rect 49812 8092 50988 8148
rect 51044 8092 51054 8148
rect 51650 8092 51660 8148
rect 51716 8092 53284 8148
rect 56018 8092 56028 8148
rect 56084 8092 57932 8148
rect 57988 8092 57998 8148
rect 49756 8036 49812 8092
rect 53228 8036 53284 8092
rect 25666 7980 25676 8036
rect 25732 7980 33180 8036
rect 33236 7980 33246 8036
rect 35074 7980 35084 8036
rect 35140 7980 37884 8036
rect 37940 7980 38332 8036
rect 38388 7980 38398 8036
rect 38612 7980 42028 8036
rect 42084 7980 42094 8036
rect 47142 7980 47180 8036
rect 47236 7980 47246 8036
rect 49074 7980 49084 8036
rect 49140 7980 49812 8036
rect 49970 7980 49980 8036
rect 50036 7980 51212 8036
rect 51268 7980 51278 8036
rect 51762 7980 51772 8036
rect 51828 7980 52780 8036
rect 52836 7980 52846 8036
rect 53218 7980 53228 8036
rect 53284 7980 55468 8036
rect 55524 7980 55534 8036
rect 55794 7980 55804 8036
rect 55860 7980 58716 8036
rect 58772 7980 58782 8036
rect 38612 7924 38668 7980
rect 22530 7868 22540 7924
rect 22596 7868 34636 7924
rect 34692 7868 34702 7924
rect 34860 7868 38668 7924
rect 41356 7868 44380 7924
rect 44436 7868 46396 7924
rect 46452 7868 46956 7924
rect 47012 7868 47022 7924
rect 53778 7868 53788 7924
rect 53844 7868 54460 7924
rect 54516 7868 55244 7924
rect 55300 7868 55310 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 34860 7812 34916 7868
rect 41356 7812 41412 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 28466 7756 28476 7812
rect 28532 7756 30940 7812
rect 30996 7756 31006 7812
rect 32162 7756 32172 7812
rect 32228 7756 34916 7812
rect 36978 7756 36988 7812
rect 37044 7756 41412 7812
rect 41570 7756 41580 7812
rect 41636 7756 42700 7812
rect 42756 7756 43820 7812
rect 43876 7756 45500 7812
rect 45556 7756 46620 7812
rect 46676 7756 46686 7812
rect 41458 7644 41468 7700
rect 41524 7644 42476 7700
rect 42532 7644 42542 7700
rect 43362 7644 43372 7700
rect 43428 7644 44380 7700
rect 44436 7644 44446 7700
rect 47506 7644 47516 7700
rect 47572 7644 48188 7700
rect 48244 7644 48254 7700
rect 50082 7644 50092 7700
rect 50148 7644 50652 7700
rect 50708 7644 50718 7700
rect 56802 7644 56812 7700
rect 56868 7644 58044 7700
rect 58100 7644 58110 7700
rect 28466 7532 28476 7588
rect 28532 7532 30044 7588
rect 30100 7532 30110 7588
rect 36530 7532 36540 7588
rect 36596 7532 37660 7588
rect 37716 7532 37726 7588
rect 45714 7532 45724 7588
rect 45780 7532 46844 7588
rect 46900 7532 46910 7588
rect 47058 7532 47068 7588
rect 47124 7532 47852 7588
rect 47908 7532 47918 7588
rect 20738 7420 20748 7476
rect 20804 7420 21644 7476
rect 21700 7420 21710 7476
rect 22082 7420 22092 7476
rect 22148 7420 23212 7476
rect 23268 7420 23436 7476
rect 23492 7420 23502 7476
rect 23650 7420 23660 7476
rect 23716 7420 24556 7476
rect 24612 7420 25676 7476
rect 25732 7420 25742 7476
rect 28130 7420 28140 7476
rect 28196 7420 28700 7476
rect 28756 7420 29036 7476
rect 29092 7420 29820 7476
rect 29876 7420 29886 7476
rect 34514 7420 34524 7476
rect 34580 7420 55804 7476
rect 55860 7420 55870 7476
rect 24658 7308 24668 7364
rect 24724 7308 25788 7364
rect 25844 7308 25854 7364
rect 27458 7308 27468 7364
rect 27524 7308 28364 7364
rect 28420 7308 28430 7364
rect 30930 7308 30940 7364
rect 30996 7308 31724 7364
rect 31780 7308 37884 7364
rect 37940 7308 37950 7364
rect 46162 7308 46172 7364
rect 46228 7308 46732 7364
rect 46788 7308 46798 7364
rect 48850 7308 48860 7364
rect 48916 7308 50204 7364
rect 50260 7308 53340 7364
rect 53396 7308 53406 7364
rect 23202 7196 23212 7252
rect 23268 7196 24556 7252
rect 24612 7196 24622 7252
rect 31266 7196 31276 7252
rect 31332 7196 35084 7252
rect 35140 7196 35150 7252
rect 47954 7196 47964 7252
rect 48020 7196 49644 7252
rect 49700 7196 49710 7252
rect 50306 7196 50316 7252
rect 50372 7196 51996 7252
rect 52052 7196 53004 7252
rect 53060 7196 54908 7252
rect 54964 7196 54974 7252
rect 22306 7084 22316 7140
rect 22372 7084 22876 7140
rect 22932 7084 29036 7140
rect 29092 7084 29102 7140
rect 45602 7084 45612 7140
rect 45668 7084 53788 7140
rect 53844 7084 54348 7140
rect 54404 7084 54414 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19394 6972 19404 7028
rect 19460 6972 20972 7028
rect 21028 6972 21038 7028
rect 39890 6972 39900 7028
rect 39956 6972 44604 7028
rect 44660 6972 47516 7028
rect 47572 6972 48076 7028
rect 48132 6972 48142 7028
rect 51090 6972 51100 7028
rect 51156 6972 51548 7028
rect 51604 6972 57148 7028
rect 57204 6972 57214 7028
rect 51314 6860 51324 6916
rect 51380 6860 53564 6916
rect 53620 6860 53630 6916
rect 59200 6804 59800 6832
rect 35298 6748 35308 6804
rect 35364 6748 36204 6804
rect 36260 6748 36270 6804
rect 36530 6748 36540 6804
rect 36596 6748 38332 6804
rect 38388 6748 38398 6804
rect 48514 6748 48524 6804
rect 48580 6748 49196 6804
rect 49252 6748 49532 6804
rect 49588 6748 49598 6804
rect 55346 6748 55356 6804
rect 55412 6748 59800 6804
rect 59200 6720 59800 6748
rect 19282 6636 19292 6692
rect 19348 6636 20412 6692
rect 20468 6636 20478 6692
rect 27458 6636 27468 6692
rect 27524 6636 28028 6692
rect 28084 6636 28094 6692
rect 30818 6636 30828 6692
rect 30884 6636 31612 6692
rect 31668 6636 31678 6692
rect 31826 6636 31836 6692
rect 31892 6636 32844 6692
rect 32900 6636 32910 6692
rect 33282 6636 33292 6692
rect 33348 6636 33740 6692
rect 33796 6636 33806 6692
rect 34626 6636 34636 6692
rect 34692 6636 36316 6692
rect 36372 6636 36382 6692
rect 37986 6636 37996 6692
rect 38052 6636 38556 6692
rect 38612 6636 38780 6692
rect 38836 6636 38846 6692
rect 43586 6636 43596 6692
rect 43652 6636 44492 6692
rect 44548 6636 44558 6692
rect 46610 6636 46620 6692
rect 46676 6636 47628 6692
rect 47684 6636 47694 6692
rect 48178 6636 48188 6692
rect 48244 6636 49308 6692
rect 49364 6636 49374 6692
rect 49858 6636 49868 6692
rect 49924 6636 50652 6692
rect 50708 6636 50718 6692
rect 52546 6636 52556 6692
rect 52612 6636 53452 6692
rect 53508 6636 53518 6692
rect 54226 6636 54236 6692
rect 54292 6636 54572 6692
rect 54628 6636 54638 6692
rect 56774 6636 56812 6692
rect 56868 6636 56878 6692
rect 27122 6524 27132 6580
rect 27188 6524 30716 6580
rect 30772 6524 31388 6580
rect 31444 6524 31454 6580
rect 37090 6524 37100 6580
rect 37156 6524 46060 6580
rect 46116 6524 46126 6580
rect 47394 6524 47404 6580
rect 47460 6524 48412 6580
rect 48468 6524 48478 6580
rect 48626 6524 48636 6580
rect 48692 6524 50988 6580
rect 51044 6524 52108 6580
rect 52164 6524 52174 6580
rect 54114 6524 54124 6580
rect 54180 6524 55356 6580
rect 55412 6524 55692 6580
rect 55748 6524 55758 6580
rect 32386 6412 32396 6468
rect 32452 6412 33068 6468
rect 33124 6412 33134 6468
rect 35074 6412 35084 6468
rect 35140 6412 35532 6468
rect 35588 6412 35980 6468
rect 36036 6412 36046 6468
rect 45378 6412 45388 6468
rect 45444 6412 48132 6468
rect 49970 6412 49980 6468
rect 50036 6412 50204 6468
rect 50260 6412 51996 6468
rect 52052 6412 52062 6468
rect 28130 6300 28140 6356
rect 28196 6300 29484 6356
rect 29540 6300 42588 6356
rect 42644 6300 44044 6356
rect 44100 6300 45276 6356
rect 45332 6300 45342 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 48076 6244 48132 6412
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 24546 6188 24556 6244
rect 24612 6188 28252 6244
rect 28308 6188 28318 6244
rect 29810 6188 29820 6244
rect 29876 6188 44380 6244
rect 44436 6188 45948 6244
rect 46004 6188 46014 6244
rect 48066 6188 48076 6244
rect 48132 6188 48142 6244
rect 19618 6076 19628 6132
rect 19684 6076 20636 6132
rect 20692 6076 21420 6132
rect 21476 6076 21486 6132
rect 31154 6076 31164 6132
rect 31220 6076 33740 6132
rect 33796 6076 33806 6132
rect 45378 6076 45388 6132
rect 45444 6076 48188 6132
rect 48244 6076 48254 6132
rect 48514 6076 48524 6132
rect 48580 6076 49756 6132
rect 49812 6076 49822 6132
rect 53778 6076 53788 6132
rect 53844 6076 54012 6132
rect 54068 6076 54078 6132
rect 32610 5964 32620 6020
rect 32676 5964 33628 6020
rect 33684 5964 33694 6020
rect 40898 5964 40908 6020
rect 40964 5964 42812 6020
rect 42868 5964 43820 6020
rect 43876 5964 44380 6020
rect 44436 5964 44446 6020
rect 52434 5964 52444 6020
rect 52500 5964 53004 6020
rect 53060 5964 54908 6020
rect 54964 5964 54974 6020
rect 32162 5852 32172 5908
rect 32228 5852 33964 5908
rect 34020 5852 35196 5908
rect 35252 5852 35262 5908
rect 35746 5852 35756 5908
rect 35812 5852 37324 5908
rect 37380 5852 49420 5908
rect 49476 5852 49486 5908
rect 50372 5852 54012 5908
rect 54068 5852 55468 5908
rect 55524 5852 57372 5908
rect 57428 5852 57438 5908
rect 31714 5740 31724 5796
rect 31780 5740 34188 5796
rect 34244 5740 35308 5796
rect 35364 5740 35374 5796
rect 35970 5740 35980 5796
rect 36036 5740 36652 5796
rect 36708 5740 37100 5796
rect 37156 5740 37166 5796
rect 43026 5740 43036 5796
rect 43092 5740 43484 5796
rect 43540 5740 47404 5796
rect 47460 5740 47470 5796
rect 50306 5740 50316 5796
rect 50372 5740 50428 5852
rect 23314 5516 23324 5572
rect 23380 5516 34636 5572
rect 34692 5516 34702 5572
rect 200 5460 800 5488
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 200 5404 1932 5460
rect 1988 5404 1998 5460
rect 46834 5404 46844 5460
rect 46900 5404 47628 5460
rect 47684 5404 48300 5460
rect 48356 5404 48366 5460
rect 200 5376 800 5404
rect 31490 5292 31500 5348
rect 31556 5292 32396 5348
rect 32452 5292 32462 5348
rect 33730 5292 33740 5348
rect 33796 5292 47964 5348
rect 48020 5292 48030 5348
rect 28354 5180 28364 5236
rect 28420 5180 31164 5236
rect 31220 5180 31230 5236
rect 34514 5180 34524 5236
rect 34580 5180 36540 5236
rect 36596 5180 37212 5236
rect 37268 5180 38220 5236
rect 38276 5180 38286 5236
rect 46722 5180 46732 5236
rect 46788 5180 47852 5236
rect 47908 5180 47918 5236
rect 54338 5180 54348 5236
rect 54404 5180 55580 5236
rect 55636 5180 55646 5236
rect 18834 5068 18844 5124
rect 18900 5068 20524 5124
rect 20580 5068 21868 5124
rect 21924 5068 21934 5124
rect 24098 5068 24108 5124
rect 24164 5068 24556 5124
rect 24612 5068 24622 5124
rect 37762 5068 37772 5124
rect 37828 5068 41916 5124
rect 41972 5068 42588 5124
rect 42644 5068 42654 5124
rect 49420 5068 50428 5124
rect 49420 5012 49476 5068
rect 50372 5012 50428 5068
rect 22418 4956 22428 5012
rect 22484 4956 23100 5012
rect 23156 4956 23772 5012
rect 23828 4956 23838 5012
rect 23986 4956 23996 5012
rect 24052 4956 25452 5012
rect 25508 4956 25518 5012
rect 33506 4956 33516 5012
rect 33572 4956 38444 5012
rect 38500 4956 38510 5012
rect 43586 4956 43596 5012
rect 43652 4956 49476 5012
rect 49634 4956 49644 5012
rect 49700 4956 50204 5012
rect 50260 4956 50270 5012
rect 50372 4956 56924 5012
rect 56980 4956 56990 5012
rect 22530 4844 22540 4900
rect 22596 4844 25116 4900
rect 25172 4844 25182 4900
rect 25330 4844 25340 4900
rect 25396 4844 54236 4900
rect 54292 4844 54302 4900
rect 21970 4732 21980 4788
rect 22036 4732 23884 4788
rect 23940 4732 23950 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 32386 4620 32396 4676
rect 32452 4620 33180 4676
rect 33236 4620 33516 4676
rect 33572 4620 50428 4676
rect 50372 4564 50428 4620
rect 2706 4508 2716 4564
rect 2772 4508 3276 4564
rect 3332 4508 9212 4564
rect 9268 4508 9278 4564
rect 29362 4508 29372 4564
rect 29428 4508 29820 4564
rect 29876 4508 32956 4564
rect 33012 4508 33022 4564
rect 37426 4508 37436 4564
rect 37492 4508 38780 4564
rect 38836 4508 40124 4564
rect 40180 4508 41132 4564
rect 41188 4508 41198 4564
rect 50372 4508 52780 4564
rect 52836 4508 52846 4564
rect 23650 4396 23660 4452
rect 23716 4396 26348 4452
rect 26404 4396 26414 4452
rect 30594 4396 30604 4452
rect 30660 4396 33852 4452
rect 33908 4396 33918 4452
rect 37538 4396 37548 4452
rect 37604 4396 39340 4452
rect 39396 4396 39406 4452
rect 48514 4396 48524 4452
rect 48580 4396 50652 4452
rect 50708 4396 50718 4452
rect 55906 4396 55916 4452
rect 55972 4396 57484 4452
rect 57540 4396 57550 4452
rect 20626 4284 20636 4340
rect 20692 4284 23100 4340
rect 23156 4284 23166 4340
rect 26674 4284 26684 4340
rect 26740 4284 31836 4340
rect 31892 4284 31902 4340
rect 34962 4284 34972 4340
rect 35028 4284 35644 4340
rect 35700 4284 36876 4340
rect 36932 4284 36942 4340
rect 37986 4284 37996 4340
rect 38052 4284 39452 4340
rect 39508 4284 40012 4340
rect 40068 4284 40078 4340
rect 54338 4284 54348 4340
rect 54404 4284 54908 4340
rect 54964 4284 54974 4340
rect 56690 4284 56700 4340
rect 56756 4284 57708 4340
rect 57764 4284 57774 4340
rect 25554 4172 25564 4228
rect 25620 4172 28588 4228
rect 28644 4172 28654 4228
rect 47954 4172 47964 4228
rect 48020 4172 48300 4228
rect 48356 4172 58604 4228
rect 58660 4172 58670 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 33618 3612 33628 3668
rect 33684 3612 34524 3668
rect 34580 3612 34590 3668
rect 36866 3612 36876 3668
rect 36932 3612 49644 3668
rect 49700 3612 49710 3668
rect 50418 3612 50428 3668
rect 50484 3612 51324 3668
rect 51380 3612 51390 3668
rect 26786 3500 26796 3556
rect 26852 3500 27356 3556
rect 27412 3500 28476 3556
rect 28532 3500 28542 3556
rect 30370 3500 30380 3556
rect 30436 3500 40012 3556
rect 40068 3500 40908 3556
rect 40964 3500 40974 3556
rect 44258 3500 44268 3556
rect 44324 3500 45164 3556
rect 45220 3500 45230 3556
rect 5058 3388 5068 3444
rect 5124 3388 5852 3444
rect 5908 3388 5918 3444
rect 16818 3388 16828 3444
rect 16884 3388 17612 3444
rect 17668 3388 17678 3444
rect 41794 3276 41804 3332
rect 41860 3276 44940 3332
rect 44996 3276 45006 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 27906 3052 27916 3108
rect 27972 3052 49644 3108
rect 49700 3052 49710 3108
rect 30930 2940 30940 2996
rect 30996 2940 49868 2996
rect 49924 2940 49934 2996
rect 32722 2828 32732 2884
rect 32788 2828 49084 2884
rect 49140 2828 49150 2884
rect 23874 2716 23884 2772
rect 23940 2716 56700 2772
rect 56756 2716 56766 2772
rect 3154 2604 3164 2660
rect 3220 2604 43372 2660
rect 43428 2604 43438 2660
rect 40226 2492 40236 2548
rect 40292 2492 53116 2548
rect 53172 2492 53182 2548
rect 18 1820 28 1876
rect 84 1820 1932 1876
rect 1988 1820 1998 1876
rect 28466 1596 28476 1652
rect 28532 1596 54124 1652
rect 54180 1596 54190 1652
rect 33282 1484 33292 1540
rect 33348 1484 48748 1540
rect 48804 1484 48814 1540
rect 59200 1428 59800 1456
rect 55234 1372 55244 1428
rect 55300 1372 59800 1428
rect 59200 1344 59800 1372
<< via3 >>
rect 6076 58492 6132 58548
rect 7868 58268 7924 58324
rect 21308 57484 21364 57540
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 31276 56364 31332 56420
rect 18508 56028 18564 56084
rect 5628 55916 5684 55972
rect 6524 55916 6580 55972
rect 10108 55916 10164 55972
rect 11676 55804 11732 55860
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 18396 55580 18452 55636
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 32396 55356 32452 55412
rect 2828 55244 2884 55300
rect 30156 55244 30212 55300
rect 15092 55132 15148 55188
rect 22316 55020 22372 55076
rect 26852 54908 26908 54964
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 18172 54796 18228 54852
rect 11452 54684 11508 54740
rect 14700 54684 14756 54740
rect 30156 54684 30212 54740
rect 18284 54572 18340 54628
rect 12684 54460 12740 54516
rect 26796 54460 26852 54516
rect 16716 54348 16772 54404
rect 9996 54236 10052 54292
rect 18172 54236 18228 54292
rect 19068 54236 19124 54292
rect 5964 54124 6020 54180
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 8204 54012 8260 54068
rect 18732 54012 18788 54068
rect 8316 53900 8372 53956
rect 8428 53788 8484 53844
rect 25004 53788 25060 53844
rect 6636 53676 6692 53732
rect 12684 53676 12740 53732
rect 14812 53676 14868 53732
rect 18284 53676 18340 53732
rect 13468 53564 13524 53620
rect 3948 53452 4004 53508
rect 12572 53452 12628 53508
rect 19628 53564 19684 53620
rect 7980 53340 8036 53396
rect 19628 53340 19684 53396
rect 11676 53228 11732 53284
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 6300 53116 6356 53172
rect 9996 53116 10052 53172
rect 9884 53004 9940 53060
rect 14812 53004 14868 53060
rect 8876 52892 8932 52948
rect 13132 52892 13188 52948
rect 15148 52892 15204 52948
rect 8540 52668 8596 52724
rect 14700 52668 14756 52724
rect 15932 52780 15988 52836
rect 16492 52780 16548 52836
rect 20300 52668 20356 52724
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19404 52332 19460 52388
rect 9436 52220 9492 52276
rect 12460 52220 12516 52276
rect 12684 52220 12740 52276
rect 6972 52108 7028 52164
rect 16380 52108 16436 52164
rect 24892 51996 24948 52052
rect 12348 51884 12404 51940
rect 15484 51884 15540 51940
rect 7532 51772 7588 51828
rect 15260 51772 15316 51828
rect 21756 51772 21812 51828
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 7868 51660 7924 51716
rect 9212 51660 9268 51716
rect 33740 51660 33796 51716
rect 6524 51548 6580 51604
rect 16716 51548 16772 51604
rect 21308 51548 21364 51604
rect 7980 51436 8036 51492
rect 12236 51436 12292 51492
rect 14252 51436 14308 51492
rect 9324 51324 9380 51380
rect 12124 51324 12180 51380
rect 16380 51324 16436 51380
rect 4844 51212 4900 51268
rect 5180 51212 5236 51268
rect 8876 51212 8932 51268
rect 33740 51212 33796 51268
rect 3724 50988 3780 51044
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 3612 50876 3668 50932
rect 5516 50876 5572 50932
rect 8764 50876 8820 50932
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 5516 50652 5572 50708
rect 16940 50652 16996 50708
rect 17836 50652 17892 50708
rect 18396 50652 18452 50708
rect 3052 50540 3108 50596
rect 4284 50540 4340 50596
rect 14028 50540 14084 50596
rect 14252 50540 14308 50596
rect 3836 50428 3892 50484
rect 5068 50428 5124 50484
rect 6748 50428 6804 50484
rect 9100 50428 9156 50484
rect 13356 50428 13412 50484
rect 13580 50428 13636 50484
rect 16940 50428 16996 50484
rect 18284 50428 18340 50484
rect 22540 50428 22596 50484
rect 27020 50428 27076 50484
rect 4956 50316 5012 50372
rect 8316 50316 8372 50372
rect 11452 50316 11508 50372
rect 14924 50316 14980 50372
rect 6860 50204 6916 50260
rect 4956 50092 5012 50148
rect 9324 50092 9380 50148
rect 14700 50092 14756 50148
rect 15036 50092 15092 50148
rect 23212 50204 23268 50260
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4172 49980 4228 50036
rect 16604 49980 16660 50036
rect 8204 49868 8260 49924
rect 9436 49868 9492 49924
rect 19516 49868 19572 49924
rect 20188 49868 20244 49924
rect 8316 49756 8372 49812
rect 16828 49756 16884 49812
rect 19628 49756 19684 49812
rect 22652 49756 22708 49812
rect 9996 49644 10052 49700
rect 10668 49644 10724 49700
rect 11676 49644 11732 49700
rect 14028 49644 14084 49700
rect 33964 49644 34020 49700
rect 18620 49532 18676 49588
rect 7084 49420 7140 49476
rect 23100 49420 23156 49476
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 21868 49308 21924 49364
rect 22092 49308 22148 49364
rect 3276 49196 3332 49252
rect 3836 49196 3892 49252
rect 4956 49196 5012 49252
rect 9436 49196 9492 49252
rect 10668 49196 10724 49252
rect 12236 49196 12292 49252
rect 36764 49420 36820 49476
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 31164 49196 31220 49252
rect 6076 49084 6132 49140
rect 7980 49084 8036 49140
rect 10108 49084 10164 49140
rect 15596 49084 15652 49140
rect 20188 49084 20244 49140
rect 24668 49084 24724 49140
rect 4060 48972 4116 49028
rect 15708 48972 15764 49028
rect 5068 48860 5124 48916
rect 8540 48860 8596 48916
rect 11676 48860 11732 48916
rect 22316 48860 22372 48916
rect 23212 48860 23268 48916
rect 27020 48860 27076 48916
rect 3724 48748 3780 48804
rect 22540 48748 22596 48804
rect 35756 48748 35812 48804
rect 3388 48636 3444 48692
rect 19516 48636 19572 48692
rect 20188 48636 20244 48692
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 15148 48524 15204 48580
rect 18284 48524 18340 48580
rect 8092 48412 8148 48468
rect 12348 48412 12404 48468
rect 23100 48412 23156 48468
rect 9884 48300 9940 48356
rect 16492 48300 16548 48356
rect 16828 48300 16884 48356
rect 6524 48188 6580 48244
rect 6860 48188 6916 48244
rect 11116 48188 11172 48244
rect 11452 48188 11508 48244
rect 12572 48188 12628 48244
rect 8540 48076 8596 48132
rect 11788 48076 11844 48132
rect 17836 48076 17892 48132
rect 18620 48076 18676 48132
rect 35644 48076 35700 48132
rect 3948 47964 4004 48020
rect 11452 47964 11508 48020
rect 18732 47964 18788 48020
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 36764 47852 36820 47908
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 15148 47740 15204 47796
rect 34300 47740 34356 47796
rect 3276 47628 3332 47684
rect 6860 47628 6916 47684
rect 4060 47516 4116 47572
rect 32396 47516 32452 47572
rect 33068 47516 33124 47572
rect 4172 47404 4228 47460
rect 18284 47404 18340 47460
rect 25004 47404 25060 47460
rect 32844 47404 32900 47460
rect 9212 47292 9268 47348
rect 9660 47292 9716 47348
rect 34300 47292 34356 47348
rect 38108 47292 38164 47348
rect 43372 47292 43428 47348
rect 16044 47180 16100 47236
rect 5852 47068 5908 47124
rect 8092 47068 8148 47124
rect 9212 47068 9268 47124
rect 24892 47068 24948 47124
rect 32844 47068 32900 47124
rect 33068 47068 33124 47124
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 21756 46956 21812 47012
rect 20188 46844 20244 46900
rect 4284 46732 4340 46788
rect 19628 46732 19684 46788
rect 3724 46620 3780 46676
rect 13244 46620 13300 46676
rect 18396 46620 18452 46676
rect 18956 46620 19012 46676
rect 11564 46508 11620 46564
rect 32060 46508 32116 46564
rect 32732 46508 32788 46564
rect 3500 46396 3556 46452
rect 6636 46396 6692 46452
rect 6972 46396 7028 46452
rect 8652 46396 8708 46452
rect 13692 46396 13748 46452
rect 14700 46396 14756 46452
rect 16156 46396 16212 46452
rect 19516 46396 19572 46452
rect 38108 46396 38164 46452
rect 3836 46284 3892 46340
rect 9436 46284 9492 46340
rect 13804 46284 13860 46340
rect 24668 46284 24724 46340
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 6748 46172 6804 46228
rect 15820 46172 15876 46228
rect 3724 46060 3780 46116
rect 4060 45948 4116 46004
rect 10108 45948 10164 46004
rect 12796 45948 12852 46004
rect 13580 45948 13636 46004
rect 33740 45948 33796 46004
rect 3388 45836 3444 45892
rect 8428 45836 8484 45892
rect 8988 45836 9044 45892
rect 16156 45836 16212 45892
rect 16940 45836 16996 45892
rect 18396 45836 18452 45892
rect 31612 45836 31668 45892
rect 3948 45724 4004 45780
rect 13804 45724 13860 45780
rect 15372 45724 15428 45780
rect 20524 45724 20580 45780
rect 4060 45612 4116 45668
rect 10108 45612 10164 45668
rect 3948 45500 4004 45556
rect 20188 45500 20244 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 8540 45388 8596 45444
rect 9772 45388 9828 45444
rect 10220 45388 10276 45444
rect 12124 45388 12180 45444
rect 15596 45388 15652 45444
rect 16716 45388 16772 45444
rect 3612 45164 3668 45220
rect 8540 45164 8596 45220
rect 9212 45164 9268 45220
rect 15372 45164 15428 45220
rect 18620 45164 18676 45220
rect 2156 45052 2212 45108
rect 7532 45052 7588 45108
rect 8652 45052 8708 45108
rect 12012 44940 12068 44996
rect 34524 45052 34580 45108
rect 19180 44828 19236 44884
rect 20188 44828 20244 44884
rect 20524 44828 20580 44884
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 13692 44716 13748 44772
rect 18844 44716 18900 44772
rect 31612 44716 31668 44772
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 35868 44604 35924 44660
rect 8204 44492 8260 44548
rect 9324 44492 9380 44548
rect 11900 44492 11956 44548
rect 14028 44492 14084 44548
rect 18956 44492 19012 44548
rect 6860 44380 6916 44436
rect 9324 44268 9380 44324
rect 9436 44156 9492 44212
rect 9772 44156 9828 44212
rect 13692 44156 13748 44212
rect 9212 44044 9268 44100
rect 9884 44044 9940 44100
rect 16604 44044 16660 44100
rect 23100 44044 23156 44100
rect 29596 44044 29652 44100
rect 12684 43932 12740 43988
rect 17164 43932 17220 43988
rect 18844 43932 18900 43988
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 6636 43820 6692 43876
rect 10332 43820 10388 43876
rect 12348 43820 12404 43876
rect 12572 43708 12628 43764
rect 13244 43708 13300 43764
rect 6748 43596 6804 43652
rect 9100 43596 9156 43652
rect 15260 43596 15316 43652
rect 18844 43596 18900 43652
rect 19404 43596 19460 43652
rect 10108 43484 10164 43540
rect 12348 43484 12404 43540
rect 17724 43484 17780 43540
rect 9660 43372 9716 43428
rect 9996 43372 10052 43428
rect 13692 43372 13748 43428
rect 18844 43260 18900 43316
rect 3500 43148 3556 43204
rect 11900 43148 11956 43204
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 3388 43036 3444 43092
rect 5292 43036 5348 43092
rect 6524 43036 6580 43092
rect 6076 42924 6132 42980
rect 6412 42924 6468 42980
rect 15260 42924 15316 42980
rect 6300 42812 6356 42868
rect 6188 42700 6244 42756
rect 26796 42700 26852 42756
rect 34860 42700 34916 42756
rect 11452 42588 11508 42644
rect 13468 42588 13524 42644
rect 15820 42588 15876 42644
rect 3388 42476 3444 42532
rect 8540 42476 8596 42532
rect 18956 42476 19012 42532
rect 22540 42476 22596 42532
rect 34860 42476 34916 42532
rect 15148 42364 15204 42420
rect 16044 42364 16100 42420
rect 3836 42252 3892 42308
rect 18620 42252 18676 42308
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 7420 42140 7476 42196
rect 9548 42140 9604 42196
rect 25228 42140 25284 42196
rect 3388 42028 3444 42084
rect 4844 42028 4900 42084
rect 5516 42028 5572 42084
rect 8540 42028 8596 42084
rect 11788 41916 11844 41972
rect 15036 41916 15092 41972
rect 2380 41804 2436 41860
rect 5292 41804 5348 41860
rect 13580 41804 13636 41860
rect 21196 41804 21252 41860
rect 6748 41692 6804 41748
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 22540 41580 22596 41636
rect 6412 41356 6468 41412
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 18956 41468 19012 41524
rect 19404 41468 19460 41524
rect 7980 41244 8036 41300
rect 6636 41132 6692 41188
rect 17164 41132 17220 41188
rect 19292 41132 19348 41188
rect 21196 41132 21252 41188
rect 17724 41020 17780 41076
rect 25228 41020 25284 41076
rect 2828 40908 2884 40964
rect 10332 40796 10388 40852
rect 15036 40796 15092 40852
rect 16604 40796 16660 40852
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 11676 40684 11732 40740
rect 26796 40572 26852 40628
rect 31164 40460 31220 40516
rect 15708 40348 15764 40404
rect 15036 40236 15092 40292
rect 18732 40236 18788 40292
rect 7308 40124 7364 40180
rect 13580 40012 13636 40068
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 8540 39788 8596 39844
rect 10668 39788 10724 39844
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 8988 39564 9044 39620
rect 22652 39452 22708 39508
rect 3612 39340 3668 39396
rect 7644 39228 7700 39284
rect 7980 39228 8036 39284
rect 9772 39228 9828 39284
rect 10220 39228 10276 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 8316 39116 8372 39172
rect 18620 39116 18676 39172
rect 3612 38892 3668 38948
rect 7196 38892 7252 38948
rect 16380 38892 16436 38948
rect 2380 38668 2436 38724
rect 31052 38668 31108 38724
rect 6076 38556 6132 38612
rect 3500 38444 3556 38500
rect 7868 38444 7924 38500
rect 13468 38444 13524 38500
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 7196 38220 7252 38276
rect 12348 38220 12404 38276
rect 16940 38220 16996 38276
rect 5404 38108 5460 38164
rect 7084 37996 7140 38052
rect 31052 37996 31108 38052
rect 5852 37884 5908 37940
rect 19292 37884 19348 37940
rect 7308 37772 7364 37828
rect 12348 37772 12404 37828
rect 6972 37660 7028 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 5964 37324 6020 37380
rect 6748 37212 6804 37268
rect 6972 37212 7028 37268
rect 7644 37212 7700 37268
rect 13356 37212 13412 37268
rect 10556 37100 10612 37156
rect 11900 37100 11956 37156
rect 6300 36988 6356 37044
rect 15820 36988 15876 37044
rect 35868 36988 35924 37044
rect 54908 36988 54964 37044
rect 7420 36876 7476 36932
rect 19068 36876 19124 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 6972 36764 7028 36820
rect 16156 36652 16212 36708
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 16492 36428 16548 36484
rect 19180 36316 19236 36372
rect 23100 36316 23156 36372
rect 7084 36204 7140 36260
rect 19068 36204 19124 36260
rect 29596 36204 29652 36260
rect 5292 36092 5348 36148
rect 15036 36092 15092 36148
rect 33740 36092 33796 36148
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 5740 35868 5796 35924
rect 6748 35868 6804 35924
rect 11564 35868 11620 35924
rect 21756 35868 21812 35924
rect 34076 35644 34132 35700
rect 3500 35420 3556 35476
rect 34076 35420 34132 35476
rect 4956 35308 5012 35364
rect 21756 35308 21812 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 2828 35196 2884 35252
rect 35756 35084 35812 35140
rect 5292 34972 5348 35028
rect 9884 34972 9940 35028
rect 16380 34860 16436 34916
rect 5852 34748 5908 34804
rect 54796 34636 54852 34692
rect 4956 34524 5012 34580
rect 50092 34524 50148 34580
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 5404 34300 5460 34356
rect 6300 34300 6356 34356
rect 10556 34300 10612 34356
rect 5740 34188 5796 34244
rect 3388 34076 3444 34132
rect 31164 33964 31220 34020
rect 2828 33852 2884 33908
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 8428 33628 8484 33684
rect 30828 33292 30884 33348
rect 3500 33180 3556 33236
rect 16044 33180 16100 33236
rect 31164 33180 31220 33236
rect 8764 33068 8820 33124
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 5628 32732 5684 32788
rect 11676 32732 11732 32788
rect 12796 32732 12852 32788
rect 16828 32732 16884 32788
rect 22092 32732 22148 32788
rect 3276 32620 3332 32676
rect 8764 32396 8820 32452
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 46396 32060 46452 32116
rect 49756 31948 49812 32004
rect 20300 31836 20356 31892
rect 12348 31612 12404 31668
rect 15932 31612 15988 31668
rect 53564 31836 53620 31892
rect 46396 31500 46452 31556
rect 19516 31388 19572 31444
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 8652 31276 8708 31332
rect 2828 31164 2884 31220
rect 14812 31164 14868 31220
rect 22540 31164 22596 31220
rect 49532 31052 49588 31108
rect 50316 30940 50372 30996
rect 10668 30716 10724 30772
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 32060 30492 32116 30548
rect 51436 30492 51492 30548
rect 15708 30268 15764 30324
rect 18396 30156 18452 30212
rect 5852 30044 5908 30100
rect 46284 29932 46340 29988
rect 55244 29820 55300 29876
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 9548 29596 9604 29652
rect 12460 29372 12516 29428
rect 2156 29260 2212 29316
rect 47068 29148 47124 29204
rect 51436 29148 51492 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 46956 28924 47012 28980
rect 12460 28812 12516 28868
rect 31276 28812 31332 28868
rect 3948 28588 4004 28644
rect 18508 28588 18564 28644
rect 2940 28476 2996 28532
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 42924 27692 42980 27748
rect 53452 27692 53508 27748
rect 47068 27580 47124 27636
rect 48636 27580 48692 27636
rect 50316 27580 50372 27636
rect 8204 27468 8260 27524
rect 42924 27468 42980 27524
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 48412 27356 48468 27412
rect 48636 27356 48692 27412
rect 49644 27356 49700 27412
rect 3052 27244 3108 27300
rect 41356 26908 41412 26964
rect 44492 26908 44548 26964
rect 49308 26908 49364 26964
rect 50316 26908 50372 26964
rect 36316 26796 36372 26852
rect 44492 26684 44548 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 53676 26460 53732 26516
rect 47404 26348 47460 26404
rect 41468 26124 41524 26180
rect 48748 26124 48804 26180
rect 44156 26012 44212 26068
rect 6188 25900 6244 25956
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 13356 25788 13412 25844
rect 48636 25788 48692 25844
rect 11116 25676 11172 25732
rect 11452 25564 11508 25620
rect 38668 25564 38724 25620
rect 45612 25452 45668 25508
rect 48636 25340 48692 25396
rect 38556 25228 38612 25284
rect 5516 25004 5572 25060
rect 18956 25004 19012 25060
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 30828 25004 30884 25060
rect 55692 25116 55748 25172
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 32732 24556 32788 24612
rect 41468 24556 41524 24612
rect 45388 24556 45444 24612
rect 48748 24556 48804 24612
rect 36540 24444 36596 24500
rect 51772 24444 51828 24500
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 34188 24332 34244 24388
rect 46508 24332 46564 24388
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 41468 23996 41524 24052
rect 50316 23996 50372 24052
rect 34748 23884 34804 23940
rect 36540 23884 36596 23940
rect 53452 23884 53508 23940
rect 47964 23772 48020 23828
rect 53676 23772 53732 23828
rect 42028 23660 42084 23716
rect 53900 23660 53956 23716
rect 34188 23548 34244 23604
rect 47964 23548 48020 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 8316 23324 8372 23380
rect 33964 23324 34020 23380
rect 46956 23324 47012 23380
rect 49196 23324 49252 23380
rect 50204 23212 50260 23268
rect 36316 23100 36372 23156
rect 46172 23100 46228 23156
rect 48972 23100 49028 23156
rect 53676 23100 53732 23156
rect 45500 22988 45556 23044
rect 49084 22988 49140 23044
rect 55020 22988 55076 23044
rect 12012 22876 12068 22932
rect 38780 22876 38836 22932
rect 46956 22876 47012 22932
rect 48748 22876 48804 22932
rect 49532 22876 49588 22932
rect 55356 22876 55412 22932
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 48860 22316 48916 22372
rect 35756 22092 35812 22148
rect 50204 22092 50260 22148
rect 51548 22092 51604 22148
rect 53340 22092 53396 22148
rect 53676 22092 53732 22148
rect 55356 22092 55412 22148
rect 50316 21980 50372 22036
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 51324 21868 51380 21924
rect 13132 21756 13188 21812
rect 48300 21756 48356 21812
rect 49644 21756 49700 21812
rect 51212 21756 51268 21812
rect 34524 21644 34580 21700
rect 43932 21644 43988 21700
rect 50316 21644 50372 21700
rect 52108 21644 52164 21700
rect 9436 21532 9492 21588
rect 21196 21532 21252 21588
rect 45612 21532 45668 21588
rect 46956 21532 47012 21588
rect 49196 21532 49252 21588
rect 51100 21532 51156 21588
rect 41020 21420 41076 21476
rect 48860 21420 48916 21476
rect 50316 21420 50372 21476
rect 51212 21420 51268 21476
rect 51548 21420 51604 21476
rect 53228 21420 53284 21476
rect 51100 21308 51156 21364
rect 52668 21308 52724 21364
rect 48748 21196 48804 21252
rect 53228 21196 53284 21252
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 41356 21084 41412 21140
rect 49980 21084 50036 21140
rect 41020 20972 41076 21028
rect 50988 20972 51044 21028
rect 43596 20860 43652 20916
rect 50316 20860 50372 20916
rect 46284 20748 46340 20804
rect 35644 20636 35700 20692
rect 47068 20636 47124 20692
rect 48636 20636 48692 20692
rect 50316 20636 50372 20692
rect 42140 20524 42196 20580
rect 48748 20524 48804 20580
rect 55580 20524 55636 20580
rect 48860 20412 48916 20468
rect 52220 20412 52276 20468
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 39452 20300 39508 20356
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 53452 20300 53508 20356
rect 35756 20188 35812 20244
rect 42252 20188 42308 20244
rect 55916 20188 55972 20244
rect 51100 20076 51156 20132
rect 52108 20076 52164 20132
rect 53676 20076 53732 20132
rect 38108 19964 38164 20020
rect 42252 19964 42308 20020
rect 43708 19964 43764 20020
rect 48524 19964 48580 20020
rect 51212 19964 51268 20020
rect 55244 19964 55300 20020
rect 44268 19852 44324 19908
rect 49084 19852 49140 19908
rect 51884 19852 51940 19908
rect 39452 19740 39508 19796
rect 40684 19740 40740 19796
rect 41468 19740 41524 19796
rect 45612 19740 45668 19796
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 46508 19628 46564 19684
rect 56028 19628 56084 19684
rect 34300 19516 34356 19572
rect 38108 19516 38164 19572
rect 39228 19516 39284 19572
rect 45276 19516 45332 19572
rect 47068 19516 47124 19572
rect 49196 19516 49252 19572
rect 55356 19516 55412 19572
rect 49980 19404 50036 19460
rect 50988 19404 51044 19460
rect 51212 19404 51268 19460
rect 51660 19404 51716 19460
rect 55468 19404 55524 19460
rect 51996 19292 52052 19348
rect 55356 19292 55412 19348
rect 43708 19180 43764 19236
rect 51212 19180 51268 19236
rect 51772 19180 51828 19236
rect 45948 19068 46004 19124
rect 48188 19068 48244 19124
rect 51100 19068 51156 19124
rect 51548 19068 51604 19124
rect 48972 18956 49028 19012
rect 51996 18956 52052 19012
rect 45724 18844 45780 18900
rect 55356 18844 55412 18900
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 49196 18732 49252 18788
rect 42252 18620 42308 18676
rect 43932 18620 43988 18676
rect 48412 18620 48468 18676
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 53900 18732 53956 18788
rect 45276 18508 45332 18564
rect 48636 18508 48692 18564
rect 48972 18508 49028 18564
rect 54460 18508 54516 18564
rect 49644 18396 49700 18452
rect 50988 18396 51044 18452
rect 53676 18396 53732 18452
rect 53900 18396 53956 18452
rect 55468 18396 55524 18452
rect 56476 18396 56532 18452
rect 33964 18284 34020 18340
rect 48860 18284 48916 18340
rect 39452 18172 39508 18228
rect 42252 18172 42308 18228
rect 46172 18172 46228 18228
rect 48524 18172 48580 18228
rect 49756 18172 49812 18228
rect 55580 18172 55636 18228
rect 42812 18060 42868 18116
rect 51324 18060 51380 18116
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 52332 17948 52388 18004
rect 53228 17948 53284 18004
rect 38780 17836 38836 17892
rect 51772 17724 51828 17780
rect 54796 17612 54852 17668
rect 55132 17612 55188 17668
rect 49756 17500 49812 17556
rect 50988 17500 51044 17556
rect 43148 17276 43204 17332
rect 44268 17276 44324 17332
rect 46060 17276 46116 17332
rect 51884 17276 51940 17332
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 34524 17164 34580 17220
rect 47516 17164 47572 17220
rect 51996 17164 52052 17220
rect 43596 17052 43652 17108
rect 45612 17052 45668 17108
rect 54012 17052 54068 17108
rect 36204 16940 36260 16996
rect 34524 16828 34580 16884
rect 36540 16828 36596 16884
rect 38780 16716 38836 16772
rect 51772 16716 51828 16772
rect 36540 16604 36596 16660
rect 42812 16604 42868 16660
rect 49532 16604 49588 16660
rect 34300 16492 34356 16548
rect 45500 16492 45556 16548
rect 56812 16492 56868 16548
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 49756 16380 49812 16436
rect 36204 16268 36260 16324
rect 42924 16268 42980 16324
rect 47180 16268 47236 16324
rect 48300 16268 48356 16324
rect 51436 16268 51492 16324
rect 54460 16268 54516 16324
rect 46060 16156 46116 16212
rect 50204 16156 50260 16212
rect 39116 16044 39172 16100
rect 43484 16044 43540 16100
rect 46172 16044 46228 16100
rect 49980 16044 50036 16100
rect 51100 16044 51156 16100
rect 51772 16044 51828 16100
rect 56700 16044 56756 16100
rect 47068 15932 47124 15988
rect 48412 15932 48468 15988
rect 49756 15932 49812 15988
rect 54012 15932 54068 15988
rect 41468 15820 41524 15876
rect 55804 15820 55860 15876
rect 56028 15820 56084 15876
rect 50204 15708 50260 15764
rect 51660 15708 51716 15764
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 40236 15596 40292 15652
rect 43708 15596 43764 15652
rect 48860 15596 48916 15652
rect 49644 15596 49700 15652
rect 51548 15596 51604 15652
rect 27916 15484 27972 15540
rect 54572 15484 54628 15540
rect 42812 15372 42868 15428
rect 48636 15372 48692 15428
rect 54460 15372 54516 15428
rect 56700 15372 56756 15428
rect 27916 15260 27972 15316
rect 43708 15260 43764 15316
rect 51548 15260 51604 15316
rect 47404 15148 47460 15204
rect 53452 15148 53508 15204
rect 55692 15148 55748 15204
rect 50204 15036 50260 15092
rect 43484 14924 43540 14980
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 50988 14812 51044 14868
rect 45948 14700 46004 14756
rect 51324 14700 51380 14756
rect 52332 14700 52388 14756
rect 39900 14588 39956 14644
rect 41580 14588 41636 14644
rect 50204 14588 50260 14644
rect 39228 14476 39284 14532
rect 43148 14476 43204 14532
rect 50092 14476 50148 14532
rect 33964 14252 34020 14308
rect 51996 14364 52052 14420
rect 57148 14364 57204 14420
rect 51548 14140 51604 14196
rect 52444 14140 52500 14196
rect 53340 14140 53396 14196
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 42140 14028 42196 14084
rect 51884 14028 51940 14084
rect 34748 13916 34804 13972
rect 39900 13692 39956 13748
rect 47068 13692 47124 13748
rect 51884 13692 51940 13748
rect 39228 13580 39284 13636
rect 49308 13580 49364 13636
rect 50988 13580 51044 13636
rect 55580 13580 55636 13636
rect 40684 13468 40740 13524
rect 45724 13468 45780 13524
rect 47964 13468 48020 13524
rect 55916 13468 55972 13524
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 41580 13356 41636 13412
rect 52220 13356 52276 13412
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 39452 13020 39508 13076
rect 46060 13020 46116 13076
rect 51100 13020 51156 13076
rect 52668 13020 52724 13076
rect 54908 13020 54964 13076
rect 55804 13020 55860 13076
rect 55020 12908 55076 12964
rect 44156 12796 44212 12852
rect 53452 12796 53508 12852
rect 39116 12572 39172 12628
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50988 12572 51044 12628
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 42700 12460 42756 12516
rect 57148 12460 57204 12516
rect 51212 12348 51268 12404
rect 49420 12124 49476 12180
rect 51212 12124 51268 12180
rect 51772 12124 51828 12180
rect 47516 12012 47572 12068
rect 48188 12012 48244 12068
rect 51324 12012 51380 12068
rect 53900 12124 53956 12180
rect 53452 12012 53508 12068
rect 46396 11900 46452 11956
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 44156 11788 44212 11844
rect 49420 11788 49476 11844
rect 53676 11788 53732 11844
rect 54460 11788 54516 11844
rect 38668 11676 38724 11732
rect 50316 11564 50372 11620
rect 49196 11452 49252 11508
rect 48748 11340 48804 11396
rect 43596 11228 43652 11284
rect 49980 11228 50036 11284
rect 42700 11116 42756 11172
rect 49644 11116 49700 11172
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 38668 10892 38724 10948
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 49532 10780 49588 10836
rect 49980 10556 50036 10612
rect 50988 10332 51044 10388
rect 25564 10220 25620 10276
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 48636 10108 48692 10164
rect 51100 10108 51156 10164
rect 51436 10108 51492 10164
rect 51996 9996 52052 10052
rect 55244 9884 55300 9940
rect 25564 9772 25620 9828
rect 48188 9772 48244 9828
rect 47068 9660 47124 9716
rect 56476 9548 56532 9604
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 55132 9212 55188 9268
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 45388 8428 45444 8484
rect 47180 8204 47236 8260
rect 53564 8204 53620 8260
rect 49756 8092 49812 8148
rect 42028 7980 42084 8036
rect 47180 7980 47236 8036
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 51548 6972 51604 7028
rect 54572 6636 54628 6692
rect 56812 6636 56868 6692
rect 55692 6524 55748 6580
rect 50204 6412 50260 6468
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 52444 5964 52500 6020
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
rect 49644 3052 49700 3108
rect 43372 2604 43428 2660
rect 40236 2492 40292 2548
rect 48748 1484 48804 1540
<< metal4 >>
rect 6076 58548 6132 58558
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 2828 55300 2884 55310
rect 2828 50428 2884 55244
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 3948 53508 4004 53518
rect 3724 51044 3780 51054
rect 3612 50932 3668 50942
rect 3052 50596 3108 50606
rect 2828 50372 2996 50428
rect 2156 45108 2212 45118
rect 2156 29316 2212 45052
rect 2380 41860 2436 41870
rect 2380 38724 2436 41804
rect 2380 38658 2436 38668
rect 2828 40964 2884 40974
rect 2828 35252 2884 40908
rect 2828 35186 2884 35196
rect 2828 33908 2884 33918
rect 2828 31220 2884 33852
rect 2828 31154 2884 31164
rect 2156 29250 2212 29260
rect 2940 28532 2996 50372
rect 2940 28466 2996 28476
rect 3052 27300 3108 50540
rect 3276 49252 3332 49262
rect 3276 47684 3332 49196
rect 3276 32676 3332 47628
rect 3388 48692 3444 48702
rect 3388 45892 3444 48636
rect 3388 45826 3444 45836
rect 3500 46452 3556 46462
rect 3500 43204 3556 46396
rect 3612 45220 3668 50876
rect 3724 48804 3780 50988
rect 3836 50484 3892 50494
rect 3836 49252 3892 50428
rect 3836 49186 3892 49196
rect 3724 48738 3780 48748
rect 3948 48020 4004 53452
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 5628 55972 5684 55982
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4284 50596 4340 50606
rect 4172 50036 4228 50046
rect 3724 46676 3780 46686
rect 3724 46116 3780 46620
rect 3724 46050 3780 46060
rect 3836 46340 3892 46350
rect 3612 45154 3668 45164
rect 3500 43138 3556 43148
rect 3388 43092 3444 43102
rect 3388 42532 3444 43036
rect 3388 42084 3444 42476
rect 3836 42308 3892 46284
rect 3948 45780 4004 47964
rect 4060 49028 4116 49038
rect 4060 47572 4116 48972
rect 4060 47506 4116 47516
rect 4172 47460 4228 49980
rect 4172 47394 4228 47404
rect 4284 46788 4340 50540
rect 4284 46722 4340 46732
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 3948 45714 4004 45724
rect 4060 46004 4116 46014
rect 4060 45668 4116 45948
rect 4060 45602 4116 45612
rect 3836 42242 3892 42252
rect 3948 45556 4004 45566
rect 3388 34132 3444 42028
rect 3612 39396 3668 39406
rect 3612 38948 3668 39340
rect 3612 38882 3668 38892
rect 3388 34066 3444 34076
rect 3500 38500 3556 38510
rect 3500 35476 3556 38444
rect 3500 33236 3556 35420
rect 3500 33170 3556 33180
rect 3276 32610 3332 32620
rect 3948 28644 4004 45500
rect 3948 28578 4004 28588
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4844 51268 4900 51278
rect 5180 51268 5236 51278
rect 4844 42084 4900 51212
rect 4956 51212 5180 51268
rect 4956 50372 5012 51212
rect 5180 51202 5236 51212
rect 5516 50932 5572 50942
rect 5516 50708 5572 50876
rect 5516 50642 5572 50652
rect 4956 50306 5012 50316
rect 5068 50484 5124 50494
rect 4956 50148 5012 50158
rect 4956 49252 5012 50092
rect 4956 49186 5012 49196
rect 5068 48916 5124 50428
rect 5068 48850 5124 48860
rect 4844 42018 4900 42028
rect 5292 43092 5348 43102
rect 5292 41860 5348 43036
rect 5292 41794 5348 41804
rect 5516 42084 5572 42094
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 5404 38164 5460 38174
rect 5292 36148 5348 36158
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4956 35364 5012 35374
rect 4956 34580 5012 35308
rect 5292 35028 5348 36092
rect 5292 34962 5348 34972
rect 4956 34514 5012 34524
rect 5404 34356 5460 38108
rect 5404 34290 5460 34300
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 3052 27234 3108 27244
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 5516 25060 5572 42028
rect 5628 32788 5684 55916
rect 5964 54180 6020 54190
rect 5852 47124 5908 47134
rect 5852 37940 5908 47068
rect 5740 35924 5796 35934
rect 5740 34244 5796 35868
rect 5740 34178 5796 34188
rect 5852 34804 5908 37884
rect 5964 37380 6020 54124
rect 6076 49140 6132 58492
rect 7868 58324 7924 58334
rect 6524 55972 6580 55982
rect 6076 49074 6132 49084
rect 6300 53172 6356 53182
rect 6076 42980 6132 42990
rect 6076 38612 6132 42924
rect 6300 42868 6356 53116
rect 6524 51604 6580 55916
rect 6524 51538 6580 51548
rect 6636 53732 6692 53742
rect 6524 48244 6580 48254
rect 6524 43092 6580 48188
rect 6636 46452 6692 53676
rect 6972 52164 7028 52174
rect 6636 46386 6692 46396
rect 6748 50484 6804 50494
rect 6748 46228 6804 50428
rect 6860 50260 6916 50270
rect 6860 48244 6916 50204
rect 6860 48178 6916 48188
rect 6748 46162 6804 46172
rect 6860 47684 6916 47694
rect 6860 44436 6916 47628
rect 6972 46452 7028 52108
rect 7532 51828 7588 51838
rect 6972 46386 7028 46396
rect 7084 49476 7140 49486
rect 6860 44370 6916 44380
rect 6524 43026 6580 43036
rect 6636 43876 6692 43886
rect 6076 38546 6132 38556
rect 6188 42756 6244 42766
rect 5964 37314 6020 37324
rect 5628 32722 5684 32732
rect 5852 30100 5908 34748
rect 5852 30034 5908 30044
rect 6188 25956 6244 42700
rect 6300 37044 6356 42812
rect 6412 42980 6468 42990
rect 6412 41412 6468 42924
rect 6412 41346 6468 41356
rect 6636 41188 6692 43820
rect 6748 43652 6804 43662
rect 7084 43652 7140 49420
rect 7532 45108 7588 51772
rect 7532 45042 7588 45052
rect 7868 51716 7924 58268
rect 21308 57540 21364 57550
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 18508 56084 18564 56094
rect 10108 55972 10164 55982
rect 9996 54292 10052 54302
rect 8204 54068 8260 54078
rect 6804 43596 7140 43652
rect 6748 41748 6804 43596
rect 6748 41682 6804 41692
rect 7420 42196 7476 42206
rect 6636 41122 6692 41132
rect 7308 40180 7364 40190
rect 7196 38948 7252 38958
rect 7196 38276 7252 38892
rect 7196 38210 7252 38220
rect 7084 38052 7140 38062
rect 6972 37716 7028 37726
rect 6300 34356 6356 36988
rect 6748 37268 6804 37278
rect 6748 35924 6804 37212
rect 6972 37268 7028 37660
rect 6972 36820 7028 37212
rect 6972 36754 7028 36764
rect 7084 36260 7140 37996
rect 7308 37828 7364 40124
rect 7308 37762 7364 37772
rect 7420 36932 7476 42140
rect 7644 39284 7700 39294
rect 7644 37268 7700 39228
rect 7868 38500 7924 51660
rect 7980 53396 8036 53406
rect 7980 51492 8036 53340
rect 7980 50428 8036 51436
rect 7980 50372 8148 50428
rect 7980 49140 8036 49150
rect 7980 41300 8036 49084
rect 8092 48468 8148 50372
rect 8204 49924 8260 54012
rect 8316 53956 8372 53966
rect 8316 50372 8372 53900
rect 8316 50306 8372 50316
rect 8428 53844 8484 53854
rect 8204 49858 8260 49868
rect 8092 47124 8148 48412
rect 8092 47058 8148 47068
rect 8316 49812 8372 49822
rect 7980 39284 8036 41244
rect 7980 39218 8036 39228
rect 8204 44548 8260 44558
rect 7868 38434 7924 38444
rect 7644 37202 7700 37212
rect 7420 36866 7476 36876
rect 7084 36194 7140 36204
rect 6748 35858 6804 35868
rect 6300 34290 6356 34300
rect 8204 27524 8260 44492
rect 8204 27458 8260 27468
rect 8316 39172 8372 49756
rect 6188 25890 6244 25900
rect 5516 24994 5572 25004
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 8316 23380 8372 39116
rect 8428 45892 8484 53788
rect 9996 53172 10052 54236
rect 9996 53106 10052 53116
rect 9884 53060 9940 53070
rect 8876 52948 8932 52958
rect 8540 52724 8596 52734
rect 8540 48916 8596 52668
rect 8876 51268 8932 52892
rect 9436 52276 9492 52286
rect 8876 51202 8932 51212
rect 9212 51716 9268 51726
rect 8540 48132 8596 48860
rect 8540 48066 8596 48076
rect 8764 50932 8820 50942
rect 8428 33684 8484 45836
rect 8652 46452 8708 46462
rect 8540 45444 8596 45454
rect 8540 45220 8596 45388
rect 8540 45154 8596 45164
rect 8652 45108 8708 46396
rect 8540 42532 8596 42542
rect 8540 42084 8596 42476
rect 8540 39844 8596 42028
rect 8540 39778 8596 39788
rect 8428 33618 8484 33628
rect 8652 31332 8708 45052
rect 8764 33124 8820 50876
rect 9100 50484 9156 50494
rect 8988 45892 9044 45902
rect 8988 39620 9044 45836
rect 9100 43652 9156 50428
rect 9212 47348 9268 51660
rect 9212 47282 9268 47292
rect 9324 51380 9380 51390
rect 9324 50148 9380 51324
rect 9212 47124 9268 47134
rect 9212 45220 9268 47068
rect 9212 44100 9268 45164
rect 9324 44548 9380 50092
rect 9436 49924 9492 52220
rect 9436 49858 9492 49868
rect 9436 49252 9492 49262
rect 9436 46340 9492 49196
rect 9884 48356 9940 53004
rect 9884 48290 9940 48300
rect 9996 49700 10052 49710
rect 9436 46274 9492 46284
rect 9660 47348 9716 47358
rect 9324 44324 9380 44492
rect 9324 44258 9380 44268
rect 9212 44034 9268 44044
rect 9436 44212 9492 44222
rect 9100 43586 9156 43596
rect 8988 39554 9044 39564
rect 8764 32452 8820 33068
rect 8764 32386 8820 32396
rect 8652 31266 8708 31276
rect 8316 23314 8372 23324
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 9436 21588 9492 44156
rect 9660 43428 9716 47292
rect 9660 43362 9716 43372
rect 9772 45444 9828 45454
rect 9772 44212 9828 45388
rect 9548 42196 9604 42206
rect 9548 29652 9604 42140
rect 9772 39284 9828 44156
rect 9772 39218 9828 39228
rect 9884 44100 9940 44110
rect 9884 35028 9940 44044
rect 9996 43428 10052 49644
rect 10108 49140 10164 55916
rect 11676 55860 11732 55870
rect 11452 54740 11508 54750
rect 11452 50372 11508 54684
rect 10108 46004 10164 49084
rect 10108 45938 10164 45948
rect 10668 49700 10724 49710
rect 10668 49252 10724 49644
rect 10108 45668 10164 45678
rect 10108 43540 10164 45612
rect 10108 43474 10164 43484
rect 10220 45444 10276 45454
rect 9996 43362 10052 43372
rect 10220 39284 10276 45388
rect 10332 43876 10388 43886
rect 10332 40852 10388 43820
rect 10332 40786 10388 40796
rect 10220 39218 10276 39228
rect 10668 39844 10724 49196
rect 9884 34962 9940 34972
rect 10556 37156 10612 37166
rect 10556 34356 10612 37100
rect 10556 34290 10612 34300
rect 10668 30772 10724 39788
rect 10668 30706 10724 30716
rect 11116 48244 11172 48254
rect 9548 29586 9604 29596
rect 11116 25732 11172 48188
rect 11452 48244 11508 50316
rect 11452 48178 11508 48188
rect 11676 53284 11732 55804
rect 18396 55636 18452 55646
rect 15092 55188 15148 55198
rect 14924 55132 15092 55188
rect 14700 54740 14756 54750
rect 14924 54740 14980 55132
rect 15092 55122 15148 55132
rect 14756 54684 14980 54740
rect 18172 54852 18228 54862
rect 12684 54516 12740 54526
rect 12684 53732 12740 54460
rect 11676 49700 11732 53228
rect 12572 53508 12628 53518
rect 12460 52276 12516 52286
rect 12348 51940 12404 51950
rect 12236 51492 12292 51502
rect 11676 48916 11732 49644
rect 11116 25666 11172 25676
rect 11452 48020 11508 48030
rect 11452 42644 11508 47964
rect 11452 25620 11508 42588
rect 11564 46564 11620 46574
rect 11564 35924 11620 46508
rect 11564 35858 11620 35868
rect 11676 40740 11732 48860
rect 12124 51380 12180 51390
rect 11788 48132 11844 48142
rect 11788 41972 11844 48076
rect 12124 45444 12180 51324
rect 12236 49252 12292 51436
rect 12236 49186 12292 49196
rect 12348 48468 12404 51884
rect 12348 48402 12404 48412
rect 12124 45378 12180 45388
rect 12012 44996 12068 45006
rect 11788 41906 11844 41916
rect 11900 44548 11956 44558
rect 11900 43204 11956 44492
rect 11676 32788 11732 40684
rect 11900 37156 11956 43148
rect 11900 37090 11956 37100
rect 11676 32722 11732 32732
rect 11452 25554 11508 25564
rect 12012 22932 12068 44940
rect 12348 43876 12404 43886
rect 12348 43540 12404 43820
rect 12348 43474 12404 43484
rect 12348 38276 12404 38286
rect 12348 37828 12404 38220
rect 12348 31668 12404 37772
rect 12348 31602 12404 31612
rect 12460 29428 12516 52220
rect 12572 48244 12628 53452
rect 12684 52276 12740 53676
rect 13468 53620 13524 53630
rect 12684 52210 12740 52220
rect 13132 52948 13188 52958
rect 12572 48178 12628 48188
rect 12796 46004 12852 46014
rect 12684 43988 12740 43998
rect 12572 43764 12628 43774
rect 12684 43764 12740 43932
rect 12628 43708 12740 43764
rect 12572 43698 12628 43708
rect 12796 32788 12852 45948
rect 12796 32722 12852 32732
rect 12460 28868 12516 29372
rect 12460 28802 12516 28812
rect 12012 22866 12068 22876
rect 13132 21812 13188 52892
rect 13356 50484 13412 50494
rect 13468 50484 13524 53564
rect 14700 52724 14756 54684
rect 16716 54404 16772 54414
rect 14252 51492 14308 51502
rect 14028 50596 14084 50606
rect 13412 50428 13524 50484
rect 13356 50418 13412 50428
rect 13244 46676 13300 46686
rect 13244 43764 13300 46620
rect 13244 43698 13300 43708
rect 13468 42868 13524 50428
rect 13580 50484 13636 50494
rect 13580 46004 13636 50428
rect 14028 49700 14084 50540
rect 14252 50596 14308 51436
rect 14252 50530 14308 50540
rect 13580 45938 13636 45948
rect 13692 46452 13748 46462
rect 13692 44772 13748 46396
rect 13804 46340 13860 46350
rect 13804 45780 13860 46284
rect 13804 45714 13860 45724
rect 13692 44212 13748 44716
rect 14028 44548 14084 49644
rect 14700 50148 14756 52668
rect 14700 46452 14756 50092
rect 14700 46386 14756 46396
rect 14812 53732 14868 53742
rect 14812 53060 14868 53676
rect 14028 44482 14084 44492
rect 13692 43428 13748 44156
rect 13692 43362 13748 43372
rect 13468 42812 13636 42868
rect 13468 42644 13524 42654
rect 13468 38500 13524 42588
rect 13580 41860 13636 42812
rect 13580 40068 13636 41804
rect 13580 40002 13636 40012
rect 13468 38434 13524 38444
rect 13356 37268 13412 37278
rect 13356 25844 13412 37212
rect 14812 31220 14868 53004
rect 15148 52948 15204 52958
rect 14924 50372 14980 50382
rect 14924 50148 14980 50316
rect 15036 50148 15092 50158
rect 14924 50092 15036 50148
rect 15036 50082 15092 50092
rect 15148 48580 15204 52892
rect 15932 52836 15988 52846
rect 15484 51940 15540 51950
rect 15148 48514 15204 48524
rect 15260 51828 15316 51838
rect 15148 47796 15204 47806
rect 15148 42420 15204 47740
rect 15260 43652 15316 51772
rect 15484 49140 15540 51884
rect 15596 49140 15652 49150
rect 15484 49084 15596 49140
rect 15260 43586 15316 43596
rect 15372 45780 15428 45790
rect 15372 45220 15428 45724
rect 15596 45444 15652 49084
rect 15596 45378 15652 45388
rect 15708 49028 15764 49038
rect 15260 42980 15316 42990
rect 15372 42980 15428 45164
rect 15316 42924 15428 42980
rect 15260 42914 15316 42924
rect 15148 42354 15204 42364
rect 15036 41972 15092 41982
rect 15036 40852 15092 41916
rect 15036 40786 15092 40796
rect 15708 40404 15764 48972
rect 15820 46228 15876 46238
rect 15932 46228 15988 52780
rect 16492 52836 16548 52846
rect 16380 52164 16436 52174
rect 16380 51380 16436 52108
rect 16380 51314 16436 51324
rect 16492 48356 16548 52780
rect 16716 51604 16772 54348
rect 18172 54292 18228 54796
rect 18172 54226 18228 54236
rect 18284 54628 18340 54638
rect 18284 53732 18340 54572
rect 18284 53666 18340 53676
rect 16716 50428 16772 51548
rect 16604 50372 16772 50428
rect 16940 50708 16996 50718
rect 16940 50484 16996 50652
rect 16604 50036 16660 50372
rect 16604 49970 16660 49980
rect 16492 48290 16548 48300
rect 16828 49812 16884 49822
rect 16828 48356 16884 49756
rect 15876 46172 15988 46228
rect 15820 46162 15876 46172
rect 15036 40292 15092 40302
rect 15036 36148 15092 40236
rect 15036 36082 15092 36092
rect 14812 31154 14868 31164
rect 15708 30324 15764 40348
rect 15820 42644 15876 42654
rect 15820 37044 15876 42588
rect 15820 36978 15876 36988
rect 15932 31668 15988 46172
rect 16044 47236 16100 47246
rect 16044 42420 16100 47180
rect 16044 33236 16100 42364
rect 16156 46452 16212 46462
rect 16156 45892 16212 46396
rect 16156 36708 16212 45836
rect 16828 45668 16884 48300
rect 16940 45892 16996 50428
rect 17836 50708 17892 50718
rect 17836 48132 17892 50652
rect 18396 50708 18452 55580
rect 18396 50642 18452 50652
rect 17836 48066 17892 48076
rect 18284 50484 18340 50494
rect 18284 48580 18340 50428
rect 18284 47460 18340 48524
rect 18284 47394 18340 47404
rect 16940 45826 16996 45836
rect 18396 46676 18452 46686
rect 18396 45892 18452 46620
rect 16828 45612 16996 45668
rect 16716 45444 16772 45454
rect 16772 45388 16884 45444
rect 16716 45378 16772 45388
rect 16604 44100 16660 44110
rect 16604 40852 16660 44044
rect 16604 40786 16660 40796
rect 16156 36642 16212 36652
rect 16380 38948 16436 38958
rect 16380 36484 16436 38892
rect 16492 36484 16548 36494
rect 16380 36428 16492 36484
rect 16380 34916 16436 36428
rect 16492 36418 16548 36428
rect 16380 34850 16436 34860
rect 16044 33170 16100 33180
rect 16828 32788 16884 45388
rect 16940 38276 16996 45612
rect 17164 43988 17220 43998
rect 17164 41188 17220 43932
rect 17164 41122 17220 41132
rect 17724 43540 17780 43550
rect 17724 41076 17780 43484
rect 17724 41010 17780 41020
rect 16940 38210 16996 38220
rect 16828 32722 16884 32732
rect 15932 31602 15988 31612
rect 15708 30258 15764 30268
rect 18396 30212 18452 45836
rect 18396 30146 18452 30156
rect 18508 28644 18564 56028
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19068 54292 19124 54302
rect 18732 54068 18788 54078
rect 18620 49588 18676 49598
rect 18620 48132 18676 49532
rect 18620 48066 18676 48076
rect 18732 48020 18788 54012
rect 18620 45220 18676 45230
rect 18620 42308 18676 45164
rect 18620 39172 18676 42252
rect 18732 40292 18788 47964
rect 18956 46676 19012 46686
rect 18844 44772 18900 44782
rect 18844 43988 18900 44716
rect 18844 43922 18900 43932
rect 18956 44548 19012 46620
rect 18844 43652 18900 43662
rect 18844 43316 18900 43596
rect 18844 43250 18900 43260
rect 18956 42532 19012 44492
rect 18956 42466 19012 42476
rect 18732 40226 18788 40236
rect 18956 41524 19012 41534
rect 18620 39106 18676 39116
rect 18508 28578 18564 28588
rect 13356 25778 13412 25788
rect 18956 25060 19012 41468
rect 19068 36932 19124 54236
rect 19628 53620 19684 53630
rect 19628 53396 19684 53564
rect 19628 53330 19684 53340
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19404 52388 19460 52398
rect 19068 36260 19124 36876
rect 19180 44884 19236 44894
rect 19180 36372 19236 44828
rect 19404 43652 19460 52332
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19516 49924 19572 49934
rect 19516 48692 19572 49868
rect 19516 48626 19572 48636
rect 19628 49812 19684 49822
rect 19628 46788 19684 49756
rect 19628 46722 19684 46732
rect 19808 48636 20128 50148
rect 20300 52724 20356 52734
rect 20188 49924 20244 49934
rect 20188 49140 20244 49868
rect 20188 49074 20244 49084
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19404 41524 19460 43596
rect 19404 41458 19460 41468
rect 19516 46452 19572 46462
rect 19292 41188 19348 41198
rect 19292 37940 19348 41132
rect 19292 37874 19348 37884
rect 19180 36306 19236 36316
rect 19068 36194 19124 36204
rect 19516 31444 19572 46396
rect 19516 31378 19572 31388
rect 19808 45500 20128 47012
rect 20188 48692 20244 48702
rect 20188 46900 20244 48636
rect 20188 46834 20244 46844
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 20188 45556 20244 45566
rect 20188 44884 20244 45500
rect 20188 44818 20244 44828
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 20300 31892 20356 52668
rect 21308 51604 21364 57484
rect 31276 56420 31332 56430
rect 30156 55300 30212 55310
rect 22316 55076 22372 55086
rect 21308 51538 21364 51548
rect 21756 51828 21812 51838
rect 21756 49140 21812 51772
rect 21868 49364 21924 49374
rect 22092 49364 22148 49374
rect 21924 49308 22092 49364
rect 21868 49298 21924 49308
rect 22092 49298 22148 49308
rect 21756 49084 21924 49140
rect 21868 47068 21924 49084
rect 22316 48916 22372 55020
rect 26852 54964 26908 54974
rect 26796 54908 26852 54964
rect 26796 54898 26908 54908
rect 26796 54516 26852 54898
rect 30156 54740 30212 55244
rect 30156 54674 30212 54684
rect 26796 54450 26852 54460
rect 25004 53844 25060 53854
rect 24892 52052 24948 52062
rect 22316 48850 22372 48860
rect 22540 50484 22596 50494
rect 22540 48804 22596 50428
rect 23212 50260 23268 50270
rect 22540 48738 22596 48748
rect 22652 49812 22708 49822
rect 21756 47012 21812 47022
rect 21868 47012 22148 47068
rect 20524 45780 20580 45790
rect 20524 44884 20580 45724
rect 20524 44818 20580 44828
rect 20300 31826 20356 31836
rect 21196 41860 21252 41870
rect 21196 41188 21252 41804
rect 18956 24994 19012 25004
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 13132 21746 13188 21756
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 9436 21522 9492 21532
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 20412 20128 21924
rect 21196 21588 21252 41132
rect 21756 35924 21812 46956
rect 21756 35364 21812 35868
rect 21756 35298 21812 35308
rect 22092 32788 22148 47012
rect 22092 32722 22148 32732
rect 22540 42532 22596 42542
rect 22540 41636 22596 42476
rect 22540 31220 22596 41580
rect 22652 39508 22708 49756
rect 23100 49476 23156 49486
rect 23100 48468 23156 49420
rect 23212 48916 23268 50204
rect 23212 48850 23268 48860
rect 24668 49140 24724 49150
rect 23100 48402 23156 48412
rect 24668 46340 24724 49084
rect 24892 47124 24948 51996
rect 25004 47460 25060 53788
rect 27020 50484 27076 50494
rect 27020 48916 27076 50428
rect 27020 48850 27076 48860
rect 31164 49252 31220 49262
rect 25004 47394 25060 47404
rect 24892 47058 24948 47068
rect 24668 46274 24724 46284
rect 22652 39442 22708 39452
rect 23100 44100 23156 44110
rect 23100 36372 23156 44044
rect 29596 44100 29652 44110
rect 26796 42756 26852 42766
rect 25228 42196 25284 42206
rect 25228 41076 25284 42140
rect 25228 41010 25284 41020
rect 26796 40628 26852 42700
rect 26796 40562 26852 40572
rect 23100 36306 23156 36316
rect 29596 36260 29652 44044
rect 31164 40516 31220 49196
rect 31164 40450 31220 40460
rect 31052 38724 31108 38734
rect 31052 38052 31108 38668
rect 31052 37986 31108 37996
rect 29596 36194 29652 36204
rect 31164 34020 31220 34030
rect 22540 31154 22596 31164
rect 30828 33348 30884 33358
rect 30828 25060 30884 33292
rect 31164 33236 31220 33964
rect 31164 33170 31220 33180
rect 31276 28868 31332 56364
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 32396 55412 32452 55422
rect 32396 47572 32452 55356
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 33740 51716 33796 51726
rect 33740 51268 33796 51660
rect 33740 51202 33796 51212
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 33964 49700 34020 49710
rect 32396 47506 32452 47516
rect 33068 47572 33124 47582
rect 32844 47460 32900 47470
rect 32844 47124 32900 47404
rect 32844 47058 32900 47068
rect 33068 47124 33124 47516
rect 33068 47058 33124 47068
rect 32060 46564 32116 46574
rect 31612 45892 31668 45902
rect 31612 44772 31668 45836
rect 31612 44706 31668 44716
rect 32060 30548 32116 46508
rect 32060 30482 32116 30492
rect 32732 46564 32788 46574
rect 31276 28802 31332 28812
rect 30828 24994 30884 25004
rect 32732 24612 32788 46508
rect 33740 46004 33796 46014
rect 33740 36148 33796 45948
rect 33740 36082 33796 36092
rect 32732 24546 32788 24556
rect 33964 23380 34020 49644
rect 35168 49420 35488 50932
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 36764 49476 36820 49486
rect 35756 48804 35812 48814
rect 34300 47796 34356 47806
rect 34300 47348 34356 47740
rect 34300 47282 34356 47292
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 34524 45108 34580 45118
rect 34076 35700 34132 35710
rect 34076 35476 34132 35644
rect 34076 35410 34132 35420
rect 34188 24388 34244 24398
rect 34188 23604 34244 24332
rect 34188 23538 34244 23548
rect 33964 23314 34020 23324
rect 34524 21700 34580 45052
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 34860 42756 34916 42766
rect 34860 42532 34916 42700
rect 34860 42466 34916 42476
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 34524 21634 34580 21644
rect 34748 23940 34804 23950
rect 21196 21522 21252 21532
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 34300 19572 34356 19582
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 33964 18340 34020 18350
rect 27916 15540 27972 15550
rect 27916 15316 27972 15484
rect 27916 15250 27972 15260
rect 33964 14308 34020 18284
rect 34300 16548 34356 19516
rect 34524 17220 34580 17230
rect 34524 16884 34580 17164
rect 34524 16818 34580 16828
rect 34300 16482 34356 16492
rect 33964 14242 34020 14252
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 34748 13972 34804 23884
rect 34748 13906 34804 13916
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35644 48132 35700 48142
rect 35644 20692 35700 48076
rect 35756 35140 35812 48748
rect 36764 47908 36820 49420
rect 36764 47842 36820 47852
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 38108 47348 38164 47358
rect 38108 46452 38164 47292
rect 38108 46386 38164 46396
rect 43372 47348 43428 47358
rect 35868 44660 35924 44670
rect 35868 37044 35924 44604
rect 35868 36978 35924 36988
rect 35756 35074 35812 35084
rect 42924 27748 42980 27758
rect 42924 27524 42980 27692
rect 41356 26964 41412 26974
rect 36316 26852 36372 26862
rect 36316 23156 36372 26796
rect 38668 25620 38724 25630
rect 38556 25284 38612 25294
rect 38668 25284 38724 25564
rect 38612 25228 38724 25284
rect 38556 25218 38612 25228
rect 36540 24500 36596 24510
rect 36540 23940 36596 24444
rect 36540 23874 36596 23884
rect 36316 23090 36372 23100
rect 38780 22932 38836 22942
rect 35644 20626 35700 20636
rect 35756 22148 35812 22158
rect 35756 20244 35812 22092
rect 35756 20178 35812 20188
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 38108 20020 38164 20030
rect 38108 19572 38164 19964
rect 38108 19506 38164 19516
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 38780 17892 38836 22876
rect 41020 21476 41076 21486
rect 41020 21028 41076 21420
rect 41356 21140 41412 26908
rect 41468 26180 41524 26190
rect 41468 24612 41524 26124
rect 41468 24052 41524 24556
rect 41468 23986 41524 23996
rect 41356 21074 41412 21084
rect 42028 23716 42084 23726
rect 41020 20962 41076 20972
rect 39452 20356 39508 20366
rect 39452 19796 39508 20300
rect 39452 19730 39508 19740
rect 40684 19796 40740 19806
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 36204 16996 36260 17006
rect 36204 16324 36260 16940
rect 36540 16884 36596 16894
rect 36540 16660 36596 16828
rect 38780 16772 38836 17836
rect 38780 16706 38836 16716
rect 39228 19572 39284 19582
rect 36540 16594 36596 16604
rect 36204 16258 36260 16268
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 39116 16100 39172 16110
rect 39116 12628 39172 16044
rect 39228 14532 39284 19516
rect 39228 13636 39284 14476
rect 39228 13570 39284 13580
rect 39452 18228 39508 18238
rect 39452 13076 39508 18172
rect 40236 15652 40292 15662
rect 39900 14644 39956 14654
rect 39900 13748 39956 14588
rect 39900 13682 39956 13692
rect 39452 13010 39508 13020
rect 39116 12562 39172 12572
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 25564 10276 25620 10286
rect 25564 9828 25620 10220
rect 25564 9762 25620 9772
rect 35168 10220 35488 11732
rect 38668 11732 38724 11742
rect 38668 10948 38724 11676
rect 38668 10882 38724 10892
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 40236 2548 40292 15596
rect 40684 13524 40740 19740
rect 41468 19796 41524 19806
rect 41468 15876 41524 19740
rect 41468 15810 41524 15820
rect 40684 13458 40740 13468
rect 41580 14644 41636 14654
rect 41580 13412 41636 14588
rect 41580 13346 41636 13356
rect 42028 8036 42084 23660
rect 42140 20580 42196 20590
rect 42140 14084 42196 20524
rect 42252 20244 42308 20254
rect 42252 20020 42308 20188
rect 42252 19954 42308 19964
rect 42252 18676 42308 18686
rect 42252 18228 42308 18620
rect 42252 18162 42308 18172
rect 42812 18116 42868 18126
rect 42812 16660 42868 18060
rect 42812 15428 42868 16604
rect 42924 16324 42980 27468
rect 42924 16258 42980 16268
rect 43148 17332 43204 17342
rect 42812 15362 42868 15372
rect 43148 14532 43204 17276
rect 43148 14466 43204 14476
rect 42140 14018 42196 14028
rect 42700 12516 42756 12526
rect 42700 11172 42756 12460
rect 42700 11106 42756 11116
rect 42028 7970 42084 7980
rect 43372 2660 43428 47292
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50092 34580 50148 34590
rect 46396 32116 46452 32126
rect 46396 31556 46452 32060
rect 46284 29988 46340 29998
rect 44492 26964 44548 26974
rect 44492 26740 44548 26908
rect 44492 26674 44548 26684
rect 44156 26068 44212 26078
rect 43932 21700 43988 21710
rect 43596 20916 43652 20926
rect 43596 20020 43652 20860
rect 43708 20020 43764 20030
rect 43596 19964 43708 20020
rect 43708 19954 43764 19964
rect 43708 19236 43764 19246
rect 43596 17108 43652 17118
rect 43484 16100 43540 16110
rect 43484 14980 43540 16044
rect 43484 14914 43540 14924
rect 43596 15316 43652 17052
rect 43708 15652 43764 19180
rect 43932 18676 43988 21644
rect 43932 18610 43988 18620
rect 43708 15586 43764 15596
rect 43708 15316 43764 15326
rect 43596 15260 43708 15316
rect 43596 11284 43652 15260
rect 43708 15250 43764 15260
rect 44156 12852 44212 26012
rect 45612 25508 45668 25518
rect 45388 24612 45444 24622
rect 44268 19908 44324 19918
rect 44268 17332 44324 19852
rect 45276 19572 45332 19582
rect 45276 18564 45332 19516
rect 45276 18498 45332 18508
rect 44268 17266 44324 17276
rect 44156 11844 44212 12796
rect 44156 11778 44212 11788
rect 43596 11218 43652 11228
rect 45388 8484 45444 24556
rect 45500 23044 45556 23054
rect 45500 16548 45556 22988
rect 45612 21588 45668 25452
rect 45612 19796 45668 21532
rect 45612 17108 45668 19740
rect 46172 23156 46228 23166
rect 45948 19124 46004 19134
rect 45612 17042 45668 17052
rect 45724 18900 45780 18910
rect 45500 16482 45556 16492
rect 45724 13524 45780 18844
rect 45948 14756 46004 19068
rect 46172 18228 46228 23100
rect 46284 20804 46340 29932
rect 46284 20738 46340 20748
rect 45948 14690 46004 14700
rect 46060 17332 46116 17342
rect 46060 16212 46116 17276
rect 45724 13458 45780 13468
rect 46060 13076 46116 16156
rect 46172 16100 46228 18172
rect 46172 16034 46228 16044
rect 46060 13010 46116 13020
rect 46396 11956 46452 31500
rect 49756 32004 49812 32014
rect 49532 31108 49588 31118
rect 47068 29204 47124 29214
rect 46956 28980 47012 28990
rect 46508 24388 46564 24398
rect 46508 19684 46564 24332
rect 46956 23380 47012 28924
rect 47068 27636 47124 29148
rect 47068 27570 47124 27580
rect 48636 27636 48692 27646
rect 48412 27412 48468 27422
rect 46956 23314 47012 23324
rect 47404 26404 47460 26414
rect 46956 22932 47012 22942
rect 46956 21588 47012 22876
rect 46956 21522 47012 21532
rect 46508 19618 46564 19628
rect 47068 20692 47124 20702
rect 47068 19572 47124 20636
rect 47068 15988 47124 19516
rect 47068 15922 47124 15932
rect 47180 16324 47236 16334
rect 47180 15148 47236 16268
rect 46396 11890 46452 11900
rect 47068 15092 47236 15148
rect 47404 15204 47460 26348
rect 47964 23828 48020 23838
rect 47964 23604 48020 23772
rect 47404 15138 47460 15148
rect 47516 17220 47572 17230
rect 47068 13748 47124 15092
rect 47068 9716 47124 13692
rect 47516 12068 47572 17164
rect 47964 13524 48020 23548
rect 48300 21812 48356 21822
rect 47964 13458 48020 13468
rect 48188 19124 48244 19134
rect 47516 12002 47572 12012
rect 48188 12068 48244 19068
rect 48300 16324 48356 21756
rect 48300 16258 48356 16268
rect 48412 18676 48468 27356
rect 48636 27412 48692 27580
rect 48636 27346 48692 27356
rect 49308 26964 49364 26974
rect 48748 26180 48804 26190
rect 48636 25844 48692 25854
rect 48636 25396 48692 25788
rect 48636 20692 48692 25340
rect 48748 24612 48804 26124
rect 48748 23548 48804 24556
rect 48748 23492 49028 23548
rect 48972 23156 49028 23492
rect 48748 22932 48804 22942
rect 48748 21252 48804 22876
rect 48748 21186 48804 21196
rect 48860 22372 48916 22382
rect 48860 21476 48916 22316
rect 48636 20626 48692 20636
rect 48748 20580 48804 20590
rect 48412 15988 48468 18620
rect 48524 20020 48580 20030
rect 48524 18228 48580 19964
rect 48636 18564 48692 18574
rect 48748 18564 48804 20524
rect 48860 20468 48916 21420
rect 48860 20402 48916 20412
rect 48692 18508 48804 18564
rect 48636 18498 48692 18508
rect 48524 18162 48580 18172
rect 48412 15922 48468 15932
rect 48188 9828 48244 12012
rect 48636 15428 48692 15438
rect 48636 10164 48692 15372
rect 48636 10098 48692 10108
rect 48748 11396 48804 18508
rect 48972 19012 49028 23100
rect 49196 23380 49252 23390
rect 49084 23044 49140 23054
rect 49084 19908 49140 22988
rect 49196 21588 49252 23324
rect 49196 21522 49252 21532
rect 49084 19842 49140 19852
rect 48972 18564 49028 18956
rect 48972 18498 49028 18508
rect 49196 19572 49252 19582
rect 49196 18788 49252 19516
rect 48860 18340 48916 18350
rect 48860 15652 48916 18284
rect 48860 15586 48916 15596
rect 49196 11508 49252 18732
rect 49308 13636 49364 26908
rect 49532 22932 49588 31052
rect 49532 22866 49588 22876
rect 49644 27412 49700 27422
rect 49644 21812 49700 27356
rect 49644 21746 49700 21756
rect 49644 18452 49700 18462
rect 49308 13570 49364 13580
rect 49532 16660 49588 16670
rect 49420 12180 49476 12190
rect 49420 11844 49476 12124
rect 49420 11778 49476 11788
rect 49196 11442 49252 11452
rect 48188 9762 48244 9772
rect 47068 9650 47124 9660
rect 45388 8418 45444 8428
rect 47180 8260 47236 8270
rect 47180 8036 47236 8204
rect 47180 7970 47236 7980
rect 43372 2594 43428 2604
rect 40236 2482 40292 2492
rect 48748 1540 48804 11340
rect 49532 10836 49588 16604
rect 49644 15652 49700 18396
rect 49756 18228 49812 31948
rect 49980 21140 50036 21150
rect 49980 19460 50036 21084
rect 49980 19394 50036 19404
rect 49756 17556 49812 18172
rect 49756 17490 49812 17500
rect 49644 15586 49700 15596
rect 49756 16436 49812 16446
rect 49756 15988 49812 16380
rect 49532 10770 49588 10780
rect 49644 11172 49700 11182
rect 49644 3108 49700 11116
rect 49756 8148 49812 15932
rect 49980 16100 50036 16110
rect 49980 11284 50036 16044
rect 50092 14532 50148 34524
rect 50528 34524 50848 36036
rect 54908 37044 54964 37054
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 54796 34692 54852 34702
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50316 30996 50372 31006
rect 50316 27636 50372 30940
rect 50316 26964 50372 27580
rect 50316 24052 50372 26908
rect 50316 23986 50372 23996
rect 50528 29820 50848 31332
rect 53564 31892 53620 31902
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50204 23268 50260 23278
rect 50204 22148 50260 23212
rect 50204 16212 50260 22092
rect 50316 22036 50372 22046
rect 50316 21700 50372 21980
rect 50316 21634 50372 21644
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 51436 30548 51492 30558
rect 51436 29204 51492 30492
rect 50204 15764 50260 16156
rect 50204 15698 50260 15708
rect 50316 21476 50372 21486
rect 50316 20916 50372 21420
rect 50316 20692 50372 20860
rect 50092 14466 50148 14476
rect 50204 15092 50260 15102
rect 50204 14644 50260 15036
rect 49980 10612 50036 11228
rect 49980 10546 50036 10556
rect 49756 8082 49812 8092
rect 50204 6468 50260 14588
rect 50316 11620 50372 20636
rect 50316 11554 50372 11564
rect 50528 20412 50848 21924
rect 51324 21924 51380 21934
rect 51212 21812 51268 21822
rect 51100 21588 51156 21598
rect 51100 21364 51156 21532
rect 51212 21476 51268 21756
rect 51212 21410 51268 21420
rect 51100 21298 51156 21308
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50988 21028 51044 21038
rect 50988 19460 51044 20972
rect 50988 19394 51044 19404
rect 51100 20132 51156 20142
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 51100 19124 51156 20076
rect 51212 20020 51268 20030
rect 51212 19460 51268 19964
rect 51212 19394 51268 19404
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50988 18452 51044 18462
rect 50988 17556 51044 18396
rect 50988 14868 51044 17500
rect 51100 16100 51156 19068
rect 51100 16034 51156 16044
rect 51212 19236 51268 19246
rect 50988 14802 51044 14812
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50204 6402 50260 6412
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50988 13636 51044 13646
rect 50988 12628 51044 13580
rect 50988 10388 51044 12572
rect 50988 10322 51044 10332
rect 51100 13076 51156 13086
rect 51100 12180 51156 13020
rect 51212 12404 51268 19180
rect 51324 18116 51380 21868
rect 51324 18050 51380 18060
rect 51436 16324 51492 29148
rect 53452 27748 53508 27758
rect 51772 24500 51828 24510
rect 51548 22148 51604 22158
rect 51548 21476 51604 22092
rect 51548 21410 51604 21420
rect 51660 19460 51716 19470
rect 51212 12338 51268 12348
rect 51324 14756 51380 14766
rect 51212 12180 51268 12190
rect 51100 12124 51212 12180
rect 51100 10164 51156 12124
rect 51212 12114 51268 12124
rect 51324 12068 51380 14700
rect 51324 12002 51380 12012
rect 51100 10098 51156 10108
rect 51436 10164 51492 16268
rect 51548 19124 51604 19134
rect 51548 15652 51604 19068
rect 51660 15764 51716 19404
rect 51772 19236 51828 24444
rect 53452 23940 53508 27692
rect 53452 23874 53508 23884
rect 53340 22148 53396 22158
rect 52108 21700 52164 21710
rect 52108 20132 52164 21644
rect 53228 21476 53284 21486
rect 52668 21364 52724 21374
rect 52108 20066 52164 20076
rect 52220 20468 52276 20478
rect 51772 19170 51828 19180
rect 51884 19908 51940 19918
rect 51772 17780 51828 17790
rect 51772 16772 51828 17724
rect 51884 17332 51940 19852
rect 51884 17266 51940 17276
rect 51996 19348 52052 19358
rect 51996 19012 52052 19292
rect 51772 16706 51828 16716
rect 51996 17220 52052 18956
rect 51660 15698 51716 15708
rect 51772 16100 51828 16110
rect 51548 15316 51604 15596
rect 51548 15250 51604 15260
rect 51436 10098 51492 10108
rect 51548 14196 51604 14206
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 51548 7028 51604 14140
rect 51772 12180 51828 16044
rect 51996 14420 52052 17164
rect 51884 14084 51940 14094
rect 51884 13748 51940 14028
rect 51884 13682 51940 13692
rect 51772 12114 51828 12124
rect 51996 10052 52052 14364
rect 52220 13412 52276 20412
rect 52332 18004 52388 18014
rect 52332 14756 52388 17948
rect 52332 14690 52388 14700
rect 52220 13346 52276 13356
rect 52444 14196 52500 14206
rect 51996 9986 52052 9996
rect 51548 6962 51604 6972
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 52444 6020 52500 14140
rect 52668 13076 52724 21308
rect 53228 21252 53284 21420
rect 53228 18004 53284 21196
rect 53228 17938 53284 17948
rect 53340 14196 53396 22092
rect 53452 20356 53508 20366
rect 53452 15204 53508 20300
rect 53452 15138 53508 15148
rect 53340 14130 53396 14140
rect 52668 13010 52724 13020
rect 53452 12852 53508 12862
rect 53452 12068 53508 12796
rect 53452 12002 53508 12012
rect 53564 8260 53620 31836
rect 53676 26516 53732 26526
rect 53676 23828 53732 26460
rect 53676 23156 53732 23772
rect 53676 22148 53732 23100
rect 53676 22082 53732 22092
rect 53900 23716 53956 23726
rect 53676 20132 53732 20142
rect 53676 18452 53732 20076
rect 53900 18788 53956 23660
rect 53900 18722 53956 18732
rect 54460 18564 54516 18574
rect 53676 11844 53732 18396
rect 53900 18452 53956 18462
rect 53900 12180 53956 18396
rect 54012 17108 54068 17118
rect 54012 15988 54068 17052
rect 54460 16324 54516 18508
rect 54796 17668 54852 34636
rect 54796 17602 54852 17612
rect 54460 16258 54516 16268
rect 54012 15922 54068 15932
rect 54572 15540 54628 15550
rect 53900 12114 53956 12124
rect 54460 15428 54516 15438
rect 53676 11778 53732 11788
rect 54460 11844 54516 15372
rect 54460 11778 54516 11788
rect 53564 8194 53620 8204
rect 54572 6692 54628 15484
rect 54908 13076 54964 36988
rect 55244 29876 55300 29886
rect 54908 13010 54964 13020
rect 55020 23044 55076 23054
rect 55020 12964 55076 22988
rect 55244 20020 55300 29820
rect 55692 25172 55748 25182
rect 55020 12898 55076 12908
rect 55132 17668 55188 17678
rect 55132 9268 55188 17612
rect 55244 9940 55300 19964
rect 55356 22932 55412 22942
rect 55356 22148 55412 22876
rect 55356 19572 55412 22092
rect 55356 19506 55412 19516
rect 55580 20580 55636 20590
rect 55468 19460 55524 19470
rect 55356 19348 55412 19358
rect 55356 18900 55412 19292
rect 55356 18834 55412 18844
rect 55468 18452 55524 19404
rect 55468 18386 55524 18396
rect 55580 18228 55636 20524
rect 55580 13636 55636 18172
rect 55580 13570 55636 13580
rect 55692 15204 55748 25116
rect 55916 20244 55972 20254
rect 55244 9874 55300 9884
rect 55132 9202 55188 9212
rect 54572 6626 54628 6636
rect 55692 6580 55748 15148
rect 55804 15876 55860 15886
rect 55804 13076 55860 15820
rect 55916 13524 55972 20188
rect 56028 19684 56084 19694
rect 56028 15876 56084 19628
rect 56028 15810 56084 15820
rect 56476 18452 56532 18462
rect 55916 13458 55972 13468
rect 55804 13010 55860 13020
rect 56476 9604 56532 18396
rect 56812 16548 56868 16558
rect 56700 16100 56756 16110
rect 56700 15428 56756 16044
rect 56700 15362 56756 15372
rect 56476 9538 56532 9548
rect 56812 6692 56868 16492
rect 57148 14420 57204 14430
rect 57148 12516 57204 14364
rect 57148 12450 57204 12460
rect 56812 6626 56868 6636
rect 55692 6514 55748 6524
rect 52444 5954 52500 5964
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 49644 3042 49700 3052
rect 48748 1474 48804 1484
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1346__I dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 57792 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1347__I
timestamp 1669390400
transform 1 0 56672 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__A2
timestamp 1669390400
transform -1 0 57568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1350__I
timestamp 1669390400
transform 1 0 55328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1352__I
timestamp 1669390400
transform 1 0 53872 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1354__I
timestamp 1669390400
transform 1 0 51072 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__A3
timestamp 1669390400
transform 1 0 52528 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1358__A1
timestamp 1669390400
transform 1 0 32592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1358__A2
timestamp 1669390400
transform -1 0 33264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1359__I
timestamp 1669390400
transform 1 0 51072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1360__I
timestamp 1669390400
transform -1 0 53984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__A1
timestamp 1669390400
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__B
timestamp 1669390400
transform 1 0 32368 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1364__I
timestamp 1669390400
transform 1 0 50288 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1366__I
timestamp 1669390400
transform 1 0 57120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1367__A3
timestamp 1669390400
transform -1 0 57008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1367__B
timestamp 1669390400
transform 1 0 57680 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1368__A1
timestamp 1669390400
transform -1 0 51856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1368__A2
timestamp 1669390400
transform -1 0 52192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1370__I
timestamp 1669390400
transform -1 0 58016 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1371__I
timestamp 1669390400
transform 1 0 57344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1372__I
timestamp 1669390400
transform 1 0 54992 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1373__I
timestamp 1669390400
transform 1 0 58016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1374__A1
timestamp 1669390400
transform 1 0 57792 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__A1
timestamp 1669390400
transform -1 0 56896 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1375__A4
timestamp 1669390400
transform -1 0 56896 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1376__A1
timestamp 1669390400
transform -1 0 35280 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1376__A2
timestamp 1669390400
transform 1 0 33264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1377__A2
timestamp 1669390400
transform 1 0 28672 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1380__I
timestamp 1669390400
transform 1 0 55664 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1381__I
timestamp 1669390400
transform 1 0 55328 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1384__A1
timestamp 1669390400
transform 1 0 57344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1384__A3
timestamp 1669390400
transform 1 0 57792 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1385__A1
timestamp 1669390400
transform 1 0 36736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1385__A2
timestamp 1669390400
transform 1 0 39312 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1386__A2
timestamp 1669390400
transform 1 0 28000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1388__I
timestamp 1669390400
transform 1 0 21840 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1389__I
timestamp 1669390400
transform 1 0 9632 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1392__I
timestamp 1669390400
transform 1 0 9632 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1393__I
timestamp 1669390400
transform 1 0 5488 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1397__I
timestamp 1669390400
transform 1 0 20832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1400__A3
timestamp 1669390400
transform 1 0 8512 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1401__A1
timestamp 1669390400
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1402__I
timestamp 1669390400
transform 1 0 19712 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1403__I
timestamp 1669390400
transform 1 0 2352 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1405__A1
timestamp 1669390400
transform 1 0 5712 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1405__A2
timestamp 1669390400
transform 1 0 8848 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1406__A2
timestamp 1669390400
transform 1 0 19040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1407__A1
timestamp 1669390400
transform 1 0 24080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1407__A2
timestamp 1669390400
transform 1 0 22064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1408__I
timestamp 1669390400
transform 1 0 25536 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__A2
timestamp 1669390400
transform 1 0 20160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1410__I
timestamp 1669390400
transform 1 0 12320 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1411__A1
timestamp 1669390400
transform 1 0 11872 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1412__A1
timestamp 1669390400
transform 1 0 12544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1412__A2
timestamp 1669390400
transform 1 0 14336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1413__A2
timestamp 1669390400
transform 1 0 25984 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1414__B
timestamp 1669390400
transform 1 0 25984 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1415__A1
timestamp 1669390400
transform -1 0 24192 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1415__A2
timestamp 1669390400
transform 1 0 23184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1415__A3
timestamp 1669390400
transform 1 0 25536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1416__I
timestamp 1669390400
transform -1 0 30688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1419__A2
timestamp 1669390400
transform 1 0 26096 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1420__I
timestamp 1669390400
transform 1 0 25536 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1422__A1
timestamp 1669390400
transform 1 0 26656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1425__I
timestamp 1669390400
transform -1 0 30016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1427__I
timestamp 1669390400
transform 1 0 26544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1428__I
timestamp 1669390400
transform 1 0 26096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1430__A2
timestamp 1669390400
transform -1 0 27664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1431__A1
timestamp 1669390400
transform 1 0 26432 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1431__A2
timestamp 1669390400
transform 1 0 27888 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1432__A1
timestamp 1669390400
transform -1 0 24864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1433__A1
timestamp 1669390400
transform -1 0 22624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1434__I
timestamp 1669390400
transform 1 0 31136 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1436__I
timestamp 1669390400
transform 1 0 27888 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1437__I
timestamp 1669390400
transform 1 0 30016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1438__A1
timestamp 1669390400
transform -1 0 31248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1439__A1
timestamp 1669390400
transform 1 0 27776 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1439__A2
timestamp 1669390400
transform -1 0 29344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1440__A1
timestamp 1669390400
transform 1 0 28672 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__A1
timestamp 1669390400
transform -1 0 31472 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__A2
timestamp 1669390400
transform 1 0 29344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1442__A1
timestamp 1669390400
transform 1 0 18480 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1442__A2
timestamp 1669390400
transform 1 0 16912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1444__A1
timestamp 1669390400
transform 1 0 20832 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1444__A2
timestamp 1669390400
transform 1 0 20384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1446__I
timestamp 1669390400
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1448__A2
timestamp 1669390400
transform -1 0 26768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1449__I
timestamp 1669390400
transform 1 0 31024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1450__I
timestamp 1669390400
transform 1 0 30240 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__I
timestamp 1669390400
transform -1 0 36400 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1452__I
timestamp 1669390400
transform 1 0 20384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1454__I
timestamp 1669390400
transform -1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1458__I
timestamp 1669390400
transform 1 0 24976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1459__A1
timestamp 1669390400
transform 1 0 15904 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1460__I
timestamp 1669390400
transform -1 0 2128 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__I
timestamp 1669390400
transform -1 0 7952 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1463__A1
timestamp 1669390400
transform 1 0 16912 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1463__B
timestamp 1669390400
transform -1 0 16688 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1464__I
timestamp 1669390400
transform 1 0 6384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1467__I
timestamp 1669390400
transform -1 0 4144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1469__I
timestamp 1669390400
transform -1 0 4032 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1472__A1
timestamp 1669390400
transform -1 0 4592 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1472__A2
timestamp 1669390400
transform -1 0 2464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1472__C
timestamp 1669390400
transform 1 0 5824 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1473__I
timestamp 1669390400
transform -1 0 14672 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__A2
timestamp 1669390400
transform 1 0 7728 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1476__I
timestamp 1669390400
transform 1 0 17584 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__A1
timestamp 1669390400
transform 1 0 17920 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__A2
timestamp 1669390400
transform 1 0 16912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__I
timestamp 1669390400
transform -1 0 16240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1481__I
timestamp 1669390400
transform 1 0 4144 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1482__I
timestamp 1669390400
transform -1 0 3808 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1485__I
timestamp 1669390400
transform -1 0 2016 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1486__I
timestamp 1669390400
transform 1 0 4592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__A2
timestamp 1669390400
transform 1 0 5936 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__B
timestamp 1669390400
transform 1 0 4480 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__A1
timestamp 1669390400
transform 1 0 19264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__A2
timestamp 1669390400
transform 1 0 20832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1489__A1
timestamp 1669390400
transform 1 0 18816 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1489__A3
timestamp 1669390400
transform 1 0 20608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1489__B2
timestamp 1669390400
transform -1 0 20048 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1493__A1
timestamp 1669390400
transform 1 0 21616 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1493__A2
timestamp 1669390400
transform 1 0 22064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__A1
timestamp 1669390400
transform 1 0 20272 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__A2
timestamp 1669390400
transform 1 0 20720 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__B
timestamp 1669390400
transform -1 0 22176 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1497__A1
timestamp 1669390400
transform -1 0 28112 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1498__I
timestamp 1669390400
transform -1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1499__I
timestamp 1669390400
transform -1 0 16576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1500__A2
timestamp 1669390400
transform 1 0 15232 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__A1
timestamp 1669390400
transform -1 0 8400 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__A2
timestamp 1669390400
transform 1 0 8624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__B
timestamp 1669390400
transform 1 0 5600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1504__I
timestamp 1669390400
transform 1 0 7168 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__A2
timestamp 1669390400
transform 1 0 11200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A2
timestamp 1669390400
transform 1 0 16016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__B1
timestamp 1669390400
transform -1 0 15792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__B2
timestamp 1669390400
transform 1 0 15568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__A1
timestamp 1669390400
transform 1 0 7280 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__A2
timestamp 1669390400
transform 1 0 12208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__A2
timestamp 1669390400
transform 1 0 9744 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1514__B
timestamp 1669390400
transform 1 0 11872 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1515__A1
timestamp 1669390400
transform 1 0 4592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1516__A2
timestamp 1669390400
transform -1 0 17808 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__I
timestamp 1669390400
transform -1 0 5824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__A1
timestamp 1669390400
transform -1 0 2016 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__A3
timestamp 1669390400
transform -1 0 2464 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1523__B
timestamp 1669390400
transform -1 0 5152 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__A1
timestamp 1669390400
transform -1 0 2464 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__A2
timestamp 1669390400
transform -1 0 2464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__A3
timestamp 1669390400
transform -1 0 1904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__B1
timestamp 1669390400
transform 1 0 19488 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__B2
timestamp 1669390400
transform -1 0 15792 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__A2
timestamp 1669390400
transform 1 0 37184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1527__I
timestamp 1669390400
transform -1 0 36960 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1529__A1
timestamp 1669390400
transform 1 0 30016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1529__A2
timestamp 1669390400
transform -1 0 32032 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1532__I
timestamp 1669390400
transform -1 0 15344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1533__I
timestamp 1669390400
transform 1 0 3136 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1535__A1
timestamp 1669390400
transform 1 0 12432 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1535__A2
timestamp 1669390400
transform 1 0 11648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1535__B
timestamp 1669390400
transform -1 0 14672 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1536__I0
timestamp 1669390400
transform 1 0 8064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1536__I1
timestamp 1669390400
transform 1 0 8400 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1537__A2
timestamp 1669390400
transform 1 0 9856 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1538__I
timestamp 1669390400
transform 1 0 12432 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1541__A1
timestamp 1669390400
transform -1 0 15680 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1541__A2
timestamp 1669390400
transform 1 0 12880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1542__A1
timestamp 1669390400
transform -1 0 15792 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1542__B1
timestamp 1669390400
transform 1 0 15008 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1542__B2
timestamp 1669390400
transform 1 0 9184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1544__A1
timestamp 1669390400
transform 1 0 3584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1545__A1
timestamp 1669390400
transform 1 0 6384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__A1
timestamp 1669390400
transform 1 0 5600 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__A2
timestamp 1669390400
transform -1 0 6384 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__B
timestamp 1669390400
transform -1 0 2016 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1547__A1
timestamp 1669390400
transform -1 0 1904 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1547__A3
timestamp 1669390400
transform 1 0 5152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1550__A1
timestamp 1669390400
transform -1 0 18816 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__A1
timestamp 1669390400
transform 1 0 18368 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__A2
timestamp 1669390400
transform 1 0 17920 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__B
timestamp 1669390400
transform 1 0 16912 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__C
timestamp 1669390400
transform 1 0 17472 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__A1
timestamp 1669390400
transform 1 0 22624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__A3
timestamp 1669390400
transform 1 0 24416 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1553__A2
timestamp 1669390400
transform -1 0 21056 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1553__B
timestamp 1669390400
transform 1 0 24080 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1553__C
timestamp 1669390400
transform 1 0 24976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1557__I
timestamp 1669390400
transform -1 0 3360 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__A2
timestamp 1669390400
transform 1 0 33936 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1563__A1
timestamp 1669390400
transform 1 0 25424 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1563__A2
timestamp 1669390400
transform 1 0 22624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1564__A2
timestamp 1669390400
transform -1 0 5040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1565__A1
timestamp 1669390400
transform 1 0 7616 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__A2
timestamp 1669390400
transform -1 0 15008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1567__A1
timestamp 1669390400
transform -1 0 18816 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1567__B1
timestamp 1669390400
transform -1 0 17136 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1567__C
timestamp 1669390400
transform 1 0 16016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1570__A1
timestamp 1669390400
transform -1 0 2016 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1570__A2
timestamp 1669390400
transform -1 0 2464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__A2
timestamp 1669390400
transform -1 0 2912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1573__A2
timestamp 1669390400
transform -1 0 4368 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1573__B
timestamp 1669390400
transform -1 0 3136 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1575__B
timestamp 1669390400
transform 1 0 4368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A2
timestamp 1669390400
transform -1 0 10416 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__B
timestamp 1669390400
transform -1 0 11984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1577__A1
timestamp 1669390400
transform -1 0 12096 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1577__A2
timestamp 1669390400
transform 1 0 12880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1577__B
timestamp 1669390400
transform 1 0 15568 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1578__I
timestamp 1669390400
transform -1 0 11536 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__A1
timestamp 1669390400
transform -1 0 9968 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__B2
timestamp 1669390400
transform -1 0 7056 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A1
timestamp 1669390400
transform 1 0 30464 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A2
timestamp 1669390400
transform 1 0 33488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1582__A1
timestamp 1669390400
transform -1 0 33264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1583__I
timestamp 1669390400
transform -1 0 12992 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1584__I
timestamp 1669390400
transform -1 0 2016 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1585__A1
timestamp 1669390400
transform -1 0 2240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1585__A2
timestamp 1669390400
transform -1 0 2688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1586__I
timestamp 1669390400
transform 1 0 35728 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1587__A1
timestamp 1669390400
transform -1 0 4592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__A1
timestamp 1669390400
transform -1 0 12208 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__A2
timestamp 1669390400
transform -1 0 15008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__A3
timestamp 1669390400
transform -1 0 14112 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1589__I
timestamp 1669390400
transform 1 0 2240 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1590__A1
timestamp 1669390400
transform -1 0 10080 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1590__A2
timestamp 1669390400
transform -1 0 12320 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1591__I
timestamp 1669390400
transform -1 0 6384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1592__A1
timestamp 1669390400
transform -1 0 10080 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1592__A2
timestamp 1669390400
transform 1 0 5824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1594__A1
timestamp 1669390400
transform 1 0 14672 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1594__A2
timestamp 1669390400
transform -1 0 6272 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1595__B
timestamp 1669390400
transform -1 0 11312 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1596__I
timestamp 1669390400
transform -1 0 5152 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A1
timestamp 1669390400
transform 1 0 14448 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A2
timestamp 1669390400
transform -1 0 18480 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1598__I
timestamp 1669390400
transform -1 0 2912 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__A1
timestamp 1669390400
transform 1 0 5936 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__A2
timestamp 1669390400
transform 1 0 5936 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1600__A2
timestamp 1669390400
transform 1 0 24864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1601__I
timestamp 1669390400
transform 1 0 21840 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1602__A1
timestamp 1669390400
transform 1 0 21504 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1602__B
timestamp 1669390400
transform -1 0 20608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1602__C
timestamp 1669390400
transform 1 0 24416 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__B
timestamp 1669390400
transform 1 0 21056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1604__A1
timestamp 1669390400
transform 1 0 27888 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__A1
timestamp 1669390400
transform -1 0 26320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__I
timestamp 1669390400
transform -1 0 27216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1608__I
timestamp 1669390400
transform 1 0 19264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1609__A1
timestamp 1669390400
transform 1 0 24080 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1609__A2
timestamp 1669390400
transform 1 0 24528 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__A1
timestamp 1669390400
transform 1 0 35280 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1612__I
timestamp 1669390400
transform -1 0 3584 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__A1
timestamp 1669390400
transform 1 0 13664 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__A2
timestamp 1669390400
transform 1 0 15344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__B
timestamp 1669390400
transform 1 0 15120 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1614__I
timestamp 1669390400
transform 1 0 30240 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1615__I
timestamp 1669390400
transform 1 0 16016 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__A1
timestamp 1669390400
transform 1 0 18368 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__A2
timestamp 1669390400
transform 1 0 16912 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__B1
timestamp 1669390400
transform 1 0 25536 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1617__A1
timestamp 1669390400
transform -1 0 7728 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1617__B
timestamp 1669390400
transform -1 0 7280 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__I
timestamp 1669390400
transform 1 0 2912 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1621__I
timestamp 1669390400
transform -1 0 6160 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__A1
timestamp 1669390400
transform 1 0 7392 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__A2
timestamp 1669390400
transform 1 0 12320 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__B
timestamp 1669390400
transform -1 0 8400 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__I
timestamp 1669390400
transform 1 0 24304 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__I
timestamp 1669390400
transform 1 0 16912 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1626__I
timestamp 1669390400
transform -1 0 17472 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__A1
timestamp 1669390400
transform 1 0 16464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__A2
timestamp 1669390400
transform -1 0 15456 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__A3
timestamp 1669390400
transform 1 0 18816 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__A1
timestamp 1669390400
transform 1 0 19040 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__A2
timestamp 1669390400
transform 1 0 27664 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__A1
timestamp 1669390400
transform -1 0 35616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A2
timestamp 1669390400
transform -1 0 34048 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1633__A1
timestamp 1669390400
transform -1 0 38528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__I
timestamp 1669390400
transform 1 0 34944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1635__B
timestamp 1669390400
transform -1 0 34608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__A3
timestamp 1669390400
transform -1 0 35728 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1638__A1
timestamp 1669390400
transform 1 0 30688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1641__I
timestamp 1669390400
transform -1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__A1
timestamp 1669390400
transform 1 0 9856 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__A2
timestamp 1669390400
transform -1 0 8736 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__A1
timestamp 1669390400
transform 1 0 12096 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__A2
timestamp 1669390400
transform 1 0 8960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__A3
timestamp 1669390400
transform 1 0 14112 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A1
timestamp 1669390400
transform 1 0 10752 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__A2
timestamp 1669390400
transform -1 0 11424 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__A1
timestamp 1669390400
transform -1 0 7616 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__B
timestamp 1669390400
transform 1 0 11424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1647__I
timestamp 1669390400
transform -1 0 3696 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1648__A2
timestamp 1669390400
transform -1 0 15792 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__A1
timestamp 1669390400
transform 1 0 16464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__A1
timestamp 1669390400
transform 1 0 16016 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__B
timestamp 1669390400
transform 1 0 18032 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__A1
timestamp 1669390400
transform 1 0 4704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__A2
timestamp 1669390400
transform -1 0 5488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__A3
timestamp 1669390400
transform -1 0 6160 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__B
timestamp 1669390400
transform -1 0 1904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A1
timestamp 1669390400
transform 1 0 22512 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A3
timestamp 1669390400
transform 1 0 19040 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1655__A1
timestamp 1669390400
transform 1 0 26768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1655__A2
timestamp 1669390400
transform -1 0 21840 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A1
timestamp 1669390400
transform 1 0 29568 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A2
timestamp 1669390400
transform -1 0 30464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A3
timestamp 1669390400
transform -1 0 30016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__A2
timestamp 1669390400
transform -1 0 34608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__A1
timestamp 1669390400
transform 1 0 38080 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__A1
timestamp 1669390400
transform 1 0 12208 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__A2
timestamp 1669390400
transform 1 0 15120 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__A1
timestamp 1669390400
transform -1 0 2240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__A2
timestamp 1669390400
transform -1 0 5040 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__B
timestamp 1669390400
transform -1 0 2352 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A1
timestamp 1669390400
transform -1 0 2352 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A2
timestamp 1669390400
transform 1 0 4032 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A3
timestamp 1669390400
transform -1 0 1904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__A2
timestamp 1669390400
transform 1 0 3248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__B
timestamp 1669390400
transform -1 0 4368 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__A1
timestamp 1669390400
transform -1 0 10640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__A2
timestamp 1669390400
transform 1 0 4928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__B
timestamp 1669390400
transform -1 0 3920 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__A1
timestamp 1669390400
transform 1 0 24528 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__B1
timestamp 1669390400
transform -1 0 16016 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__B2
timestamp 1669390400
transform 1 0 21392 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__C
timestamp 1669390400
transform -1 0 15568 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__A2
timestamp 1669390400
transform 1 0 25648 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A1
timestamp 1669390400
transform -1 0 26432 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__A1
timestamp 1669390400
transform 1 0 25760 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__I
timestamp 1669390400
transform -1 0 27440 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__A2
timestamp 1669390400
transform -1 0 26432 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__A1
timestamp 1669390400
transform -1 0 17808 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__I0
timestamp 1669390400
transform 1 0 17920 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__I1
timestamp 1669390400
transform 1 0 15568 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__S
timestamp 1669390400
transform 1 0 16016 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1676__A2
timestamp 1669390400
transform 1 0 8624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A1
timestamp 1669390400
transform 1 0 10304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__A2
timestamp 1669390400
transform -1 0 6608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A1
timestamp 1669390400
transform 1 0 6496 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A2
timestamp 1669390400
transform 1 0 5376 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__B
timestamp 1669390400
transform -1 0 4032 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__A2
timestamp 1669390400
transform -1 0 5264 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__I
timestamp 1669390400
transform 1 0 38192 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__A1
timestamp 1669390400
transform -1 0 5264 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__B1
timestamp 1669390400
transform 1 0 12096 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__C
timestamp 1669390400
transform -1 0 2576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__A1
timestamp 1669390400
transform 1 0 8512 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__A2
timestamp 1669390400
transform 1 0 9744 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__A3
timestamp 1669390400
transform 1 0 10192 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A1
timestamp 1669390400
transform -1 0 15232 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A2
timestamp 1669390400
transform 1 0 11536 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__A1
timestamp 1669390400
transform -1 0 15232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__A2
timestamp 1669390400
transform 1 0 14896 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__A2
timestamp 1669390400
transform -1 0 28560 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__B
timestamp 1669390400
transform 1 0 30576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A2
timestamp 1669390400
transform -1 0 29008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__A2
timestamp 1669390400
transform -1 0 37744 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__A3
timestamp 1669390400
transform 1 0 36736 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__I
timestamp 1669390400
transform 1 0 40208 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__A1
timestamp 1669390400
transform -1 0 41216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__A2
timestamp 1669390400
transform 1 0 37520 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__I
timestamp 1669390400
transform 1 0 40432 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__A2
timestamp 1669390400
transform 1 0 39984 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A1
timestamp 1669390400
transform -1 0 4144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__A1
timestamp 1669390400
transform -1 0 3696 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__A2
timestamp 1669390400
transform -1 0 3248 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__A1
timestamp 1669390400
transform -1 0 2128 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__A4
timestamp 1669390400
transform 1 0 9072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__B1
timestamp 1669390400
transform 1 0 5824 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__B2
timestamp 1669390400
transform -1 0 4928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__A1
timestamp 1669390400
transform -1 0 7616 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__I
timestamp 1669390400
transform 1 0 17584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__A1
timestamp 1669390400
transform 1 0 13552 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__A2
timestamp 1669390400
transform 1 0 14896 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__A1
timestamp 1669390400
transform -1 0 5152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__A2
timestamp 1669390400
transform -1 0 9072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__A1
timestamp 1669390400
transform -1 0 3472 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__A2
timestamp 1669390400
transform -1 0 2800 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__A3
timestamp 1669390400
transform -1 0 4256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__A2
timestamp 1669390400
transform 1 0 12768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__A1
timestamp 1669390400
transform -1 0 5824 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1714__A2
timestamp 1669390400
transform -1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__I
timestamp 1669390400
transform 1 0 39536 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__I
timestamp 1669390400
transform -1 0 4816 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__A2
timestamp 1669390400
transform 1 0 38640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__B
timestamp 1669390400
transform -1 0 14224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__A1
timestamp 1669390400
transform 1 0 38640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__B
timestamp 1669390400
transform 1 0 32256 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__A3
timestamp 1669390400
transform 1 0 5376 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__A1
timestamp 1669390400
transform -1 0 6160 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__A2
timestamp 1669390400
transform -1 0 7056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__A1
timestamp 1669390400
transform 1 0 8512 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__A2
timestamp 1669390400
transform 1 0 8960 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__A1
timestamp 1669390400
transform -1 0 6272 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__A2
timestamp 1669390400
transform -1 0 5376 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__B2
timestamp 1669390400
transform -1 0 4256 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__A1
timestamp 1669390400
transform 1 0 20608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__B1
timestamp 1669390400
transform -1 0 17024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__B2
timestamp 1669390400
transform -1 0 15904 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__A3
timestamp 1669390400
transform 1 0 25200 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__A1
timestamp 1669390400
transform 1 0 27104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__B
timestamp 1669390400
transform 1 0 28896 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1729__A1
timestamp 1669390400
transform 1 0 26656 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__I
timestamp 1669390400
transform 1 0 38416 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__I
timestamp 1669390400
transform -1 0 2464 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1733__A1
timestamp 1669390400
transform 1 0 6048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__A1
timestamp 1669390400
transform 1 0 10752 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__B
timestamp 1669390400
transform 1 0 12096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__A1
timestamp 1669390400
transform -1 0 3248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__A2
timestamp 1669390400
transform 1 0 8960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__B1
timestamp 1669390400
transform -1 0 7504 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__B2
timestamp 1669390400
transform -1 0 3696 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__C
timestamp 1669390400
transform -1 0 2016 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__A2
timestamp 1669390400
transform 1 0 21168 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__A1
timestamp 1669390400
transform 1 0 29568 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__A2
timestamp 1669390400
transform 1 0 30016 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__A3
timestamp 1669390400
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__A1
timestamp 1669390400
transform 1 0 17584 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__A2
timestamp 1669390400
transform 1 0 12544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__A1
timestamp 1669390400
transform -1 0 2016 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__A2
timestamp 1669390400
transform -1 0 9072 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A1
timestamp 1669390400
transform -1 0 16464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A2
timestamp 1669390400
transform 1 0 25984 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__A2
timestamp 1669390400
transform 1 0 21392 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__A3
timestamp 1669390400
transform -1 0 18368 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__A1
timestamp 1669390400
transform 1 0 4256 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__A2
timestamp 1669390400
transform -1 0 7056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__A3
timestamp 1669390400
transform -1 0 4144 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__A2
timestamp 1669390400
transform 1 0 4144 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__B
timestamp 1669390400
transform -1 0 1904 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__A2
timestamp 1669390400
transform -1 0 2352 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__B1
timestamp 1669390400
transform -1 0 3920 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__B2
timestamp 1669390400
transform -1 0 2240 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__C
timestamp 1669390400
transform -1 0 8736 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__B
timestamp 1669390400
transform -1 0 10416 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__A1
timestamp 1669390400
transform 1 0 29456 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__A2
timestamp 1669390400
transform 1 0 30128 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__A1
timestamp 1669390400
transform 1 0 31024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__A1
timestamp 1669390400
transform 1 0 33488 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__A2
timestamp 1669390400
transform 1 0 31472 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1750__A2
timestamp 1669390400
transform 1 0 32816 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__B
timestamp 1669390400
transform 1 0 32816 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__A1
timestamp 1669390400
transform 1 0 36624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__I
timestamp 1669390400
transform -1 0 26320 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__A1
timestamp 1669390400
transform 1 0 28336 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__B
timestamp 1669390400
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__A1
timestamp 1669390400
transform 1 0 5824 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__A2
timestamp 1669390400
transform 1 0 6384 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__A2
timestamp 1669390400
transform 1 0 35616 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__B1
timestamp 1669390400
transform 1 0 34384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__B2
timestamp 1669390400
transform -1 0 31360 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__C
timestamp 1669390400
transform 1 0 33936 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__A2
timestamp 1669390400
transform -1 0 4704 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A2
timestamp 1669390400
transform -1 0 3360 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A3
timestamp 1669390400
transform 1 0 5712 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__A4
timestamp 1669390400
transform -1 0 5152 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A1
timestamp 1669390400
transform -1 0 2240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__A1
timestamp 1669390400
transform -1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__A2
timestamp 1669390400
transform -1 0 2016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__B
timestamp 1669390400
transform -1 0 11088 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1769__A1
timestamp 1669390400
transform -1 0 2016 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__A2
timestamp 1669390400
transform -1 0 2912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__A2
timestamp 1669390400
transform 1 0 25872 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__A4
timestamp 1669390400
transform 1 0 38528 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__B
timestamp 1669390400
transform 1 0 38640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__A2
timestamp 1669390400
transform 1 0 39984 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__I
timestamp 1669390400
transform -1 0 3360 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__A3
timestamp 1669390400
transform -1 0 25088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__A1
timestamp 1669390400
transform 1 0 25312 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__B
timestamp 1669390400
transform -1 0 26432 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__I
timestamp 1669390400
transform -1 0 4256 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1784__A2
timestamp 1669390400
transform -1 0 12656 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__A1
timestamp 1669390400
transform 1 0 8176 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__A2
timestamp 1669390400
transform -1 0 13776 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1786__I
timestamp 1669390400
transform 1 0 12992 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__A1
timestamp 1669390400
transform 1 0 14560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__A2
timestamp 1669390400
transform -1 0 10752 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A1
timestamp 1669390400
transform 1 0 15568 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A2
timestamp 1669390400
transform 1 0 16464 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__I
timestamp 1669390400
transform -1 0 22400 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__A1
timestamp 1669390400
transform -1 0 16016 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__A2
timestamp 1669390400
transform -1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__A1
timestamp 1669390400
transform 1 0 8064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__A2
timestamp 1669390400
transform -1 0 3024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__B
timestamp 1669390400
transform -1 0 2800 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__A1
timestamp 1669390400
transform 1 0 12880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__A2
timestamp 1669390400
transform -1 0 14560 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__A1
timestamp 1669390400
transform -1 0 16240 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__A2
timestamp 1669390400
transform 1 0 10640 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__B
timestamp 1669390400
transform -1 0 15344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__A1
timestamp 1669390400
transform 1 0 11984 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__B2
timestamp 1669390400
transform -1 0 7952 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__A2
timestamp 1669390400
transform 1 0 27552 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__B
timestamp 1669390400
transform 1 0 28672 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__A2
timestamp 1669390400
transform -1 0 25984 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__A1
timestamp 1669390400
transform -1 0 31248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__A2
timestamp 1669390400
transform 1 0 29904 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__A3
timestamp 1669390400
transform 1 0 30576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__I
timestamp 1669390400
transform -1 0 19040 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__I
timestamp 1669390400
transform -1 0 8064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__A1
timestamp 1669390400
transform -1 0 4928 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__A2
timestamp 1669390400
transform -1 0 10304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__B1
timestamp 1669390400
transform -1 0 10752 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__I0
timestamp 1669390400
transform 1 0 29792 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__S
timestamp 1669390400
transform 1 0 32928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__A1
timestamp 1669390400
transform -1 0 34048 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__A2
timestamp 1669390400
transform 1 0 33936 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__I
timestamp 1669390400
transform 1 0 37856 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__I
timestamp 1669390400
transform 1 0 41888 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__I
timestamp 1669390400
transform 1 0 40320 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__I
timestamp 1669390400
transform 1 0 40768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__A1
timestamp 1669390400
transform -1 0 37632 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__A2
timestamp 1669390400
transform 1 0 40432 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__B
timestamp 1669390400
transform -1 0 38080 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__A1
timestamp 1669390400
transform 1 0 31584 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__A2
timestamp 1669390400
transform 1 0 36512 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__B1
timestamp 1669390400
transform 1 0 37408 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__C
timestamp 1669390400
transform 1 0 33376 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__A1
timestamp 1669390400
transform -1 0 2576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__A2
timestamp 1669390400
transform -1 0 4704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__B2
timestamp 1669390400
transform -1 0 33264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__B
timestamp 1669390400
transform 1 0 33936 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__A3
timestamp 1669390400
transform 1 0 33600 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__A2
timestamp 1669390400
transform 1 0 25424 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__A3
timestamp 1669390400
transform -1 0 26096 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__A4
timestamp 1669390400
transform 1 0 26320 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__A1
timestamp 1669390400
transform 1 0 30688 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__A2
timestamp 1669390400
transform 1 0 31136 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__A1
timestamp 1669390400
transform 1 0 25872 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__B
timestamp 1669390400
transform -1 0 31808 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__A1
timestamp 1669390400
transform -1 0 5152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__A2
timestamp 1669390400
transform -1 0 8736 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__A2
timestamp 1669390400
transform 1 0 25984 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__A2
timestamp 1669390400
transform 1 0 34832 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__A1
timestamp 1669390400
transform 1 0 39984 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__A1
timestamp 1669390400
transform 1 0 30688 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__A2
timestamp 1669390400
transform 1 0 32032 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__B2
timestamp 1669390400
transform 1 0 32480 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__A1
timestamp 1669390400
transform -1 0 3808 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1827__B2
timestamp 1669390400
transform -1 0 2352 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1828__A2
timestamp 1669390400
transform 1 0 29456 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__A1
timestamp 1669390400
transform 1 0 40432 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1829__A4
timestamp 1669390400
transform 1 0 36736 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__I
timestamp 1669390400
transform 1 0 38976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__A1
timestamp 1669390400
transform -1 0 37296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__B
timestamp 1669390400
transform 1 0 39872 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1832__A1
timestamp 1669390400
transform 1 0 41776 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__B
timestamp 1669390400
transform -1 0 43344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1835__A1
timestamp 1669390400
transform -1 0 41104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1835__A4
timestamp 1669390400
transform 1 0 40320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1836__A1
timestamp 1669390400
transform 1 0 41440 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__A1
timestamp 1669390400
transform 1 0 40768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1845__I
timestamp 1669390400
transform -1 0 3360 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1846__A1
timestamp 1669390400
transform 1 0 42336 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__A2
timestamp 1669390400
transform 1 0 31920 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__B2
timestamp 1669390400
transform 1 0 35280 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1850__A1
timestamp 1669390400
transform 1 0 15792 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1850__A2
timestamp 1669390400
transform 1 0 18816 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1850__B
timestamp 1669390400
transform 1 0 18928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1851__A1
timestamp 1669390400
transform 1 0 23856 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1851__A3
timestamp 1669390400
transform 1 0 22512 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__A1
timestamp 1669390400
transform 1 0 9744 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__A2
timestamp 1669390400
transform -1 0 11984 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__B
timestamp 1669390400
transform 1 0 5600 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__I
timestamp 1669390400
transform -1 0 22288 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__A1
timestamp 1669390400
transform 1 0 23632 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__A2
timestamp 1669390400
transform 1 0 30240 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__I0
timestamp 1669390400
transform 1 0 33488 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1857__A1
timestamp 1669390400
transform 1 0 32928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1858__A1
timestamp 1669390400
transform 1 0 37632 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__I
timestamp 1669390400
transform -1 0 6720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__A1
timestamp 1669390400
transform 1 0 25424 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__A2
timestamp 1669390400
transform -1 0 25200 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__C
timestamp 1669390400
transform -1 0 19488 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__A2
timestamp 1669390400
transform 1 0 17696 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1863__A1
timestamp 1669390400
transform -1 0 5152 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1863__A2
timestamp 1669390400
transform -1 0 4144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1863__B
timestamp 1669390400
transform -1 0 2688 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1863__C
timestamp 1669390400
transform -1 0 2016 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__A1
timestamp 1669390400
transform 1 0 20832 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__B1
timestamp 1669390400
transform -1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1864__B2
timestamp 1669390400
transform -1 0 18368 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1865__A1
timestamp 1669390400
transform 1 0 31136 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1865__A2
timestamp 1669390400
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1865__B
timestamp 1669390400
transform 1 0 30688 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A1
timestamp 1669390400
transform 1 0 31472 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1867__I
timestamp 1669390400
transform 1 0 24080 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__I
timestamp 1669390400
transform -1 0 22064 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1869__A1
timestamp 1669390400
transform 1 0 19712 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1869__A2
timestamp 1669390400
transform 1 0 19824 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A1
timestamp 1669390400
transform 1 0 22288 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__I
timestamp 1669390400
transform 1 0 21280 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1873__A1
timestamp 1669390400
transform 1 0 25536 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1873__A2
timestamp 1669390400
transform 1 0 17584 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1873__C
timestamp 1669390400
transform 1 0 15568 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A1
timestamp 1669390400
transform -1 0 15344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A2
timestamp 1669390400
transform -1 0 14448 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__B1
timestamp 1669390400
transform -1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__C
timestamp 1669390400
transform -1 0 12208 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1875__A3
timestamp 1669390400
transform 1 0 21616 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A3
timestamp 1669390400
transform -1 0 12656 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1878__A1
timestamp 1669390400
transform 1 0 25648 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1878__A3
timestamp 1669390400
transform -1 0 28000 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1880__A1
timestamp 1669390400
transform 1 0 27664 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__A1
timestamp 1669390400
transform 1 0 29008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__A2
timestamp 1669390400
transform 1 0 40768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__A3
timestamp 1669390400
transform 1 0 38080 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__A2
timestamp 1669390400
transform 1 0 30688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__A2
timestamp 1669390400
transform 1 0 39088 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__A3
timestamp 1669390400
transform -1 0 27440 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__A2
timestamp 1669390400
transform -1 0 15568 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1893__A1
timestamp 1669390400
transform -1 0 11760 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__A1
timestamp 1669390400
transform 1 0 12432 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__A2
timestamp 1669390400
transform 1 0 5600 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__B
timestamp 1669390400
transform 1 0 12880 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1894__C
timestamp 1669390400
transform 1 0 5488 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__A1
timestamp 1669390400
transform 1 0 15456 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1896__A1
timestamp 1669390400
transform -1 0 15120 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1896__A2
timestamp 1669390400
transform 1 0 14112 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1896__A3
timestamp 1669390400
transform -1 0 20272 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__A1
timestamp 1669390400
transform -1 0 14672 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__B
timestamp 1669390400
transform -1 0 11200 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__B
timestamp 1669390400
transform -1 0 33712 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__A3
timestamp 1669390400
transform 1 0 34832 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__A1
timestamp 1669390400
transform 1 0 28224 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__A2
timestamp 1669390400
transform 1 0 28560 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__A3
timestamp 1669390400
transform 1 0 26096 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__B
timestamp 1669390400
transform 1 0 30688 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1903__A2
timestamp 1669390400
transform 1 0 8064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1904__A1
timestamp 1669390400
transform 1 0 12880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1904__A2
timestamp 1669390400
transform -1 0 2464 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1905__A2
timestamp 1669390400
transform -1 0 21952 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1905__A3
timestamp 1669390400
transform -1 0 21168 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1905__B1
timestamp 1669390400
transform 1 0 21280 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__I1
timestamp 1669390400
transform 1 0 31472 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1907__A4
timestamp 1669390400
transform 1 0 38976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1908__B
timestamp 1669390400
transform 1 0 36512 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__I
timestamp 1669390400
transform 1 0 32032 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1911__A1
timestamp 1669390400
transform -1 0 13776 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1911__A3
timestamp 1669390400
transform -1 0 14224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__A1
timestamp 1669390400
transform 1 0 29792 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__A2
timestamp 1669390400
transform 1 0 29344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__B
timestamp 1669390400
transform -1 0 5152 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__B1
timestamp 1669390400
transform 1 0 23072 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__A1
timestamp 1669390400
transform 1 0 22512 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__A3
timestamp 1669390400
transform 1 0 22064 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__A1
timestamp 1669390400
transform -1 0 25200 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__A3
timestamp 1669390400
transform 1 0 25424 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__A1
timestamp 1669390400
transform -1 0 36960 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__A4
timestamp 1669390400
transform 1 0 38864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__B1
timestamp 1669390400
transform 1 0 36288 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__B2
timestamp 1669390400
transform 1 0 37296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__A1
timestamp 1669390400
transform 1 0 38304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__B
timestamp 1669390400
transform 1 0 39200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1925__A3
timestamp 1669390400
transform 1 0 38976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A2
timestamp 1669390400
transform 1 0 39648 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1933__I
timestamp 1669390400
transform -1 0 42896 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1934__A1
timestamp 1669390400
transform -1 0 37632 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1936__A3
timestamp 1669390400
transform 1 0 35840 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1938__A1
timestamp 1669390400
transform 1 0 34384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1938__A2
timestamp 1669390400
transform 1 0 36960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1939__A1
timestamp 1669390400
transform 1 0 38752 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1939__A2
timestamp 1669390400
transform 1 0 40432 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1941__A1
timestamp 1669390400
transform 1 0 40880 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1941__A2
timestamp 1669390400
transform 1 0 43568 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1942__A1
timestamp 1669390400
transform 1 0 39984 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1942__A2
timestamp 1669390400
transform 1 0 39536 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1943__A1
timestamp 1669390400
transform 1 0 34272 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1943__A2
timestamp 1669390400
transform 1 0 35504 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1944__A1
timestamp 1669390400
transform 1 0 39088 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1944__B2
timestamp 1669390400
transform 1 0 39536 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1945__I0
timestamp 1669390400
transform 1 0 31136 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1945__S
timestamp 1669390400
transform -1 0 31136 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__A1
timestamp 1669390400
transform 1 0 35056 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__A1
timestamp 1669390400
transform 1 0 37296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__B
timestamp 1669390400
transform 1 0 34720 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__C
timestamp 1669390400
transform 1 0 37408 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__A1
timestamp 1669390400
transform -1 0 3808 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__B1
timestamp 1669390400
transform 1 0 34608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__B2
timestamp 1669390400
transform -1 0 31360 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__C
timestamp 1669390400
transform -1 0 2128 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1951__A1
timestamp 1669390400
transform 1 0 20272 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__A1
timestamp 1669390400
transform 1 0 25536 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__A2
timestamp 1669390400
transform 1 0 24416 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1953__A2
timestamp 1669390400
transform 1 0 24752 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1957__I
timestamp 1669390400
transform -1 0 25424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__A2
timestamp 1669390400
transform -1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__A2
timestamp 1669390400
transform -1 0 8176 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__A3
timestamp 1669390400
transform -1 0 6608 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__B1
timestamp 1669390400
transform -1 0 5264 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__B2
timestamp 1669390400
transform -1 0 4816 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__A1
timestamp 1669390400
transform 1 0 28448 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1962__B
timestamp 1669390400
transform 1 0 28224 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__A3
timestamp 1669390400
transform -1 0 37968 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__I
timestamp 1669390400
transform 1 0 3136 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__A1
timestamp 1669390400
transform 1 0 20608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__A2
timestamp 1669390400
transform 1 0 20720 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__B
timestamp 1669390400
transform 1 0 24752 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1976__A1
timestamp 1669390400
transform 1 0 25424 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1977__A1
timestamp 1669390400
transform 1 0 30240 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1977__A2
timestamp 1669390400
transform 1 0 26320 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__A1
timestamp 1669390400
transform 1 0 38304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__A2
timestamp 1669390400
transform 1 0 40320 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1979__A2
timestamp 1669390400
transform -1 0 32256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__A2
timestamp 1669390400
transform -1 0 5936 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__B1
timestamp 1669390400
transform -1 0 6832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__B2
timestamp 1669390400
transform 1 0 30576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__B2
timestamp 1669390400
transform 1 0 26208 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1982__A2
timestamp 1669390400
transform 1 0 32592 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__A1
timestamp 1669390400
transform 1 0 34384 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__A2
timestamp 1669390400
transform 1 0 31248 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__A1
timestamp 1669390400
transform 1 0 35168 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A1
timestamp 1669390400
transform -1 0 18032 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A2
timestamp 1669390400
transform -1 0 17584 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1987__A2
timestamp 1669390400
transform -1 0 16912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__A1
timestamp 1669390400
transform 1 0 26992 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1989__A1
timestamp 1669390400
transform -1 0 25872 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1990__A1
timestamp 1669390400
transform 1 0 28896 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1990__A2
timestamp 1669390400
transform 1 0 29344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1991__A2
timestamp 1669390400
transform 1 0 40768 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__I
timestamp 1669390400
transform -1 0 26656 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1993__A2
timestamp 1669390400
transform 1 0 24528 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__A1
timestamp 1669390400
transform 1 0 26656 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__A2
timestamp 1669390400
transform 1 0 26096 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1996__A2
timestamp 1669390400
transform 1 0 25760 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__C
timestamp 1669390400
transform -1 0 30016 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__A2
timestamp 1669390400
transform 1 0 41552 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__A2
timestamp 1669390400
transform -1 0 39312 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2009__I
timestamp 1669390400
transform -1 0 48048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__A2
timestamp 1669390400
transform 1 0 42448 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__A2
timestamp 1669390400
transform 1 0 41664 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__I
timestamp 1669390400
transform 1 0 21280 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__A1
timestamp 1669390400
transform -1 0 17472 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__A2
timestamp 1669390400
transform 1 0 17472 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__B
timestamp 1669390400
transform 1 0 18592 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__A2
timestamp 1669390400
transform -1 0 6384 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2016__A2
timestamp 1669390400
transform 1 0 22736 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2017__A1
timestamp 1669390400
transform 1 0 24976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__B
timestamp 1669390400
transform -1 0 31920 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__A1
timestamp 1669390400
transform 1 0 32592 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__A2
timestamp 1669390400
transform 1 0 33488 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__C
timestamp 1669390400
transform 1 0 35056 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__A1
timestamp 1669390400
transform -1 0 20272 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__A2
timestamp 1669390400
transform 1 0 24528 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__A3
timestamp 1669390400
transform 1 0 20496 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__A2
timestamp 1669390400
transform -1 0 24528 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__A1
timestamp 1669390400
transform 1 0 29344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__I
timestamp 1669390400
transform 1 0 31584 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2028__A1
timestamp 1669390400
transform 1 0 27104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2028__A2
timestamp 1669390400
transform 1 0 26544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2030__A1
timestamp 1669390400
transform -1 0 6608 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2030__A2
timestamp 1669390400
transform -1 0 5712 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2031__A1
timestamp 1669390400
transform 1 0 8848 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2031__B
timestamp 1669390400
transform -1 0 8624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2032__A1
timestamp 1669390400
transform -1 0 20832 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__A1
timestamp 1669390400
transform -1 0 32704 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__A2
timestamp 1669390400
transform 1 0 44016 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__A1
timestamp 1669390400
transform -1 0 34608 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__A1
timestamp 1669390400
transform -1 0 35280 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2044__A1
timestamp 1669390400
transform 1 0 4480 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2044__B
timestamp 1669390400
transform -1 0 9856 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__A1
timestamp 1669390400
transform 1 0 23520 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__B2
timestamp 1669390400
transform 1 0 21728 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2046__A2
timestamp 1669390400
transform 1 0 36736 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__A1
timestamp 1669390400
transform 1 0 38192 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2048__A1
timestamp 1669390400
transform -1 0 26208 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__A1
timestamp 1669390400
transform 1 0 28448 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__A2
timestamp 1669390400
transform 1 0 28896 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__B
timestamp 1669390400
transform 1 0 25536 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__A2
timestamp 1669390400
transform 1 0 36736 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__A1
timestamp 1669390400
transform 1 0 20832 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2052__A2
timestamp 1669390400
transform -1 0 22176 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2055__A1
timestamp 1669390400
transform 1 0 30800 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2058__A1
timestamp 1669390400
transform -1 0 32256 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2060__A2
timestamp 1669390400
transform -1 0 42000 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2061__A2
timestamp 1669390400
transform 1 0 43008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__A2
timestamp 1669390400
transform -1 0 44240 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2066__A2
timestamp 1669390400
transform 1 0 38640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2068__A1
timestamp 1669390400
transform 1 0 24864 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2069__A1
timestamp 1669390400
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2070__A1
timestamp 1669390400
transform 1 0 31248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2072__A1
timestamp 1669390400
transform 1 0 33376 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2073__A1
timestamp 1669390400
transform 1 0 33488 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2077__A2
timestamp 1669390400
transform 1 0 44128 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__B
timestamp 1669390400
transform 1 0 35056 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2087__B2
timestamp 1669390400
transform 1 0 40768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2088__A1
timestamp 1669390400
transform 1 0 41776 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2089__I
timestamp 1669390400
transform 1 0 47824 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__A1
timestamp 1669390400
transform 1 0 46592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__A2
timestamp 1669390400
transform 1 0 46144 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2092__I
timestamp 1669390400
transform 1 0 49056 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2096__A2
timestamp 1669390400
transform -1 0 50512 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2097__A1
timestamp 1669390400
transform 1 0 54208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2097__A2
timestamp 1669390400
transform 1 0 52304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2098__I
timestamp 1669390400
transform 1 0 49840 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2101__I
timestamp 1669390400
transform 1 0 44688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2102__I
timestamp 1669390400
transform 1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2103__A1
timestamp 1669390400
transform 1 0 45360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2103__B
timestamp 1669390400
transform -1 0 46592 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2106__I
timestamp 1669390400
transform 1 0 46144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2107__I
timestamp 1669390400
transform 1 0 57344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2108__A1
timestamp 1669390400
transform -1 0 56000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__I
timestamp 1669390400
transform 1 0 58016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2111__A2
timestamp 1669390400
transform -1 0 47264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2111__B
timestamp 1669390400
transform 1 0 46592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2113__I
timestamp 1669390400
transform 1 0 57792 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2114__A1
timestamp 1669390400
transform 1 0 49392 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2114__A2
timestamp 1669390400
transform 1 0 49840 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2114__C
timestamp 1669390400
transform 1 0 49504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2115__A2
timestamp 1669390400
transform 1 0 57792 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2116__A1
timestamp 1669390400
transform 1 0 56000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2122__A1
timestamp 1669390400
transform 1 0 54880 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2123__A1
timestamp 1669390400
transform 1 0 51744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2123__A2
timestamp 1669390400
transform 1 0 56112 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__A1
timestamp 1669390400
transform 1 0 55552 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__B
timestamp 1669390400
transform 1 0 56000 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2128__A2
timestamp 1669390400
transform -1 0 56896 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2128__B
timestamp 1669390400
transform -1 0 56448 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__A1
timestamp 1669390400
transform -1 0 50960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__A2
timestamp 1669390400
transform -1 0 51408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2130__I
timestamp 1669390400
transform 1 0 41888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2132__I
timestamp 1669390400
transform -1 0 46256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2133__A2
timestamp 1669390400
transform 1 0 57232 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2135__I
timestamp 1669390400
transform 1 0 54432 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2136__I
timestamp 1669390400
transform 1 0 43680 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__A1
timestamp 1669390400
transform 1 0 47376 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2138__A2
timestamp 1669390400
transform -1 0 44576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2139__A1
timestamp 1669390400
transform -1 0 38864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2139__A2
timestamp 1669390400
transform -1 0 46592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2139__B1
timestamp 1669390400
transform -1 0 45136 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2141__I
timestamp 1669390400
transform -1 0 43904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__A2
timestamp 1669390400
transform 1 0 45920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2143__I
timestamp 1669390400
transform 1 0 52416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2144__I
timestamp 1669390400
transform -1 0 55776 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2145__A1
timestamp 1669390400
transform -1 0 53088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2145__A2
timestamp 1669390400
transform -1 0 52640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2147__A1
timestamp 1669390400
transform -1 0 55328 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2147__B
timestamp 1669390400
transform -1 0 55776 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2148__I
timestamp 1669390400
transform -1 0 57456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__A1
timestamp 1669390400
transform -1 0 56000 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2150__A3
timestamp 1669390400
transform -1 0 54992 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2151__A2
timestamp 1669390400
transform -1 0 54880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2151__B
timestamp 1669390400
transform -1 0 54544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2151__C
timestamp 1669390400
transform -1 0 55328 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2154__B
timestamp 1669390400
transform -1 0 54432 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2155__I
timestamp 1669390400
transform 1 0 55552 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2156__I
timestamp 1669390400
transform 1 0 56000 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2157__A1
timestamp 1669390400
transform 1 0 57792 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2157__A2
timestamp 1669390400
transform 1 0 55776 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2157__B
timestamp 1669390400
transform 1 0 56448 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2159__A1
timestamp 1669390400
transform 1 0 57344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2159__B
timestamp 1669390400
transform 1 0 57680 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2161__A1
timestamp 1669390400
transform 1 0 53760 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2161__A2
timestamp 1669390400
transform 1 0 56112 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2161__B
timestamp 1669390400
transform 1 0 57792 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2163__A1
timestamp 1669390400
transform -1 0 53760 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2163__A2
timestamp 1669390400
transform -1 0 48944 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2164__A1
timestamp 1669390400
transform 1 0 58016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__A1
timestamp 1669390400
transform 1 0 56448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__A2
timestamp 1669390400
transform 1 0 56000 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__B1
timestamp 1669390400
transform 1 0 54096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__B2
timestamp 1669390400
transform 1 0 57344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__C
timestamp 1669390400
transform -1 0 56448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2170__I
timestamp 1669390400
transform -1 0 52976 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__A1
timestamp 1669390400
transform -1 0 55664 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__A2
timestamp 1669390400
transform 1 0 55888 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__B
timestamp 1669390400
transform 1 0 55104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__C
timestamp 1669390400
transform 1 0 57680 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2174__I
timestamp 1669390400
transform 1 0 52976 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2175__A1
timestamp 1669390400
transform 1 0 53200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2175__A2
timestamp 1669390400
transform 1 0 54096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2176__A1
timestamp 1669390400
transform 1 0 53312 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2176__A2
timestamp 1669390400
transform 1 0 56560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2176__B
timestamp 1669390400
transform 1 0 56336 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2177__I
timestamp 1669390400
transform -1 0 50288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2178__I
timestamp 1669390400
transform 1 0 57568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2179__A1
timestamp 1669390400
transform 1 0 53648 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2179__B2
timestamp 1669390400
transform 1 0 55552 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2179__C
timestamp 1669390400
transform 1 0 53760 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__A1
timestamp 1669390400
transform 1 0 48720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__A2
timestamp 1669390400
transform 1 0 49168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__B
timestamp 1669390400
transform 1 0 48720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2182__A1
timestamp 1669390400
transform -1 0 53984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2182__A2
timestamp 1669390400
transform 1 0 57904 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2182__C
timestamp 1669390400
transform 1 0 51072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2183__I
timestamp 1669390400
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2184__A1
timestamp 1669390400
transform -1 0 47600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2186__A1
timestamp 1669390400
transform -1 0 54432 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2189__A1
timestamp 1669390400
transform 1 0 55552 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2190__I
timestamp 1669390400
transform 1 0 47152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__I
timestamp 1669390400
transform 1 0 48160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__A1
timestamp 1669390400
transform -1 0 48272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__A2
timestamp 1669390400
transform 1 0 48496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__B
timestamp 1669390400
transform -1 0 48720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2194__A1
timestamp 1669390400
transform -1 0 47824 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2194__A2
timestamp 1669390400
transform 1 0 48048 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2196__A2
timestamp 1669390400
transform 1 0 48496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2196__B
timestamp 1669390400
transform 1 0 48944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2197__I
timestamp 1669390400
transform 1 0 48272 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2198__B
timestamp 1669390400
transform -1 0 48160 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2203__A1
timestamp 1669390400
transform -1 0 45808 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2203__A2
timestamp 1669390400
transform 1 0 47488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2205__A1
timestamp 1669390400
transform 1 0 49280 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2205__A2
timestamp 1669390400
transform 1 0 51520 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2205__C
timestamp 1669390400
transform 1 0 51968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2207__A2
timestamp 1669390400
transform 1 0 57904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2208__A1
timestamp 1669390400
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2208__A2
timestamp 1669390400
transform -1 0 46032 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2208__B
timestamp 1669390400
transform 1 0 48832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2208__C
timestamp 1669390400
transform 1 0 49056 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2209__A1
timestamp 1669390400
transform 1 0 45360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2211__A1
timestamp 1669390400
transform -1 0 43680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2213__A1
timestamp 1669390400
transform 1 0 45360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2217__I
timestamp 1669390400
transform -1 0 49616 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__A1
timestamp 1669390400
transform -1 0 49168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__A2
timestamp 1669390400
transform -1 0 48720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2219__A1
timestamp 1669390400
transform -1 0 54656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2219__A2
timestamp 1669390400
transform 1 0 54656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2221__A1
timestamp 1669390400
transform -1 0 50960 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2221__A2
timestamp 1669390400
transform 1 0 50176 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2222__A1
timestamp 1669390400
transform 1 0 52640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2222__A2
timestamp 1669390400
transform 1 0 51744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2222__A3
timestamp 1669390400
transform -1 0 53984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2223__A1
timestamp 1669390400
transform -1 0 53312 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2223__A2
timestamp 1669390400
transform -1 0 56336 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2224__A2
timestamp 1669390400
transform -1 0 54880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2224__A3
timestamp 1669390400
transform -1 0 53536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2225__A1
timestamp 1669390400
transform 1 0 55216 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2226__A1
timestamp 1669390400
transform 1 0 53312 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2226__B1
timestamp 1669390400
transform 1 0 53760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2226__B2
timestamp 1669390400
transform 1 0 52416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2227__A3
timestamp 1669390400
transform -1 0 47824 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2229__A1
timestamp 1669390400
transform -1 0 46480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2229__B
timestamp 1669390400
transform 1 0 47824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2230__A1
timestamp 1669390400
transform -1 0 47376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2231__A1
timestamp 1669390400
transform 1 0 57344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2231__A2
timestamp 1669390400
transform -1 0 54432 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2232__A1
timestamp 1669390400
transform 1 0 54208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2232__A2
timestamp 1669390400
transform 1 0 53760 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2234__A1
timestamp 1669390400
transform 1 0 52080 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2234__B
timestamp 1669390400
transform 1 0 52528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__A1
timestamp 1669390400
transform 1 0 56336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__A2
timestamp 1669390400
transform 1 0 56784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__A3
timestamp 1669390400
transform -1 0 51744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__B
timestamp 1669390400
transform -1 0 51072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2236__A1
timestamp 1669390400
transform 1 0 57344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2236__A2
timestamp 1669390400
transform 1 0 53312 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2237__A1
timestamp 1669390400
transform -1 0 51968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2237__A2
timestamp 1669390400
transform -1 0 51520 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2237__A3
timestamp 1669390400
transform 1 0 53760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2238__A1
timestamp 1669390400
transform 1 0 51968 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2240__A1
timestamp 1669390400
transform 1 0 50400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2247__I
timestamp 1669390400
transform 1 0 29456 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2249__A1
timestamp 1669390400
transform 1 0 25088 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2251__I
timestamp 1669390400
transform 1 0 46704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__A1
timestamp 1669390400
transform -1 0 40880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__A2
timestamp 1669390400
transform -1 0 40432 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2255__B
timestamp 1669390400
transform -1 0 49392 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2256__I
timestamp 1669390400
transform 1 0 43680 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2257__A1
timestamp 1669390400
transform 1 0 46592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2257__B
timestamp 1669390400
transform 1 0 43344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2257__C
timestamp 1669390400
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2258__A2
timestamp 1669390400
transform 1 0 42112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2260__A1
timestamp 1669390400
transform -1 0 44800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2260__A2
timestamp 1669390400
transform 1 0 44128 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2261__A2
timestamp 1669390400
transform 1 0 48160 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2262__A1
timestamp 1669390400
transform 1 0 51408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2262__A2
timestamp 1669390400
transform 1 0 51744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2263__A2
timestamp 1669390400
transform 1 0 47712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2263__B
timestamp 1669390400
transform -1 0 48272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2264__A1
timestamp 1669390400
transform 1 0 43568 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2264__A3
timestamp 1669390400
transform -1 0 44240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2265__A1
timestamp 1669390400
transform 1 0 48048 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2265__A2
timestamp 1669390400
transform 1 0 47040 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2265__B
timestamp 1669390400
transform 1 0 45920 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2266__I
timestamp 1669390400
transform 1 0 52640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2267__A1
timestamp 1669390400
transform 1 0 45360 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2267__A2
timestamp 1669390400
transform -1 0 43680 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2267__B
timestamp 1669390400
transform 1 0 45024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2268__A1
timestamp 1669390400
transform 1 0 45472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2269__A1
timestamp 1669390400
transform 1 0 46032 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2269__A2
timestamp 1669390400
transform 1 0 46480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2270__A1
timestamp 1669390400
transform 1 0 46480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2271__A1
timestamp 1669390400
transform 1 0 33152 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2271__A2
timestamp 1669390400
transform -1 0 30688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2272__A1
timestamp 1669390400
transform -1 0 29120 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2272__A2
timestamp 1669390400
transform 1 0 32144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2275__A1
timestamp 1669390400
transform -1 0 57120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2275__A2
timestamp 1669390400
transform 1 0 56896 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2275__C
timestamp 1669390400
transform -1 0 57568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2276__A1
timestamp 1669390400
transform -1 0 55888 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2277__A1
timestamp 1669390400
transform 1 0 51856 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2278__A1
timestamp 1669390400
transform 1 0 52304 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2278__A3
timestamp 1669390400
transform -1 0 52416 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2279__A1
timestamp 1669390400
transform 1 0 54208 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2279__A2
timestamp 1669390400
transform -1 0 54880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2280__A1
timestamp 1669390400
transform 1 0 58016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2280__B
timestamp 1669390400
transform 1 0 58016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2281__A1
timestamp 1669390400
transform -1 0 57904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2282__A1
timestamp 1669390400
transform 1 0 54544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2282__A2
timestamp 1669390400
transform -1 0 55216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2282__B1
timestamp 1669390400
transform -1 0 54432 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2282__B2
timestamp 1669390400
transform 1 0 53312 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2282__C
timestamp 1669390400
transform -1 0 56672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2283__A1
timestamp 1669390400
transform 1 0 54656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2284__A2
timestamp 1669390400
transform 1 0 46704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2285__A1
timestamp 1669390400
transform -1 0 46928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2286__B
timestamp 1669390400
transform 1 0 49616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2287__I
timestamp 1669390400
transform -1 0 56896 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2288__A1
timestamp 1669390400
transform 1 0 57344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2288__B
timestamp 1669390400
transform 1 0 57232 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2289__A2
timestamp 1669390400
transform 1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A1
timestamp 1669390400
transform -1 0 51744 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A2
timestamp 1669390400
transform 1 0 54656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__B
timestamp 1669390400
transform 1 0 52640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__C
timestamp 1669390400
transform 1 0 52192 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2291__A1
timestamp 1669390400
transform 1 0 55104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2292__A1
timestamp 1669390400
transform 1 0 57344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2292__A2
timestamp 1669390400
transform 1 0 56784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2292__B1
timestamp 1669390400
transform 1 0 54656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2292__B2
timestamp 1669390400
transform 1 0 54544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2293__B
timestamp 1669390400
transform 1 0 55104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2294__I
timestamp 1669390400
transform 1 0 42448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2295__A2
timestamp 1669390400
transform 1 0 42560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2296__A1
timestamp 1669390400
transform 1 0 50176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2296__A2
timestamp 1669390400
transform 1 0 50624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2296__A3
timestamp 1669390400
transform 1 0 51968 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2297__A1
timestamp 1669390400
transform -1 0 51744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2299__A1
timestamp 1669390400
transform 1 0 38304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2299__A2
timestamp 1669390400
transform -1 0 37184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2299__A3
timestamp 1669390400
transform -1 0 37632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2300__I
timestamp 1669390400
transform -1 0 34720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2301__A2
timestamp 1669390400
transform 1 0 36624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2301__B
timestamp 1669390400
transform 1 0 37408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2303__A1
timestamp 1669390400
transform -1 0 33824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2304__A1
timestamp 1669390400
transform -1 0 33264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2308__A1
timestamp 1669390400
transform 1 0 30912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2309__A1
timestamp 1669390400
transform 1 0 33824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2310__A1
timestamp 1669390400
transform 1 0 33488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2311__A2
timestamp 1669390400
transform -1 0 36064 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2311__A3
timestamp 1669390400
transform 1 0 37408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2313__I
timestamp 1669390400
transform 1 0 32816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2314__A2
timestamp 1669390400
transform 1 0 42000 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__A2
timestamp 1669390400
transform 1 0 41552 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__B
timestamp 1669390400
transform 1 0 40096 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__C
timestamp 1669390400
transform 1 0 40544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2316__A1
timestamp 1669390400
transform 1 0 40320 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2316__A2
timestamp 1669390400
transform 1 0 40768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2317__I
timestamp 1669390400
transform 1 0 47600 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2318__A1
timestamp 1669390400
transform 1 0 44464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2319__A1
timestamp 1669390400
transform 1 0 43232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2319__B
timestamp 1669390400
transform -1 0 43904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__A1
timestamp 1669390400
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__A2
timestamp 1669390400
transform 1 0 39648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__A3
timestamp 1669390400
transform -1 0 40320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2322__A1
timestamp 1669390400
transform 1 0 38752 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2322__A2
timestamp 1669390400
transform -1 0 39424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2325__A2
timestamp 1669390400
transform 1 0 33600 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2325__C
timestamp 1669390400
transform -1 0 34272 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2326__I
timestamp 1669390400
transform 1 0 42336 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2327__A1
timestamp 1669390400
transform -1 0 41888 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2327__A2
timestamp 1669390400
transform 1 0 43232 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2328__A2
timestamp 1669390400
transform -1 0 43568 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2328__B
timestamp 1669390400
transform 1 0 47936 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__A1
timestamp 1669390400
transform 1 0 44688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__B
timestamp 1669390400
transform 1 0 42784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2330__A1
timestamp 1669390400
transform 1 0 45360 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2330__A2
timestamp 1669390400
transform -1 0 43008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2330__B
timestamp 1669390400
transform 1 0 46032 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2331__I
timestamp 1669390400
transform 1 0 45360 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2332__A1
timestamp 1669390400
transform -1 0 44464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2335__A1
timestamp 1669390400
transform 1 0 33936 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2336__A2
timestamp 1669390400
transform 1 0 33488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2337__A1
timestamp 1669390400
transform -1 0 26880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2338__I
timestamp 1669390400
transform -1 0 24752 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2340__A1
timestamp 1669390400
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2342__A1
timestamp 1669390400
transform 1 0 48720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2342__A2
timestamp 1669390400
transform 1 0 49168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2342__A3
timestamp 1669390400
transform 1 0 48272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2344__I
timestamp 1669390400
transform 1 0 31808 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2345__A1
timestamp 1669390400
transform -1 0 50848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2345__A2
timestamp 1669390400
transform 1 0 52080 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2346__A1
timestamp 1669390400
transform -1 0 49168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2347__A2
timestamp 1669390400
transform 1 0 47264 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2347__B
timestamp 1669390400
transform 1 0 46816 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2349__A2
timestamp 1669390400
transform 1 0 50288 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2350__I
timestamp 1669390400
transform 1 0 48160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2351__A1
timestamp 1669390400
transform 1 0 50400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2351__A2
timestamp 1669390400
transform 1 0 51296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2351__B1
timestamp 1669390400
transform 1 0 48944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2351__B2
timestamp 1669390400
transform 1 0 48720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2351__C
timestamp 1669390400
transform 1 0 50848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2352__A1
timestamp 1669390400
transform 1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2352__B
timestamp 1669390400
transform 1 0 47488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__A1
timestamp 1669390400
transform 1 0 49952 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__A2
timestamp 1669390400
transform -1 0 48832 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__B1
timestamp 1669390400
transform 1 0 52752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__B2
timestamp 1669390400
transform 1 0 50960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__C
timestamp 1669390400
transform 1 0 53200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2355__A1
timestamp 1669390400
transform 1 0 47600 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2356__I
timestamp 1669390400
transform 1 0 42112 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2358__A2
timestamp 1669390400
transform -1 0 42784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2359__A1
timestamp 1669390400
transform 1 0 43008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2360__I
timestamp 1669390400
transform 1 0 36736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2361__I
timestamp 1669390400
transform 1 0 48384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2362__A1
timestamp 1669390400
transform 1 0 52416 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2362__A2
timestamp 1669390400
transform 1 0 54208 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2363__A1
timestamp 1669390400
transform 1 0 56560 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2363__A2
timestamp 1669390400
transform -1 0 52640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2363__B2
timestamp 1669390400
transform -1 0 52192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2364__B
timestamp 1669390400
transform -1 0 47712 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2365__A1
timestamp 1669390400
transform 1 0 49840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2365__A2
timestamp 1669390400
transform 1 0 48496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2366__A1
timestamp 1669390400
transform 1 0 52304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2366__A2
timestamp 1669390400
transform -1 0 51520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2368__A1
timestamp 1669390400
transform 1 0 52640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2368__A2
timestamp 1669390400
transform 1 0 52192 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2368__B
timestamp 1669390400
transform 1 0 51968 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2368__C
timestamp 1669390400
transform 1 0 52416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2369__B
timestamp 1669390400
transform 1 0 51744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2370__A1
timestamp 1669390400
transform 1 0 55104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2370__A2
timestamp 1669390400
transform 1 0 49392 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2371__A3
timestamp 1669390400
transform -1 0 51072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2372__A2
timestamp 1669390400
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2373__A1
timestamp 1669390400
transform 1 0 26544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2374__A1
timestamp 1669390400
transform 1 0 27104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2374__A2
timestamp 1669390400
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2379__I
timestamp 1669390400
transform 1 0 37856 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__A1
timestamp 1669390400
transform 1 0 40768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__A2
timestamp 1669390400
transform -1 0 41664 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2381__A1
timestamp 1669390400
transform -1 0 42560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2381__A2
timestamp 1669390400
transform -1 0 41664 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2382__A1
timestamp 1669390400
transform -1 0 49616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2382__B
timestamp 1669390400
transform 1 0 49840 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2384__A1
timestamp 1669390400
transform 1 0 36736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2384__A2
timestamp 1669390400
transform 1 0 37184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__A1
timestamp 1669390400
transform 1 0 46256 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__A2
timestamp 1669390400
transform 1 0 47152 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2386__I
timestamp 1669390400
transform 1 0 49504 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2387__A1
timestamp 1669390400
transform 1 0 48048 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2387__A2
timestamp 1669390400
transform 1 0 49392 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2388__A2
timestamp 1669390400
transform -1 0 38528 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2388__B2
timestamp 1669390400
transform -1 0 37632 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2388__C
timestamp 1669390400
transform -1 0 35840 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2389__B
timestamp 1669390400
transform -1 0 32480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2395__A1
timestamp 1669390400
transform 1 0 42784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2395__A2
timestamp 1669390400
transform 1 0 42336 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2396__I
timestamp 1669390400
transform 1 0 41440 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2397__A2
timestamp 1669390400
transform 1 0 40320 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2397__B1
timestamp 1669390400
transform 1 0 40768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2398__A1
timestamp 1669390400
transform -1 0 39872 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2399__A1
timestamp 1669390400
transform 1 0 45360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2399__A2
timestamp 1669390400
transform -1 0 45024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2399__B
timestamp 1669390400
transform 1 0 45360 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2400__A1
timestamp 1669390400
transform 1 0 43232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2401__A1
timestamp 1669390400
transform 1 0 47152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2401__A2
timestamp 1669390400
transform 1 0 47824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2402__A2
timestamp 1669390400
transform 1 0 41440 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2402__A3
timestamp 1669390400
transform 1 0 41104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2404__A1
timestamp 1669390400
transform -1 0 43792 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2404__A2
timestamp 1669390400
transform -1 0 42672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2405__A1
timestamp 1669390400
transform -1 0 42112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2407__B
timestamp 1669390400
transform -1 0 39984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2409__A1
timestamp 1669390400
transform -1 0 23520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2409__A2
timestamp 1669390400
transform 1 0 24752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2410__A1
timestamp 1669390400
transform 1 0 23744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2411__I
timestamp 1669390400
transform 1 0 32144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2412__I
timestamp 1669390400
transform 1 0 43120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2413__A1
timestamp 1669390400
transform 1 0 41440 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2413__A2
timestamp 1669390400
transform 1 0 44016 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2414__A1
timestamp 1669390400
transform 1 0 42560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2414__A2
timestamp 1669390400
transform 1 0 43680 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2416__A1
timestamp 1669390400
transform 1 0 42672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2416__A2
timestamp 1669390400
transform 1 0 43008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2417__A1
timestamp 1669390400
transform 1 0 50512 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2417__A2
timestamp 1669390400
transform 1 0 50848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2417__C
timestamp 1669390400
transform 1 0 51296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2418__A1
timestamp 1669390400
transform -1 0 29008 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2418__A2
timestamp 1669390400
transform 1 0 30576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2419__A2
timestamp 1669390400
transform 1 0 30688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2420__A2
timestamp 1669390400
transform -1 0 23184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2421__A1
timestamp 1669390400
transform 1 0 23408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2421__A2
timestamp 1669390400
transform 1 0 22960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2424__A1
timestamp 1669390400
transform 1 0 26656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2424__A2
timestamp 1669390400
transform 1 0 26656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2425__A2
timestamp 1669390400
transform -1 0 23632 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2428__A2
timestamp 1669390400
transform -1 0 22512 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2430__A1
timestamp 1669390400
transform 1 0 20832 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2430__A2
timestamp 1669390400
transform 1 0 23408 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2434__A1
timestamp 1669390400
transform 1 0 46704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2434__B
timestamp 1669390400
transform 1 0 45136 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2435__I
timestamp 1669390400
transform 1 0 38304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2436__A1
timestamp 1669390400
transform 1 0 41552 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2436__A2
timestamp 1669390400
transform 1 0 43568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2437__I
timestamp 1669390400
transform 1 0 38304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2438__A1
timestamp 1669390400
transform -1 0 41328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2438__C
timestamp 1669390400
transform 1 0 41552 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2439__A1
timestamp 1669390400
transform 1 0 51072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2439__A2
timestamp 1669390400
transform -1 0 45584 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2439__C
timestamp 1669390400
transform 1 0 49392 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2440__A1
timestamp 1669390400
transform 1 0 41888 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2442__A2
timestamp 1669390400
transform 1 0 30240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2443__A1
timestamp 1669390400
transform -1 0 27888 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2443__A2
timestamp 1669390400
transform 1 0 27328 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__I
timestamp 1669390400
transform 1 0 37856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2447__I
timestamp 1669390400
transform 1 0 32816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2448__A2
timestamp 1669390400
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2449__A1
timestamp 1669390400
transform 1 0 30800 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2450__A1
timestamp 1669390400
transform 1 0 37856 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2451__A1
timestamp 1669390400
transform 1 0 53312 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2451__B
timestamp 1669390400
transform 1 0 54656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2452__A1
timestamp 1669390400
transform 1 0 44576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2452__A2
timestamp 1669390400
transform -1 0 44352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2453__A1
timestamp 1669390400
transform 1 0 44352 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2453__A2
timestamp 1669390400
transform 1 0 44800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2453__B1
timestamp 1669390400
transform 1 0 45696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2453__B2
timestamp 1669390400
transform 1 0 45248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2454__I
timestamp 1669390400
transform -1 0 46032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2455__A2
timestamp 1669390400
transform 1 0 42896 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2455__B2
timestamp 1669390400
transform 1 0 50288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2455__C
timestamp 1669390400
transform 1 0 46144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2457__I
timestamp 1669390400
transform 1 0 36960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2460__A1
timestamp 1669390400
transform 1 0 39088 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2462__A2
timestamp 1669390400
transform 1 0 24752 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2462__B
timestamp 1669390400
transform 1 0 24304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2463__A1
timestamp 1669390400
transform 1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2463__A2
timestamp 1669390400
transform 1 0 41776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2463__B
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2464__A1
timestamp 1669390400
transform 1 0 39424 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2464__B
timestamp 1669390400
transform 1 0 39872 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2465__A1
timestamp 1669390400
transform 1 0 49840 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2465__A2
timestamp 1669390400
transform -1 0 47936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2467__A1
timestamp 1669390400
transform 1 0 37408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2467__A2
timestamp 1669390400
transform 1 0 37856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2469__A2
timestamp 1669390400
transform -1 0 23632 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2470__A2
timestamp 1669390400
transform 1 0 21952 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2470__A3
timestamp 1669390400
transform 1 0 21504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2471__A2
timestamp 1669390400
transform -1 0 19936 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2472__A2
timestamp 1669390400
transform 1 0 22624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2474__I
timestamp 1669390400
transform -1 0 3360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2476__A1
timestamp 1669390400
transform 1 0 35952 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2476__A2
timestamp 1669390400
transform 1 0 33488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__I
timestamp 1669390400
transform 1 0 39088 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2481__A2
timestamp 1669390400
transform -1 0 40432 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2482__A2
timestamp 1669390400
transform 1 0 37744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2483__A1
timestamp 1669390400
transform 1 0 46816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2483__A2
timestamp 1669390400
transform 1 0 46368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2483__B1
timestamp 1669390400
transform 1 0 48496 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2483__B2
timestamp 1669390400
transform 1 0 47264 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2484__A2
timestamp 1669390400
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2484__A3
timestamp 1669390400
transform 1 0 32816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2484__B
timestamp 1669390400
transform 1 0 30800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2485__A1
timestamp 1669390400
transform 1 0 37296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2485__B1
timestamp 1669390400
transform -1 0 34944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2486__A1
timestamp 1669390400
transform -1 0 31024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2486__A2
timestamp 1669390400
transform -1 0 30576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2488__A1
timestamp 1669390400
transform 1 0 30016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2490__I
timestamp 1669390400
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2491__I
timestamp 1669390400
transform 1 0 36288 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2492__I
timestamp 1669390400
transform 1 0 39760 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2494__A2
timestamp 1669390400
transform 1 0 36960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2495__I
timestamp 1669390400
transform 1 0 37408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2497__A2
timestamp 1669390400
transform 1 0 38192 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2498__A2
timestamp 1669390400
transform -1 0 37184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2499__A1
timestamp 1669390400
transform 1 0 38640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2500__A1
timestamp 1669390400
transform 1 0 35168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2500__A2
timestamp 1669390400
transform 1 0 36512 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2502__A4
timestamp 1669390400
transform -1 0 40432 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__I
timestamp 1669390400
transform 1 0 37184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2505__A4
timestamp 1669390400
transform -1 0 40992 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2506__A2
timestamp 1669390400
transform -1 0 34832 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2507__A1
timestamp 1669390400
transform 1 0 35168 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__A1
timestamp 1669390400
transform 1 0 30240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__A2
timestamp 1669390400
transform 1 0 30016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2509__I0
timestamp 1669390400
transform -1 0 30128 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2509__S
timestamp 1669390400
transform -1 0 29008 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2510__A1
timestamp 1669390400
transform -1 0 28336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2510__A2
timestamp 1669390400
transform -1 0 28784 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2510__A4
timestamp 1669390400
transform -1 0 30016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2513__I
timestamp 1669390400
transform -1 0 36960 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2514__A2
timestamp 1669390400
transform 1 0 41440 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2514__B
timestamp 1669390400
transform 1 0 41440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2515__A1
timestamp 1669390400
transform 1 0 36512 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2515__A2
timestamp 1669390400
transform 1 0 36960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__A1
timestamp 1669390400
transform 1 0 45360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2518__A1
timestamp 1669390400
transform -1 0 37408 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2518__B1
timestamp 1669390400
transform 1 0 37408 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__I1
timestamp 1669390400
transform 1 0 27104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__S
timestamp 1669390400
transform -1 0 23296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__A1
timestamp 1669390400
transform 1 0 17024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__A2
timestamp 1669390400
transform 1 0 16576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__A3
timestamp 1669390400
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2521__A1
timestamp 1669390400
transform 1 0 20160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2521__A2
timestamp 1669390400
transform 1 0 19712 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2522__A1
timestamp 1669390400
transform 1 0 20384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2522__A2
timestamp 1669390400
transform 1 0 19936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__A2
timestamp 1669390400
transform 1 0 26656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2526__B2
timestamp 1669390400
transform 1 0 25536 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2529__I
timestamp 1669390400
transform -1 0 56784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2530__A1
timestamp 1669390400
transform -1 0 13888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2530__A2
timestamp 1669390400
transform -1 0 14336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2531__A1
timestamp 1669390400
transform 1 0 17920 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2531__A2
timestamp 1669390400
transform -1 0 17696 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__A1
timestamp 1669390400
transform -1 0 14000 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2534__A1
timestamp 1669390400
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__A1
timestamp 1669390400
transform 1 0 41440 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__B2
timestamp 1669390400
transform 1 0 42224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__A1
timestamp 1669390400
transform -1 0 39536 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__A2
timestamp 1669390400
transform 1 0 40208 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2539__A2
timestamp 1669390400
transform 1 0 40096 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2540__A1
timestamp 1669390400
transform 1 0 38752 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2542__I
timestamp 1669390400
transform 1 0 36512 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2543__A1
timestamp 1669390400
transform -1 0 31472 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2544__A1
timestamp 1669390400
transform 1 0 33936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2544__B
timestamp 1669390400
transform 1 0 33488 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2544__C
timestamp 1669390400
transform -1 0 32256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2545__A1
timestamp 1669390400
transform 1 0 33152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2546__A2
timestamp 1669390400
transform 1 0 29568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2547__A2
timestamp 1669390400
transform 1 0 30240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2548__A1
timestamp 1669390400
transform 1 0 30576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2549__A1
timestamp 1669390400
transform 1 0 42000 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2551__A1
timestamp 1669390400
transform 1 0 36512 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2552__A1
timestamp 1669390400
transform -1 0 34272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2552__A3
timestamp 1669390400
transform 1 0 35840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2553__B
timestamp 1669390400
transform -1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2554__B
timestamp 1669390400
transform 1 0 36512 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2555__I
timestamp 1669390400
transform 1 0 36736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2556__B
timestamp 1669390400
transform 1 0 39312 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2557__A1
timestamp 1669390400
transform 1 0 24080 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2557__A2
timestamp 1669390400
transform -1 0 23856 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2558__A2
timestamp 1669390400
transform 1 0 32592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2559__A1
timestamp 1669390400
transform 1 0 36512 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2559__A2
timestamp 1669390400
transform 1 0 37856 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2560__A1
timestamp 1669390400
transform 1 0 36064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2560__B
timestamp 1669390400
transform -1 0 35840 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2561__A2
timestamp 1669390400
transform -1 0 32816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__A1
timestamp 1669390400
transform 1 0 32256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__A2
timestamp 1669390400
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2573__I
timestamp 1669390400
transform -1 0 3360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2574__A1
timestamp 1669390400
transform -1 0 28560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2575__A1
timestamp 1669390400
transform 1 0 39760 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__A1
timestamp 1669390400
transform 1 0 41888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__A2
timestamp 1669390400
transform 1 0 39536 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__B1
timestamp 1669390400
transform 1 0 42112 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2576__C
timestamp 1669390400
transform 1 0 38752 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2577__A1
timestamp 1669390400
transform 1 0 40768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2577__C
timestamp 1669390400
transform 1 0 37520 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2578__A2
timestamp 1669390400
transform 1 0 39536 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2578__A3
timestamp 1669390400
transform 1 0 39984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2579__A1
timestamp 1669390400
transform 1 0 29232 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2579__A2
timestamp 1669390400
transform -1 0 29904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2579__B
timestamp 1669390400
transform 1 0 28784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2580__A2
timestamp 1669390400
transform 1 0 27216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__A1
timestamp 1669390400
transform -1 0 39088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__A2
timestamp 1669390400
transform 1 0 39648 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__B2
timestamp 1669390400
transform 1 0 38416 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2583__C
timestamp 1669390400
transform 1 0 38864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__A2
timestamp 1669390400
transform 1 0 27664 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2586__A1
timestamp 1669390400
transform -1 0 37520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2587__A2
timestamp 1669390400
transform -1 0 38304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2587__A3
timestamp 1669390400
transform -1 0 37856 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__A2
timestamp 1669390400
transform -1 0 37184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2590__A1
timestamp 1669390400
transform 1 0 36736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2592__A1
timestamp 1669390400
transform 1 0 21504 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2592__A2
timestamp 1669390400
transform -1 0 21952 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2593__A1
timestamp 1669390400
transform -1 0 20608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__A1
timestamp 1669390400
transform 1 0 25200 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__A2
timestamp 1669390400
transform -1 0 24976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2604__A1
timestamp 1669390400
transform 1 0 20832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2604__A2
timestamp 1669390400
transform -1 0 20608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2605__A1
timestamp 1669390400
transform -1 0 18592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2606__I
timestamp 1669390400
transform 1 0 29568 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2607__I
timestamp 1669390400
transform -1 0 34160 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2608__A1
timestamp 1669390400
transform 1 0 33488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2608__B
timestamp 1669390400
transform 1 0 34608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2609__A1
timestamp 1669390400
transform -1 0 34832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2609__B1
timestamp 1669390400
transform 1 0 34160 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2610__I
timestamp 1669390400
transform 1 0 29904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__A1
timestamp 1669390400
transform -1 0 30464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__A2
timestamp 1669390400
transform 1 0 30688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2612__A1
timestamp 1669390400
transform -1 0 29680 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2613__A1
timestamp 1669390400
transform -1 0 29008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2614__A1
timestamp 1669390400
transform 1 0 29232 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2616__A1
timestamp 1669390400
transform 1 0 33488 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2617__A1
timestamp 1669390400
transform -1 0 35728 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2618__C
timestamp 1669390400
transform 1 0 33712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2621__A2
timestamp 1669390400
transform -1 0 33040 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2621__A3
timestamp 1669390400
transform -1 0 30576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2621__B
timestamp 1669390400
transform 1 0 31248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2623__A1
timestamp 1669390400
transform -1 0 25648 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2624__A1
timestamp 1669390400
transform 1 0 21504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2624__A2
timestamp 1669390400
transform -1 0 22624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2624__A3
timestamp 1669390400
transform 1 0 21952 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2632__I
timestamp 1669390400
transform 1 0 3136 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2633__A1
timestamp 1669390400
transform 1 0 35952 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2633__A2
timestamp 1669390400
transform 1 0 36400 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2634__A1
timestamp 1669390400
transform 1 0 32480 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2634__A3
timestamp 1669390400
transform 1 0 33712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__A1
timestamp 1669390400
transform 1 0 32816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2635__A4
timestamp 1669390400
transform 1 0 36736 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2637__A1
timestamp 1669390400
transform -1 0 26432 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__A1
timestamp 1669390400
transform 1 0 26432 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__A2
timestamp 1669390400
transform -1 0 22848 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2639__A1
timestamp 1669390400
transform 1 0 27440 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2639__A3
timestamp 1669390400
transform -1 0 25088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2641__A1
timestamp 1669390400
transform -1 0 24528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2641__B
timestamp 1669390400
transform 1 0 25872 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2643__A1
timestamp 1669390400
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__A1
timestamp 1669390400
transform -1 0 33488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__A2
timestamp 1669390400
transform 1 0 33712 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2645__A1
timestamp 1669390400
transform 1 0 34384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2645__B2
timestamp 1669390400
transform 1 0 30800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2646__A2
timestamp 1669390400
transform -1 0 31248 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2647__A1
timestamp 1669390400
transform 1 0 29792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2649__A1
timestamp 1669390400
transform -1 0 23072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2649__A2
timestamp 1669390400
transform -1 0 22848 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2650__A1
timestamp 1669390400
transform -1 0 21056 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2650__A2
timestamp 1669390400
transform -1 0 19712 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2651__A1
timestamp 1669390400
transform -1 0 21728 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2656__I
timestamp 1669390400
transform -1 0 3360 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2659__A1
timestamp 1669390400
transform 1 0 33936 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2659__B
timestamp 1669390400
transform 1 0 32816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__A1
timestamp 1669390400
transform 1 0 26096 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2669__I
timestamp 1669390400
transform 1 0 56672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2672__A1
timestamp 1669390400
transform 1 0 28672 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2679__I
timestamp 1669390400
transform -1 0 56784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__A2
timestamp 1669390400
transform 1 0 32480 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2682__A1
timestamp 1669390400
transform 1 0 30240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2682__A2
timestamp 1669390400
transform -1 0 30912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2683__I
timestamp 1669390400
transform 1 0 23968 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2684__I
timestamp 1669390400
transform 1 0 16016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2685__A1
timestamp 1669390400
transform 1 0 19712 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2685__A2
timestamp 1669390400
transform 1 0 17920 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2687__I
timestamp 1669390400
transform 1 0 26432 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2688__A2
timestamp 1669390400
transform 1 0 34496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2689__A1
timestamp 1669390400
transform -1 0 35504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2689__A2
timestamp 1669390400
transform 1 0 37408 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2689__A3
timestamp 1669390400
transform -1 0 35952 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__A2
timestamp 1669390400
transform 1 0 36064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__A3
timestamp 1669390400
transform 1 0 36176 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__A4
timestamp 1669390400
transform 1 0 36512 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2692__A1
timestamp 1669390400
transform 1 0 38192 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2692__A2
timestamp 1669390400
transform -1 0 37632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2693__A1
timestamp 1669390400
transform -1 0 30128 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2693__A2
timestamp 1669390400
transform -1 0 29904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2694__A1
timestamp 1669390400
transform 1 0 32704 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2696__A2
timestamp 1669390400
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2696__A3
timestamp 1669390400
transform 1 0 26992 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2697__A1
timestamp 1669390400
transform 1 0 32704 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2697__A2
timestamp 1669390400
transform 1 0 32480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2698__B
timestamp 1669390400
transform -1 0 35840 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2700__A1
timestamp 1669390400
transform 1 0 33488 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2701__A1
timestamp 1669390400
transform -1 0 31360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2702__A1
timestamp 1669390400
transform -1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2703__A1
timestamp 1669390400
transform -1 0 15568 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2703__A2
timestamp 1669390400
transform -1 0 13440 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__A1
timestamp 1669390400
transform 1 0 20272 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__A2
timestamp 1669390400
transform 1 0 21952 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__A1
timestamp 1669390400
transform 1 0 21504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__A2
timestamp 1669390400
transform -1 0 18368 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__A3
timestamp 1669390400
transform 1 0 19936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__A1
timestamp 1669390400
transform -1 0 16352 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__A3
timestamp 1669390400
transform 1 0 17584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__A4
timestamp 1669390400
transform 1 0 16912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2708__A1
timestamp 1669390400
transform -1 0 14672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2708__A2
timestamp 1669390400
transform 1 0 16016 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2708__B
timestamp 1669390400
transform -1 0 14224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__A1
timestamp 1669390400
transform -1 0 10528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2713__A1
timestamp 1669390400
transform -1 0 22064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2713__A2
timestamp 1669390400
transform 1 0 24080 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2714__A1
timestamp 1669390400
transform 1 0 23744 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2714__A2
timestamp 1669390400
transform -1 0 23520 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2715__A1
timestamp 1669390400
transform -1 0 18256 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2717__A1
timestamp 1669390400
transform 1 0 21616 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2718__A1
timestamp 1669390400
transform -1 0 22176 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2721__A1
timestamp 1669390400
transform 1 0 39984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2722__CLK
timestamp 1669390400
transform 1 0 37968 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2723__CLK
timestamp 1669390400
transform 1 0 37520 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2724__RN
timestamp 1669390400
transform 1 0 25872 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2725__RN
timestamp 1669390400
transform -1 0 25760 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2726__RN
timestamp 1669390400
transform 1 0 21504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2727__CLK
timestamp 1669390400
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2727__RN
timestamp 1669390400
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2730__CLK
timestamp 1669390400
transform -1 0 20832 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2731__CLK
timestamp 1669390400
transform 1 0 41440 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2732__CLK
timestamp 1669390400
transform 1 0 41104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2733__CLK
timestamp 1669390400
transform 1 0 30912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2733__RN
timestamp 1669390400
transform 1 0 31360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__CLK
timestamp 1669390400
transform 1 0 39424 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__D
timestamp 1669390400
transform 1 0 38976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2736__D
timestamp 1669390400
transform -1 0 35728 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2737__CLK
timestamp 1669390400
transform 1 0 28448 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2737__D
timestamp 1669390400
transform 1 0 28224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2737__RN
timestamp 1669390400
transform 1 0 28896 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2739__SETN
timestamp 1669390400
transform 1 0 18032 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2740__CLK
timestamp 1669390400
transform 1 0 22624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2740__RN
timestamp 1669390400
transform 1 0 22400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2741__RN
timestamp 1669390400
transform 1 0 17136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2742__SETN
timestamp 1669390400
transform 1 0 16240 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__CLK
timestamp 1669390400
transform 1 0 22400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__SETN
timestamp 1669390400
transform -1 0 24416 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2744__CLK
timestamp 1669390400
transform 1 0 22848 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2744__RN
timestamp 1669390400
transform 1 0 27328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2745__CLK
timestamp 1669390400
transform 1 0 31584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2745__D
timestamp 1669390400
transform 1 0 27104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2745__RN
timestamp 1669390400
transform 1 0 32032 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2747__D
timestamp 1669390400
transform -1 0 38080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout44_I
timestamp 1669390400
transform 1 0 29456 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout45_I
timestamp 1669390400
transform 1 0 27888 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout46_I
timestamp 1669390400
transform 1 0 34608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout47_I
timestamp 1669390400
transform -1 0 24192 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout48_I
timestamp 1669390400
transform -1 0 27888 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout49_I
timestamp 1669390400
transform -1 0 33824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout50_I
timestamp 1669390400
transform 1 0 24528 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout51_I
timestamp 1669390400
transform 1 0 13664 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout54_I
timestamp 1669390400
transform -1 0 20384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout55_I
timestamp 1669390400
transform 1 0 15792 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout58_I
timestamp 1669390400
transform -1 0 36848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout59_I
timestamp 1669390400
transform -1 0 30128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout60_I
timestamp 1669390400
transform -1 0 38528 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout61_I
timestamp 1669390400
transform 1 0 30352 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout62_I
timestamp 1669390400
transform -1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout63_I
timestamp 1669390400
transform -1 0 15344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout64_I
timestamp 1669390400
transform -1 0 21504 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout66_I
timestamp 1669390400
transform -1 0 38752 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout67_I
timestamp 1669390400
transform 1 0 41440 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout68_I
timestamp 1669390400
transform 1 0 43232 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform -1 0 27552 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform 1 0 43568 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform -1 0 44352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform -1 0 56448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform -1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output7_I
timestamp 1669390400
transform -1 0 2016 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output9_I
timestamp 1669390400
transform 1 0 54320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output13_I
timestamp 1669390400
transform -1 0 46256 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output18_I
timestamp 1669390400
transform 1 0 3696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output22_I
timestamp 1669390400
transform 1 0 56448 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output24_I
timestamp 1669390400
transform -1 0 33712 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output27_I
timestamp 1669390400
transform 1 0 54320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output32_I
timestamp 1669390400
transform -1 0 19376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output33_I
timestamp 1669390400
transform 1 0 35280 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output34_I
timestamp 1669390400
transform -1 0 56784 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output35_I
timestamp 1669390400
transform -1 0 26880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output36_I
timestamp 1669390400
transform 1 0 53872 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output37_I
timestamp 1669390400
transform 1 0 54320 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output38_I
timestamp 1669390400
transform -1 0 6160 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output39_I
timestamp 1669390400
transform 1 0 25648 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output40_I
timestamp 1669390400
transform 1 0 40880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output41_I
timestamp 1669390400
transform 1 0 3472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output42_I
timestamp 1669390400
transform 1 0 43120 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output43_I
timestamp 1669390400
transform 1 0 53536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3248 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4592 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31
timestamp 1669390400
transform 1 0 4816 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34
timestamp 1669390400
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1669390400
transform 1 0 5488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7392 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72
timestamp 1669390400
transform 1 0 9408 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80
timestamp 1669390400
transform 1 0 10304 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84
timestamp 1669390400
transform 1 0 10752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_99
timestamp 1669390400
transform 1 0 12432 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103
timestamp 1669390400
transform 1 0 12880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_107 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13328 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_157
timestamp 1669390400
transform 1 0 18928 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_161
timestamp 1669390400
transform 1 0 19376 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_169
timestamp 1669390400
transform 1 0 20272 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_173
timestamp 1669390400
transform 1 0 20720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_185
timestamp 1669390400
transform 1 0 22064 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_201
timestamp 1669390400
transform 1 0 23856 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_220
timestamp 1669390400
transform 1 0 25984 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_224
timestamp 1669390400
transform 1 0 26432 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_228
timestamp 1669390400
transform 1 0 26880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1669390400
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_260
timestamp 1669390400
transform 1 0 30464 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_276
timestamp 1669390400
transform 1 0 32256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_285
timestamp 1669390400
transform 1 0 33264 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_303
timestamp 1669390400
transform 1 0 35280 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_307
timestamp 1669390400
transform 1 0 35728 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_320
timestamp 1669390400
transform 1 0 37184 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_324
timestamp 1669390400
transform 1 0 37632 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_328
timestamp 1669390400
transform 1 0 38080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_332
timestamp 1669390400
transform 1 0 38528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_334
timestamp 1669390400
transform 1 0 38752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1669390400
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_355
timestamp 1669390400
transform 1 0 41104 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_371
timestamp 1669390400
transform 1 0 42896 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_379
timestamp 1669390400
transform 1 0 43792 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_381
timestamp 1669390400
transform 1 0 44016 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_384
timestamp 1669390400
transform 1 0 44352 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_394
timestamp 1669390400
transform 1 0 45472 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_410
timestamp 1669390400
transform 1 0 47264 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_414
timestamp 1669390400
transform 1 0 47712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_417
timestamp 1669390400
transform 1 0 48048 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1669390400
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_422
timestamp 1669390400
transform 1 0 48608 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_438
timestamp 1669390400
transform 1 0 50400 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_453
timestamp 1669390400
transform 1 0 52080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_457
timestamp 1669390400
transform 1 0 52528 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_473
timestamp 1669390400
transform 1 0 54320 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1669390400
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_492
timestamp 1669390400
transform 1 0 56448 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_508
timestamp 1669390400
transform 1 0 58240 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_2
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_6
timestamp 1669390400
transform 1 0 2016 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_14
timestamp 1669390400
transform 1 0 2912 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_18
timestamp 1669390400
transform 1 0 3360 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_50
timestamp 1669390400
transform 1 0 6944 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_66
timestamp 1669390400
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_73 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1669390400
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1669390400
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_176
timestamp 1669390400
transform 1 0 21056 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_178
timestamp 1669390400
transform 1 0 21280 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_203
timestamp 1669390400
transform 1 0 24080 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_211
timestamp 1669390400
transform 1 0 24976 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_219
timestamp 1669390400
transform 1 0 25872 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_221
timestamp 1669390400
transform 1 0 26096 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_228
timestamp 1669390400
transform 1 0 26880 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_236
timestamp 1669390400
transform 1 0 27776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_255
timestamp 1669390400
transform 1 0 29904 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_263
timestamp 1669390400
transform 1 0 30800 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_289
timestamp 1669390400
transform 1 0 33712 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_293
timestamp 1669390400
transform 1 0 34160 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_328
timestamp 1669390400
transform 1 0 38080 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_336
timestamp 1669390400
transform 1 0 38976 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_343
timestamp 1669390400
transform 1 0 39760 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_347
timestamp 1669390400
transform 1 0 40208 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_389
timestamp 1669390400
transform 1 0 44912 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_407
timestamp 1669390400
transform 1 0 46928 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_411
timestamp 1669390400
transform 1 0 47376 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_415
timestamp 1669390400
transform 1 0 47824 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_423
timestamp 1669390400
transform 1 0 48720 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1669390400
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_428
timestamp 1669390400
transform 1 0 49280 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_460
timestamp 1669390400
transform 1 0 52864 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_468
timestamp 1669390400
transform 1 0 53760 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_472
timestamp 1669390400
transform 1 0 54208 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_475
timestamp 1669390400
transform 1 0 54544 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_491
timestamp 1669390400
transform 1 0 56336 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_493
timestamp 1669390400
transform 1 0 56560 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1669390400
transform 1 0 56896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_499
timestamp 1669390400
transform 1 0 57232 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_506
timestamp 1669390400
transform 1 0 58016 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_508
timestamp 1669390400
transform 1 0 58240 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1669390400
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_140
timestamp 1669390400
transform 1 0 17024 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_156
timestamp 1669390400
transform 1 0 18816 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_164
timestamp 1669390400
transform 1 0 19712 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_168
timestamp 1669390400
transform 1 0 20160 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_190
timestamp 1669390400
transform 1 0 22624 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_207
timestamp 1669390400
transform 1 0 24528 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_217
timestamp 1669390400
transform 1 0 25648 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_233
timestamp 1669390400
transform 1 0 27440 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_258
timestamp 1669390400
transform 1 0 30240 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_262
timestamp 1669390400
transform 1 0 30688 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_264
timestamp 1669390400
transform 1 0 30912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_271
timestamp 1669390400
transform 1 0 31696 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_286
timestamp 1669390400
transform 1 0 33376 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_290
timestamp 1669390400
transform 1 0 33824 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_292
timestamp 1669390400
transform 1 0 34048 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_327
timestamp 1669390400
transform 1 0 37968 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_363
timestamp 1669390400
transform 1 0 42000 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_371
timestamp 1669390400
transform 1 0 42896 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_375
timestamp 1669390400
transform 1 0 43344 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_377
timestamp 1669390400
transform 1 0 43568 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_380
timestamp 1669390400
transform 1 0 43904 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_388
timestamp 1669390400
transform 1 0 44800 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_395
timestamp 1669390400
transform 1 0 45584 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_399
timestamp 1669390400
transform 1 0 46032 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_403
timestamp 1669390400
transform 1 0 46480 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_407
timestamp 1669390400
transform 1 0 46928 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_413
timestamp 1669390400
transform 1 0 47600 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_417
timestamp 1669390400
transform 1 0 48048 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_421
timestamp 1669390400
transform 1 0 48496 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_425
timestamp 1669390400
transform 1 0 48944 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_429
timestamp 1669390400
transform 1 0 49392 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_433
timestamp 1669390400
transform 1 0 49840 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_437
timestamp 1669390400
transform 1 0 50288 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_440
timestamp 1669390400
transform 1 0 50624 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_444
timestamp 1669390400
transform 1 0 51072 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_450
timestamp 1669390400
transform 1 0 51744 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_454
timestamp 1669390400
transform 1 0 52192 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_458
timestamp 1669390400
transform 1 0 52640 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1669390400
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_463
timestamp 1669390400
transform 1 0 53200 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_467
timestamp 1669390400
transform 1 0 53648 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_470
timestamp 1669390400
transform 1 0 53984 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_474
timestamp 1669390400
transform 1 0 54432 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_478
timestamp 1669390400
transform 1 0 54880 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_482
timestamp 1669390400
transform 1 0 55328 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_486
timestamp 1669390400
transform 1 0 55776 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_502
timestamp 1669390400
transform 1 0 57568 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_506
timestamp 1669390400
transform 1 0 58016 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_508
timestamp 1669390400
transform 1 0 58240 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_17
timestamp 1669390400
transform 1 0 3248 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_49
timestamp 1669390400
transform 1 0 6832 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_65
timestamp 1669390400
transform 1 0 8624 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_69
timestamp 1669390400
transform 1 0 9072 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1669390400
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_160
timestamp 1669390400
transform 1 0 19264 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_168
timestamp 1669390400
transform 1 0 20160 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_175
timestamp 1669390400
transform 1 0 20944 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_183
timestamp 1669390400
transform 1 0 21840 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_190
timestamp 1669390400
transform 1 0 22624 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_198
timestamp 1669390400
transform 1 0 23520 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_202
timestamp 1669390400
transform 1 0 23968 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_210
timestamp 1669390400
transform 1 0 24864 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_223
timestamp 1669390400
transform 1 0 26320 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_227
timestamp 1669390400
transform 1 0 26768 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_229
timestamp 1669390400
transform 1 0 26992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_236
timestamp 1669390400
transform 1 0 27776 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_246
timestamp 1669390400
transform 1 0 28896 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_254
timestamp 1669390400
transform 1 0 29792 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_258
timestamp 1669390400
transform 1 0 30240 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1669390400
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_295
timestamp 1669390400
transform 1 0 34384 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_299
timestamp 1669390400
transform 1 0 34832 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_313
timestamp 1669390400
transform 1 0 36400 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_317
timestamp 1669390400
transform 1 0 36848 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_319
timestamp 1669390400
transform 1 0 37072 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1669390400
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_365
timestamp 1669390400
transform 1 0 42224 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_373
timestamp 1669390400
transform 1 0 43120 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_381
timestamp 1669390400
transform 1 0 44016 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_387
timestamp 1669390400
transform 1 0 44688 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_389
timestamp 1669390400
transform 1 0 44912 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_396
timestamp 1669390400
transform 1 0 45696 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_400
timestamp 1669390400
transform 1 0 46144 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_404
timestamp 1669390400
transform 1 0 46592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_408
timestamp 1669390400
transform 1 0 47040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_411
timestamp 1669390400
transform 1 0 47376 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_415
timestamp 1669390400
transform 1 0 47824 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_418
timestamp 1669390400
transform 1 0 48160 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_422
timestamp 1669390400
transform 1 0 48608 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_428
timestamp 1669390400
transform 1 0 49280 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_435
timestamp 1669390400
transform 1 0 50064 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_439
timestamp 1669390400
transform 1 0 50512 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_443
timestamp 1669390400
transform 1 0 50960 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_447
timestamp 1669390400
transform 1 0 51408 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_451
timestamp 1669390400
transform 1 0 51856 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_455
timestamp 1669390400
transform 1 0 52304 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_458
timestamp 1669390400
transform 1 0 52640 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_462
timestamp 1669390400
transform 1 0 53088 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_466
timestamp 1669390400
transform 1 0 53536 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_470
timestamp 1669390400
transform 1 0 53984 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_472
timestamp 1669390400
transform 1 0 54208 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_475
timestamp 1669390400
transform 1 0 54544 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_479
timestamp 1669390400
transform 1 0 54992 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_483
timestamp 1669390400
transform 1 0 55440 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_485
timestamp 1669390400
transform 1 0 55664 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_488
timestamp 1669390400
transform 1 0 56000 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_492
timestamp 1669390400
transform 1 0 56448 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1669390400
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_499
timestamp 1669390400
transform 1 0 57232 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_502
timestamp 1669390400
transform 1 0 57568 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_506
timestamp 1669390400
transform 1 0 58016 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_508
timestamp 1669390400
transform 1 0 58240 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_6
timestamp 1669390400
transform 1 0 2016 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_14
timestamp 1669390400
transform 1 0 2912 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_18
timestamp 1669390400
transform 1 0 3360 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1669390400
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_140
timestamp 1669390400
transform 1 0 17024 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_156
timestamp 1669390400
transform 1 0 18816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_170
timestamp 1669390400
transform 1 0 20384 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_182
timestamp 1669390400
transform 1 0 21728 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_190
timestamp 1669390400
transform 1 0 22624 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_199
timestamp 1669390400
transform 1 0 23632 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_209
timestamp 1669390400
transform 1 0 24752 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_225
timestamp 1669390400
transform 1 0 26544 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_235
timestamp 1669390400
transform 1 0 27664 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_241
timestamp 1669390400
transform 1 0 28336 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_243
timestamp 1669390400
transform 1 0 28560 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_246
timestamp 1669390400
transform 1 0 28896 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_253
timestamp 1669390400
transform 1 0 29680 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_257
timestamp 1669390400
transform 1 0 30128 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_259
timestamp 1669390400
transform 1 0 30352 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_265
timestamp 1669390400
transform 1 0 31024 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_278
timestamp 1669390400
transform 1 0 32480 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_288
timestamp 1669390400
transform 1 0 33600 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_292
timestamp 1669390400
transform 1 0 34048 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_298
timestamp 1669390400
transform 1 0 34720 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_308
timestamp 1669390400
transform 1 0 35840 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_316
timestamp 1669390400
transform 1 0 36736 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1669390400
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_324
timestamp 1669390400
transform 1 0 37632 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_328
timestamp 1669390400
transform 1 0 38080 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_363
timestamp 1669390400
transform 1 0 42000 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_367
timestamp 1669390400
transform 1 0 42448 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_370
timestamp 1669390400
transform 1 0 42784 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_374
timestamp 1669390400
transform 1 0 43232 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_378
timestamp 1669390400
transform 1 0 43680 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_386
timestamp 1669390400
transform 1 0 44576 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_395
timestamp 1669390400
transform 1 0 45584 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_397
timestamp 1669390400
transform 1 0 45808 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_410
timestamp 1669390400
transform 1 0 47264 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_414
timestamp 1669390400
transform 1 0 47712 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_423
timestamp 1669390400
transform 1 0 48720 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_449
timestamp 1669390400
transform 1 0 51632 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_451
timestamp 1669390400
transform 1 0 51856 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_454
timestamp 1669390400
transform 1 0 52192 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_458
timestamp 1669390400
transform 1 0 52640 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1669390400
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_463
timestamp 1669390400
transform 1 0 53200 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_466
timestamp 1669390400
transform 1 0 53536 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_470
timestamp 1669390400
transform 1 0 53984 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_474
timestamp 1669390400
transform 1 0 54432 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_478
timestamp 1669390400
transform 1 0 54880 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_484
timestamp 1669390400
transform 1 0 55552 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_492
timestamp 1669390400
transform 1 0 56448 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_496
timestamp 1669390400
transform 1 0 56896 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_500
timestamp 1669390400
transform 1 0 57344 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_502
timestamp 1669390400
transform 1 0 57568 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_505
timestamp 1669390400
transform 1 0 57904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1669390400
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1669390400
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1669390400
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_153
timestamp 1669390400
transform 1 0 18480 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_161
timestamp 1669390400
transform 1 0 19376 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_165
timestamp 1669390400
transform 1 0 19824 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_174
timestamp 1669390400
transform 1 0 20832 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_190
timestamp 1669390400
transform 1 0 22624 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_204
timestamp 1669390400
transform 1 0 24192 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1669390400
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_220
timestamp 1669390400
transform 1 0 25984 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_222
timestamp 1669390400
transform 1 0 26208 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_235
timestamp 1669390400
transform 1 0 27664 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_237
timestamp 1669390400
transform 1 0 27888 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_244
timestamp 1669390400
transform 1 0 28672 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_252
timestamp 1669390400
transform 1 0 29568 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_256
timestamp 1669390400
transform 1 0 30016 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_266
timestamp 1669390400
transform 1 0 31136 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_277
timestamp 1669390400
transform 1 0 32368 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_281
timestamp 1669390400
transform 1 0 32816 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1669390400
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_294
timestamp 1669390400
transform 1 0 34272 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_298
timestamp 1669390400
transform 1 0 34720 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_308
timestamp 1669390400
transform 1 0 35840 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_316
timestamp 1669390400
transform 1 0 36736 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_320
timestamp 1669390400
transform 1 0 37184 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_324
timestamp 1669390400
transform 1 0 37632 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_328
timestamp 1669390400
transform 1 0 38080 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_332
timestamp 1669390400
transform 1 0 38528 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_348
timestamp 1669390400
transform 1 0 40320 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_352
timestamp 1669390400
transform 1 0 40768 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_373
timestamp 1669390400
transform 1 0 43120 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_381
timestamp 1669390400
transform 1 0 44016 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_385
timestamp 1669390400
transform 1 0 44464 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_391
timestamp 1669390400
transform 1 0 45136 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_401
timestamp 1669390400
transform 1 0 46256 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_413
timestamp 1669390400
transform 1 0 47600 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_422
timestamp 1669390400
transform 1 0 48608 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_428
timestamp 1669390400
transform 1 0 49280 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_434
timestamp 1669390400
transform 1 0 49952 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_438
timestamp 1669390400
transform 1 0 50400 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_442
timestamp 1669390400
transform 1 0 50848 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_446
timestamp 1669390400
transform 1 0 51296 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_450
timestamp 1669390400
transform 1 0 51744 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_454
timestamp 1669390400
transform 1 0 52192 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_456
timestamp 1669390400
transform 1 0 52416 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_470
timestamp 1669390400
transform 1 0 53984 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_474
timestamp 1669390400
transform 1 0 54432 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_476
timestamp 1669390400
transform 1 0 54656 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_491
timestamp 1669390400
transform 1 0 56336 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_493
timestamp 1669390400
transform 1 0 56560 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1669390400
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_499
timestamp 1669390400
transform 1 0 57232 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_501
timestamp 1669390400
transform 1 0 57456 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_504
timestamp 1669390400
transform 1 0 57792 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_508
timestamp 1669390400
transform 1 0 58240 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1669390400
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_124
timestamp 1669390400
transform 1 0 15232 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_132
timestamp 1669390400
transform 1 0 16128 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_146
timestamp 1669390400
transform 1 0 17696 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_158
timestamp 1669390400
transform 1 0 19040 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_164
timestamp 1669390400
transform 1 0 19712 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_174
timestamp 1669390400
transform 1 0 20832 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_188
timestamp 1669390400
transform 1 0 22400 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_192
timestamp 1669390400
transform 1 0 22848 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_202
timestamp 1669390400
transform 1 0 23968 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_204
timestamp 1669390400
transform 1 0 24192 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_207
timestamp 1669390400
transform 1 0 24528 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_217
timestamp 1669390400
transform 1 0 25648 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_221
timestamp 1669390400
transform 1 0 26096 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_232
timestamp 1669390400
transform 1 0 27328 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_239
timestamp 1669390400
transform 1 0 28112 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1669390400
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1669390400
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_263
timestamp 1669390400
transform 1 0 30800 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_267
timestamp 1669390400
transform 1 0 31248 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_275
timestamp 1669390400
transform 1 0 32144 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_279
timestamp 1669390400
transform 1 0 32592 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_287
timestamp 1669390400
transform 1 0 33488 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_306
timestamp 1669390400
transform 1 0 35616 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_310
timestamp 1669390400
transform 1 0 36064 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_316
timestamp 1669390400
transform 1 0 36736 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_328
timestamp 1669390400
transform 1 0 38080 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_332
timestamp 1669390400
transform 1 0 38528 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_341
timestamp 1669390400
transform 1 0 39536 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_345
timestamp 1669390400
transform 1 0 39984 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_361
timestamp 1669390400
transform 1 0 41776 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_363
timestamp 1669390400
transform 1 0 42000 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_366
timestamp 1669390400
transform 1 0 42336 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_378
timestamp 1669390400
transform 1 0 43680 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_386
timestamp 1669390400
transform 1 0 44576 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_399
timestamp 1669390400
transform 1 0 46032 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_411
timestamp 1669390400
transform 1 0 47376 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_419
timestamp 1669390400
transform 1 0 48272 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_423
timestamp 1669390400
transform 1 0 48720 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_427
timestamp 1669390400
transform 1 0 49168 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_431
timestamp 1669390400
transform 1 0 49616 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_435
timestamp 1669390400
transform 1 0 50064 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_439
timestamp 1669390400
transform 1 0 50512 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_441
timestamp 1669390400
transform 1 0 50736 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_444
timestamp 1669390400
transform 1 0 51072 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_453
timestamp 1669390400
transform 1 0 52080 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1669390400
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_463
timestamp 1669390400
transform 1 0 53200 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_477
timestamp 1669390400
transform 1 0 54768 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_484
timestamp 1669390400
transform 1 0 55552 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_488
timestamp 1669390400
transform 1 0 56000 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_492
timestamp 1669390400
transform 1 0 56448 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_498
timestamp 1669390400
transform 1 0 57120 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_502
timestamp 1669390400
transform 1 0 57568 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_508
timestamp 1669390400
transform 1 0 58240 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1669390400
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_89
timestamp 1669390400
transform 1 0 11312 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_97
timestamp 1669390400
transform 1 0 12208 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_99
timestamp 1669390400
transform 1 0 12432 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_106
timestamp 1669390400
transform 1 0 13216 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_138
timestamp 1669390400
transform 1 0 16800 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_152
timestamp 1669390400
transform 1 0 18368 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_180
timestamp 1669390400
transform 1 0 21504 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_186
timestamp 1669390400
transform 1 0 22176 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_190
timestamp 1669390400
transform 1 0 22624 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_194
timestamp 1669390400
transform 1 0 23072 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_223
timestamp 1669390400
transform 1 0 26320 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_231
timestamp 1669390400
transform 1 0 27216 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_235
timestamp 1669390400
transform 1 0 27664 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_243
timestamp 1669390400
transform 1 0 28560 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_245
timestamp 1669390400
transform 1 0 28784 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_248
timestamp 1669390400
transform 1 0 29120 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_273
timestamp 1669390400
transform 1 0 31920 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_277
timestamp 1669390400
transform 1 0 32368 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_297
timestamp 1669390400
transform 1 0 34608 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_307
timestamp 1669390400
transform 1 0 35728 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_314
timestamp 1669390400
transform 1 0 36512 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_318
timestamp 1669390400
transform 1 0 36960 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_322
timestamp 1669390400
transform 1 0 37408 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_326
timestamp 1669390400
transform 1 0 37856 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_335
timestamp 1669390400
transform 1 0 38864 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_345
timestamp 1669390400
transform 1 0 39984 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_349
timestamp 1669390400
transform 1 0 40432 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_351
timestamp 1669390400
transform 1 0 40656 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_365
timestamp 1669390400
transform 1 0 42224 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_380
timestamp 1669390400
transform 1 0 43904 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_384
timestamp 1669390400
transform 1 0 44352 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_397
timestamp 1669390400
transform 1 0 45808 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_401
timestamp 1669390400
transform 1 0 46256 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_405
timestamp 1669390400
transform 1 0 46704 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_419
timestamp 1669390400
transform 1 0 48272 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_423
timestamp 1669390400
transform 1 0 48720 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1669390400
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_428
timestamp 1669390400
transform 1 0 49280 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_444
timestamp 1669390400
transform 1 0 51072 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_448
timestamp 1669390400
transform 1 0 51520 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_452
timestamp 1669390400
transform 1 0 51968 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_468
timestamp 1669390400
transform 1 0 53760 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_482
timestamp 1669390400
transform 1 0 55328 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_486
timestamp 1669390400
transform 1 0 55776 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_490
timestamp 1669390400
transform 1 0 56224 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_494
timestamp 1669390400
transform 1 0 56672 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1669390400
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_499
timestamp 1669390400
transform 1 0 57232 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_502
timestamp 1669390400
transform 1 0 57568 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_508
timestamp 1669390400
transform 1 0 58240 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_6
timestamp 1669390400
transform 1 0 2016 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_14
timestamp 1669390400
transform 1 0 2912 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_18
timestamp 1669390400
transform 1 0 3360 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1669390400
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_123
timestamp 1669390400
transform 1 0 15120 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_125
timestamp 1669390400
transform 1 0 15344 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_138
timestamp 1669390400
transform 1 0 16800 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_142
timestamp 1669390400
transform 1 0 17248 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_149
timestamp 1669390400
transform 1 0 18032 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_165
timestamp 1669390400
transform 1 0 19824 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_173
timestamp 1669390400
transform 1 0 20720 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_182
timestamp 1669390400
transform 1 0 21728 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_190
timestamp 1669390400
transform 1 0 22624 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_197
timestamp 1669390400
transform 1 0 23408 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_201
timestamp 1669390400
transform 1 0 23856 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_205
timestamp 1669390400
transform 1 0 24304 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_211
timestamp 1669390400
transform 1 0 24976 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_215
timestamp 1669390400
transform 1 0 25424 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_224
timestamp 1669390400
transform 1 0 26432 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_228
timestamp 1669390400
transform 1 0 26880 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_232
timestamp 1669390400
transform 1 0 27328 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_240
timestamp 1669390400
transform 1 0 28224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_244
timestamp 1669390400
transform 1 0 28672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_259
timestamp 1669390400
transform 1 0 30352 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_263
timestamp 1669390400
transform 1 0 30800 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_271
timestamp 1669390400
transform 1 0 31696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_275
timestamp 1669390400
transform 1 0 32144 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_277
timestamp 1669390400
transform 1 0 32368 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_280
timestamp 1669390400
transform 1 0 32704 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_293
timestamp 1669390400
transform 1 0 34160 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_301
timestamp 1669390400
transform 1 0 35056 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_314
timestamp 1669390400
transform 1 0 36512 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1669390400
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_337
timestamp 1669390400
transform 1 0 39088 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_341
timestamp 1669390400
transform 1 0 39536 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_343
timestamp 1669390400
transform 1 0 39760 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_360
timestamp 1669390400
transform 1 0 41664 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_373
timestamp 1669390400
transform 1 0 43120 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_381
timestamp 1669390400
transform 1 0 44016 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1669390400
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_395
timestamp 1669390400
transform 1 0 45584 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_401
timestamp 1669390400
transform 1 0 46256 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_405
timestamp 1669390400
transform 1 0 46704 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_415
timestamp 1669390400
transform 1 0 47824 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_419
timestamp 1669390400
transform 1 0 48272 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_423
timestamp 1669390400
transform 1 0 48720 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_427
timestamp 1669390400
transform 1 0 49168 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_442
timestamp 1669390400
transform 1 0 50848 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_450
timestamp 1669390400
transform 1 0 51744 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_454
timestamp 1669390400
transform 1 0 52192 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_458
timestamp 1669390400
transform 1 0 52640 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1669390400
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_463
timestamp 1669390400
transform 1 0 53200 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_466
timestamp 1669390400
transform 1 0 53536 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_470
timestamp 1669390400
transform 1 0 53984 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_474
timestamp 1669390400
transform 1 0 54432 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_478
timestamp 1669390400
transform 1 0 54880 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_482
timestamp 1669390400
transform 1 0 55328 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_486
timestamp 1669390400
transform 1 0 55776 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_490
timestamp 1669390400
transform 1 0 56224 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_494
timestamp 1669390400
transform 1 0 56672 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_498
timestamp 1669390400
transform 1 0 57120 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_502
timestamp 1669390400
transform 1 0 57568 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_508
timestamp 1669390400
transform 1 0 58240 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_6
timestamp 1669390400
transform 1 0 2016 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_14
timestamp 1669390400
transform 1 0 2912 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_18
timestamp 1669390400
transform 1 0 3360 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_50
timestamp 1669390400
transform 1 0 6944 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1669390400
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_105
timestamp 1669390400
transform 1 0 13104 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_113
timestamp 1669390400
transform 1 0 14000 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_117
timestamp 1669390400
transform 1 0 14448 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_124
timestamp 1669390400
transform 1 0 15232 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_134
timestamp 1669390400
transform 1 0 16352 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_153
timestamp 1669390400
transform 1 0 18480 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_157
timestamp 1669390400
transform 1 0 18928 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_166
timestamp 1669390400
transform 1 0 19936 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_182
timestamp 1669390400
transform 1 0 21728 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_186
timestamp 1669390400
transform 1 0 22176 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_207
timestamp 1669390400
transform 1 0 24528 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_209
timestamp 1669390400
transform 1 0 24752 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1669390400
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_228
timestamp 1669390400
transform 1 0 26880 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_238
timestamp 1669390400
transform 1 0 28000 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_240
timestamp 1669390400
transform 1 0 28224 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_255
timestamp 1669390400
transform 1 0 29904 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_271
timestamp 1669390400
transform 1 0 31696 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_279
timestamp 1669390400
transform 1 0 32592 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_288
timestamp 1669390400
transform 1 0 33600 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_291
timestamp 1669390400
transform 1 0 33936 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_301
timestamp 1669390400
transform 1 0 35056 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_305
timestamp 1669390400
transform 1 0 35504 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_312
timestamp 1669390400
transform 1 0 36288 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_316
timestamp 1669390400
transform 1 0 36736 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_320
timestamp 1669390400
transform 1 0 37184 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_327
timestamp 1669390400
transform 1 0 37968 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_335
timestamp 1669390400
transform 1 0 38864 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_342
timestamp 1669390400
transform 1 0 39648 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_352
timestamp 1669390400
transform 1 0 40768 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_360
timestamp 1669390400
transform 1 0 41664 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_364
timestamp 1669390400
transform 1 0 42112 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_368
timestamp 1669390400
transform 1 0 42560 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_372
timestamp 1669390400
transform 1 0 43008 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_376
timestamp 1669390400
transform 1 0 43456 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_380
timestamp 1669390400
transform 1 0 43904 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_386
timestamp 1669390400
transform 1 0 44576 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_393
timestamp 1669390400
transform 1 0 45360 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_397
timestamp 1669390400
transform 1 0 45808 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_401
timestamp 1669390400
transform 1 0 46256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_407
timestamp 1669390400
transform 1 0 46928 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_411
timestamp 1669390400
transform 1 0 47376 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_415
timestamp 1669390400
transform 1 0 47824 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_419
timestamp 1669390400
transform 1 0 48272 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_423
timestamp 1669390400
transform 1 0 48720 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1669390400
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_428
timestamp 1669390400
transform 1 0 49280 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_431
timestamp 1669390400
transform 1 0 49616 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_441
timestamp 1669390400
transform 1 0 50736 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_448
timestamp 1669390400
transform 1 0 51520 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_452
timestamp 1669390400
transform 1 0 51968 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_456
timestamp 1669390400
transform 1 0 52416 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_462
timestamp 1669390400
transform 1 0 53088 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_469
timestamp 1669390400
transform 1 0 53872 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_473
timestamp 1669390400
transform 1 0 54320 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_477
timestamp 1669390400
transform 1 0 54768 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_479
timestamp 1669390400
transform 1 0 54992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_482
timestamp 1669390400
transform 1 0 55328 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_486
timestamp 1669390400
transform 1 0 55776 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_490
timestamp 1669390400
transform 1 0 56224 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_494
timestamp 1669390400
transform 1 0 56672 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1669390400
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_499
timestamp 1669390400
transform 1 0 57232 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_502
timestamp 1669390400
transform 1 0 57568 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_506
timestamp 1669390400
transform 1 0 58016 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_508
timestamp 1669390400
transform 1 0 58240 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_17
timestamp 1669390400
transform 1 0 3248 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_33
timestamp 1669390400
transform 1 0 5040 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1669390400
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_112
timestamp 1669390400
transform 1 0 13888 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_126
timestamp 1669390400
transform 1 0 15456 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_133
timestamp 1669390400
transform 1 0 16240 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_153
timestamp 1669390400
transform 1 0 18480 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_157
timestamp 1669390400
transform 1 0 18928 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_168
timestamp 1669390400
transform 1 0 20160 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1669390400
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1669390400
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_181
timestamp 1669390400
transform 1 0 21616 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_184
timestamp 1669390400
transform 1 0 21952 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_199
timestamp 1669390400
transform 1 0 23632 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_206
timestamp 1669390400
transform 1 0 24416 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_208
timestamp 1669390400
transform 1 0 24640 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_224
timestamp 1669390400
transform 1 0 26432 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_228
timestamp 1669390400
transform 1 0 26880 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_232
timestamp 1669390400
transform 1 0 27328 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_241
timestamp 1669390400
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_257
timestamp 1669390400
transform 1 0 30128 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_259
timestamp 1669390400
transform 1 0 30352 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_262
timestamp 1669390400
transform 1 0 30688 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_270
timestamp 1669390400
transform 1 0 31584 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_282
timestamp 1669390400
transform 1 0 32928 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_286
timestamp 1669390400
transform 1 0 33376 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_290
timestamp 1669390400
transform 1 0 33824 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_294
timestamp 1669390400
transform 1 0 34272 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_302
timestamp 1669390400
transform 1 0 35168 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_314
timestamp 1669390400
transform 1 0 36512 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1669390400
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_328
timestamp 1669390400
transform 1 0 38080 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_332
timestamp 1669390400
transform 1 0 38528 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_335
timestamp 1669390400
transform 1 0 38864 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_339
timestamp 1669390400
transform 1 0 39312 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_341
timestamp 1669390400
transform 1 0 39536 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_344
timestamp 1669390400
transform 1 0 39872 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_348
timestamp 1669390400
transform 1 0 40320 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_352
timestamp 1669390400
transform 1 0 40768 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_354
timestamp 1669390400
transform 1 0 40992 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_357
timestamp 1669390400
transform 1 0 41328 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_361
timestamp 1669390400
transform 1 0 41776 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_365
timestamp 1669390400
transform 1 0 42224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_377
timestamp 1669390400
transform 1 0 43568 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1669390400
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_402
timestamp 1669390400
transform 1 0 46368 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_404
timestamp 1669390400
transform 1 0 46592 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_409
timestamp 1669390400
transform 1 0 47152 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_413
timestamp 1669390400
transform 1 0 47600 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_417
timestamp 1669390400
transform 1 0 48048 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_421
timestamp 1669390400
transform 1 0 48496 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_425
timestamp 1669390400
transform 1 0 48944 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_429
timestamp 1669390400
transform 1 0 49392 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_442
timestamp 1669390400
transform 1 0 50848 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_446
timestamp 1669390400
transform 1 0 51296 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_450
timestamp 1669390400
transform 1 0 51744 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_454
timestamp 1669390400
transform 1 0 52192 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_459
timestamp 1669390400
transform 1 0 52752 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_463
timestamp 1669390400
transform 1 0 53200 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_473
timestamp 1669390400
transform 1 0 54320 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_477
timestamp 1669390400
transform 1 0 54768 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_481
timestamp 1669390400
transform 1 0 55216 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_485
timestamp 1669390400
transform 1 0 55664 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_489
timestamp 1669390400
transform 1 0 56112 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_493
timestamp 1669390400
transform 1 0 56560 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_497
timestamp 1669390400
transform 1 0 57008 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_501
timestamp 1669390400
transform 1 0 57456 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_505
timestamp 1669390400
transform 1 0 57904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_6
timestamp 1669390400
transform 1 0 2016 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_14
timestamp 1669390400
transform 1 0 2912 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_18
timestamp 1669390400
transform 1 0 3360 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_50
timestamp 1669390400
transform 1 0 6944 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1669390400
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1669390400
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_105
timestamp 1669390400
transform 1 0 13104 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_121
timestamp 1669390400
transform 1 0 14896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_130
timestamp 1669390400
transform 1 0 15904 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_138
timestamp 1669390400
transform 1 0 16800 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_152
timestamp 1669390400
transform 1 0 18368 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_166
timestamp 1669390400
transform 1 0 19936 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_180
timestamp 1669390400
transform 1 0 21504 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_182
timestamp 1669390400
transform 1 0 21728 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_195
timestamp 1669390400
transform 1 0 23184 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_203
timestamp 1669390400
transform 1 0 24080 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_207
timestamp 1669390400
transform 1 0 24528 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_209
timestamp 1669390400
transform 1 0 24752 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_217
timestamp 1669390400
transform 1 0 25648 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_228
timestamp 1669390400
transform 1 0 26880 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_236
timestamp 1669390400
transform 1 0 27776 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_238
timestamp 1669390400
transform 1 0 28000 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_247
timestamp 1669390400
transform 1 0 29008 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_251
timestamp 1669390400
transform 1 0 29456 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_253
timestamp 1669390400
transform 1 0 29680 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_256
timestamp 1669390400
transform 1 0 30016 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_262
timestamp 1669390400
transform 1 0 30688 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_274
timestamp 1669390400
transform 1 0 32032 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_282
timestamp 1669390400
transform 1 0 32928 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_289
timestamp 1669390400
transform 1 0 33712 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_293
timestamp 1669390400
transform 1 0 34160 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_299
timestamp 1669390400
transform 1 0 34832 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_312
timestamp 1669390400
transform 1 0 36288 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_324
timestamp 1669390400
transform 1 0 37632 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_332
timestamp 1669390400
transform 1 0 38528 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_336
timestamp 1669390400
transform 1 0 38976 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_340
timestamp 1669390400
transform 1 0 39424 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_344
timestamp 1669390400
transform 1 0 39872 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_348
timestamp 1669390400
transform 1 0 40320 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_352
timestamp 1669390400
transform 1 0 40768 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_360
timestamp 1669390400
transform 1 0 41664 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_364
timestamp 1669390400
transform 1 0 42112 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_366
timestamp 1669390400
transform 1 0 42336 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_375
timestamp 1669390400
transform 1 0 43344 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_379
timestamp 1669390400
transform 1 0 43792 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_406
timestamp 1669390400
transform 1 0 46816 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_416
timestamp 1669390400
transform 1 0 47936 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_420
timestamp 1669390400
transform 1 0 48384 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_422
timestamp 1669390400
transform 1 0 48608 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1669390400
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_428
timestamp 1669390400
transform 1 0 49280 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_437
timestamp 1669390400
transform 1 0 50288 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_445
timestamp 1669390400
transform 1 0 51184 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_452
timestamp 1669390400
transform 1 0 51968 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_456
timestamp 1669390400
transform 1 0 52416 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_460
timestamp 1669390400
transform 1 0 52864 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_462
timestamp 1669390400
transform 1 0 53088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_468
timestamp 1669390400
transform 1 0 53760 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_474
timestamp 1669390400
transform 1 0 54432 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_478
timestamp 1669390400
transform 1 0 54880 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_482
timestamp 1669390400
transform 1 0 55328 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_486
timestamp 1669390400
transform 1 0 55776 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_490
timestamp 1669390400
transform 1 0 56224 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_494
timestamp 1669390400
transform 1 0 56672 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1669390400
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_499
timestamp 1669390400
transform 1 0 57232 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_502
timestamp 1669390400
transform 1 0 57568 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_506
timestamp 1669390400
transform 1 0 58016 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_508
timestamp 1669390400
transform 1 0 58240 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1669390400
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1669390400
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1669390400
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_116
timestamp 1669390400
transform 1 0 14336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_120
timestamp 1669390400
transform 1 0 14784 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_131
timestamp 1669390400
transform 1 0 16016 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_137
timestamp 1669390400
transform 1 0 16688 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_145
timestamp 1669390400
transform 1 0 17584 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_149
timestamp 1669390400
transform 1 0 18032 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_151
timestamp 1669390400
transform 1 0 18256 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_154
timestamp 1669390400
transform 1 0 18592 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_161
timestamp 1669390400
transform 1 0 19376 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_168
timestamp 1669390400
transform 1 0 20160 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_172
timestamp 1669390400
transform 1 0 20608 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_182
timestamp 1669390400
transform 1 0 21728 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_198
timestamp 1669390400
transform 1 0 23520 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_206
timestamp 1669390400
transform 1 0 24416 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_209
timestamp 1669390400
transform 1 0 24752 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_217
timestamp 1669390400
transform 1 0 25648 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_227
timestamp 1669390400
transform 1 0 26768 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_235
timestamp 1669390400
transform 1 0 27664 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_257
timestamp 1669390400
transform 1 0 30128 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_261
timestamp 1669390400
transform 1 0 30576 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_265
timestamp 1669390400
transform 1 0 31024 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_267
timestamp 1669390400
transform 1 0 31248 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_276
timestamp 1669390400
transform 1 0 32256 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_286
timestamp 1669390400
transform 1 0 33376 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_293
timestamp 1669390400
transform 1 0 34160 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_305
timestamp 1669390400
transform 1 0 35504 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_315
timestamp 1669390400
transform 1 0 36624 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_324
timestamp 1669390400
transform 1 0 37632 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_328
timestamp 1669390400
transform 1 0 38080 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_332
timestamp 1669390400
transform 1 0 38528 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_336
timestamp 1669390400
transform 1 0 38976 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_345
timestamp 1669390400
transform 1 0 39984 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_353
timestamp 1669390400
transform 1 0 40880 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_357
timestamp 1669390400
transform 1 0 41328 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_361
timestamp 1669390400
transform 1 0 41776 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_373
timestamp 1669390400
transform 1 0 43120 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_377
timestamp 1669390400
transform 1 0 43568 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1669390400
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_395
timestamp 1669390400
transform 1 0 45584 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_399
timestamp 1669390400
transform 1 0 46032 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_401
timestamp 1669390400
transform 1 0 46256 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_410
timestamp 1669390400
transform 1 0 47264 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_414
timestamp 1669390400
transform 1 0 47712 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_456
timestamp 1669390400
transform 1 0 52416 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1669390400
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_463
timestamp 1669390400
transform 1 0 53200 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_474
timestamp 1669390400
transform 1 0 54432 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_476
timestamp 1669390400
transform 1 0 54656 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_493
timestamp 1669390400
transform 1 0 56560 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_497
timestamp 1669390400
transform 1 0 57008 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_501
timestamp 1669390400
transform 1 0 57456 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_505
timestamp 1669390400
transform 1 0 57904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1669390400
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_105
timestamp 1669390400
transform 1 0 13104 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_109
timestamp 1669390400
transform 1 0 13552 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_113
timestamp 1669390400
transform 1 0 14000 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_123
timestamp 1669390400
transform 1 0 15120 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_133
timestamp 1669390400
transform 1 0 16240 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_140
timestamp 1669390400
transform 1 0 17024 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_152
timestamp 1669390400
transform 1 0 18368 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_162
timestamp 1669390400
transform 1 0 19488 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_166
timestamp 1669390400
transform 1 0 19936 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_170
timestamp 1669390400
transform 1 0 20384 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_176
timestamp 1669390400
transform 1 0 21056 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_191
timestamp 1669390400
transform 1 0 22736 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_195
timestamp 1669390400
transform 1 0 23184 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_199
timestamp 1669390400
transform 1 0 23632 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_203
timestamp 1669390400
transform 1 0 24080 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_205
timestamp 1669390400
transform 1 0 24304 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1669390400
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_224
timestamp 1669390400
transform 1 0 26432 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_232
timestamp 1669390400
transform 1 0 27328 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_234
timestamp 1669390400
transform 1 0 27552 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_237
timestamp 1669390400
transform 1 0 27888 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_256
timestamp 1669390400
transform 1 0 30016 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_260
timestamp 1669390400
transform 1 0 30464 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_264
timestamp 1669390400
transform 1 0 30912 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_271
timestamp 1669390400
transform 1 0 31696 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_275
timestamp 1669390400
transform 1 0 32144 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_278
timestamp 1669390400
transform 1 0 32480 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_282
timestamp 1669390400
transform 1 0 32928 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_304
timestamp 1669390400
transform 1 0 35392 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_308
timestamp 1669390400
transform 1 0 35840 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_316
timestamp 1669390400
transform 1 0 36736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_322
timestamp 1669390400
transform 1 0 37408 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_326
timestamp 1669390400
transform 1 0 37856 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_334
timestamp 1669390400
transform 1 0 38752 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_346
timestamp 1669390400
transform 1 0 40096 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_353
timestamp 1669390400
transform 1 0 40880 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_359
timestamp 1669390400
transform 1 0 41552 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_365
timestamp 1669390400
transform 1 0 42224 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_369
timestamp 1669390400
transform 1 0 42672 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_373
timestamp 1669390400
transform 1 0 43120 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_382
timestamp 1669390400
transform 1 0 44128 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_386
timestamp 1669390400
transform 1 0 44576 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_390
timestamp 1669390400
transform 1 0 45024 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_394
timestamp 1669390400
transform 1 0 45472 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_398
timestamp 1669390400
transform 1 0 45920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_412
timestamp 1669390400
transform 1 0 47488 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_422
timestamp 1669390400
transform 1 0 48608 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_428
timestamp 1669390400
transform 1 0 49280 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_436
timestamp 1669390400
transform 1 0 50176 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_444
timestamp 1669390400
transform 1 0 51072 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_452
timestamp 1669390400
transform 1 0 51968 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_459
timestamp 1669390400
transform 1 0 52752 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_467
timestamp 1669390400
transform 1 0 53648 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_469
timestamp 1669390400
transform 1 0 53872 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_476
timestamp 1669390400
transform 1 0 54656 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_483
timestamp 1669390400
transform 1 0 55440 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_487
timestamp 1669390400
transform 1 0 55888 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_491
timestamp 1669390400
transform 1 0 56336 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_495
timestamp 1669390400
transform 1 0 56784 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_499
timestamp 1669390400
transform 1 0 57232 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_502
timestamp 1669390400
transform 1 0 57568 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_506
timestamp 1669390400
transform 1 0 58016 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_508
timestamp 1669390400
transform 1 0 58240 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1669390400
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1669390400
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_112
timestamp 1669390400
transform 1 0 13888 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_116
timestamp 1669390400
transform 1 0 14336 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_126
timestamp 1669390400
transform 1 0 15456 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_134
timestamp 1669390400
transform 1 0 16352 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_138
timestamp 1669390400
transform 1 0 16800 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_142
timestamp 1669390400
transform 1 0 17248 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_146
timestamp 1669390400
transform 1 0 17696 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_150
timestamp 1669390400
transform 1 0 18144 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_162
timestamp 1669390400
transform 1 0 19488 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_166
timestamp 1669390400
transform 1 0 19936 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1669390400
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_195
timestamp 1669390400
transform 1 0 23184 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_199
timestamp 1669390400
transform 1 0 23632 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_201
timestamp 1669390400
transform 1 0 23856 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_210
timestamp 1669390400
transform 1 0 24864 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_220
timestamp 1669390400
transform 1 0 25984 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_224
timestamp 1669390400
transform 1 0 26432 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_233
timestamp 1669390400
transform 1 0 27440 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_256
timestamp 1669390400
transform 1 0 30016 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_260
timestamp 1669390400
transform 1 0 30464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_277
timestamp 1669390400
transform 1 0 32368 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_287
timestamp 1669390400
transform 1 0 33488 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_291
timestamp 1669390400
transform 1 0 33936 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_299
timestamp 1669390400
transform 1 0 34832 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_301
timestamp 1669390400
transform 1 0 35056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_314
timestamp 1669390400
transform 1 0 36512 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_324
timestamp 1669390400
transform 1 0 37632 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_328
timestamp 1669390400
transform 1 0 38080 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_332
timestamp 1669390400
transform 1 0 38528 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_334
timestamp 1669390400
transform 1 0 38752 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_342
timestamp 1669390400
transform 1 0 39648 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_353
timestamp 1669390400
transform 1 0 40880 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_364
timestamp 1669390400
transform 1 0 42112 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_374
timestamp 1669390400
transform 1 0 43232 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_378
timestamp 1669390400
transform 1 0 43680 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_387
timestamp 1669390400
transform 1 0 44688 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1669390400
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_399
timestamp 1669390400
transform 1 0 46032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_403
timestamp 1669390400
transform 1 0 46480 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_410
timestamp 1669390400
transform 1 0 47264 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_418
timestamp 1669390400
transform 1 0 48160 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_422
timestamp 1669390400
transform 1 0 48608 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_426
timestamp 1669390400
transform 1 0 49056 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_430
timestamp 1669390400
transform 1 0 49504 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_434
timestamp 1669390400
transform 1 0 49952 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_441
timestamp 1669390400
transform 1 0 50736 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_449
timestamp 1669390400
transform 1 0 51632 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_453
timestamp 1669390400
transform 1 0 52080 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1669390400
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_463
timestamp 1669390400
transform 1 0 53200 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_477
timestamp 1669390400
transform 1 0 54768 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_486
timestamp 1669390400
transform 1 0 55776 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_494
timestamp 1669390400
transform 1 0 56672 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_502
timestamp 1669390400
transform 1 0 57568 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_508
timestamp 1669390400
transform 1 0 58240 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1669390400
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_105
timestamp 1669390400
transform 1 0 13104 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_109
timestamp 1669390400
transform 1 0 13552 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_134
timestamp 1669390400
transform 1 0 16352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_140
timestamp 1669390400
transform 1 0 17024 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_176
timestamp 1669390400
transform 1 0 21056 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_196
timestamp 1669390400
transform 1 0 23296 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_211
timestamp 1669390400
transform 1 0 24976 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_218
timestamp 1669390400
transform 1 0 25760 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_220
timestamp 1669390400
transform 1 0 25984 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_227
timestamp 1669390400
transform 1 0 26768 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_231
timestamp 1669390400
transform 1 0 27216 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_234
timestamp 1669390400
transform 1 0 27552 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_242
timestamp 1669390400
transform 1 0 28448 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_250
timestamp 1669390400
transform 1 0 29344 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_254
timestamp 1669390400
transform 1 0 29792 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_258
timestamp 1669390400
transform 1 0 30240 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_274
timestamp 1669390400
transform 1 0 32032 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_278
timestamp 1669390400
transform 1 0 32480 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_282
timestamp 1669390400
transform 1 0 32928 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_304
timestamp 1669390400
transform 1 0 35392 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_318
timestamp 1669390400
transform 1 0 36960 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_322
timestamp 1669390400
transform 1 0 37408 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_326
timestamp 1669390400
transform 1 0 37856 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_330
timestamp 1669390400
transform 1 0 38304 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_346
timestamp 1669390400
transform 1 0 40096 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_350
timestamp 1669390400
transform 1 0 40544 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_360
timestamp 1669390400
transform 1 0 41664 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_364
timestamp 1669390400
transform 1 0 42112 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_368
timestamp 1669390400
transform 1 0 42560 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_372
timestamp 1669390400
transform 1 0 43008 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_376
timestamp 1669390400
transform 1 0 43456 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_380
timestamp 1669390400
transform 1 0 43904 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_384
timestamp 1669390400
transform 1 0 44352 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_388
timestamp 1669390400
transform 1 0 44800 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_398
timestamp 1669390400
transform 1 0 45920 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_402
timestamp 1669390400
transform 1 0 46368 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_414
timestamp 1669390400
transform 1 0 47712 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_418
timestamp 1669390400
transform 1 0 48160 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_422
timestamp 1669390400
transform 1 0 48608 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_428
timestamp 1669390400
transform 1 0 49280 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_431
timestamp 1669390400
transform 1 0 49616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_452
timestamp 1669390400
transform 1 0 51968 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_456
timestamp 1669390400
transform 1 0 52416 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_464
timestamp 1669390400
transform 1 0 53312 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_473
timestamp 1669390400
transform 1 0 54320 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_481
timestamp 1669390400
transform 1 0 55216 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_483
timestamp 1669390400
transform 1 0 55440 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_488
timestamp 1669390400
transform 1 0 56000 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1669390400
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_499
timestamp 1669390400
transform 1 0 57232 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_506
timestamp 1669390400
transform 1 0 58016 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_508
timestamp 1669390400
transform 1 0 58240 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1669390400
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_116
timestamp 1669390400
transform 1 0 14336 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_123
timestamp 1669390400
transform 1 0 15120 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_137
timestamp 1669390400
transform 1 0 16688 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_143
timestamp 1669390400
transform 1 0 17360 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_151
timestamp 1669390400
transform 1 0 18256 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_155
timestamp 1669390400
transform 1 0 18704 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_164
timestamp 1669390400
transform 1 0 19712 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_168
timestamp 1669390400
transform 1 0 20160 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1669390400
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_182
timestamp 1669390400
transform 1 0 21728 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_186
timestamp 1669390400
transform 1 0 22176 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_196
timestamp 1669390400
transform 1 0 23296 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_213
timestamp 1669390400
transform 1 0 25200 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_217
timestamp 1669390400
transform 1 0 25648 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_221
timestamp 1669390400
transform 1 0 26096 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_224
timestamp 1669390400
transform 1 0 26432 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_228
timestamp 1669390400
transform 1 0 26880 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_232
timestamp 1669390400
transform 1 0 27328 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_236
timestamp 1669390400
transform 1 0 27776 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_243
timestamp 1669390400
transform 1 0 28560 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_253
timestamp 1669390400
transform 1 0 29680 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_257
timestamp 1669390400
transform 1 0 30128 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_265
timestamp 1669390400
transform 1 0 31024 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_267
timestamp 1669390400
transform 1 0 31248 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_276
timestamp 1669390400
transform 1 0 32256 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_283
timestamp 1669390400
transform 1 0 33040 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_287
timestamp 1669390400
transform 1 0 33488 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_291
timestamp 1669390400
transform 1 0 33936 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_295
timestamp 1669390400
transform 1 0 34384 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_299
timestamp 1669390400
transform 1 0 34832 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_303
timestamp 1669390400
transform 1 0 35280 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_307
timestamp 1669390400
transform 1 0 35728 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_311
timestamp 1669390400
transform 1 0 36176 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_323
timestamp 1669390400
transform 1 0 37520 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_330
timestamp 1669390400
transform 1 0 38304 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_355
timestamp 1669390400
transform 1 0 41104 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_359
timestamp 1669390400
transform 1 0 41552 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_366
timestamp 1669390400
transform 1 0 42336 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_378
timestamp 1669390400
transform 1 0 43680 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_386
timestamp 1669390400
transform 1 0 44576 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_395
timestamp 1669390400
transform 1 0 45584 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_405
timestamp 1669390400
transform 1 0 46704 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_412
timestamp 1669390400
transform 1 0 47488 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_416
timestamp 1669390400
transform 1 0 47936 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_418
timestamp 1669390400
transform 1 0 48160 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_424
timestamp 1669390400
transform 1 0 48832 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_428
timestamp 1669390400
transform 1 0 49280 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_430
timestamp 1669390400
transform 1 0 49504 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_442
timestamp 1669390400
transform 1 0 50848 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_446
timestamp 1669390400
transform 1 0 51296 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_450
timestamp 1669390400
transform 1 0 51744 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_454
timestamp 1669390400
transform 1 0 52192 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_458
timestamp 1669390400
transform 1 0 52640 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1669390400
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_463
timestamp 1669390400
transform 1 0 53200 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_466
timestamp 1669390400
transform 1 0 53536 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_470
timestamp 1669390400
transform 1 0 53984 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_472
timestamp 1669390400
transform 1 0 54208 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_479
timestamp 1669390400
transform 1 0 54992 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_489
timestamp 1669390400
transform 1 0 56112 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_497
timestamp 1669390400
transform 1 0 57008 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_505
timestamp 1669390400
transform 1 0 57904 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_6
timestamp 1669390400
transform 1 0 2016 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_14
timestamp 1669390400
transform 1 0 2912 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_18
timestamp 1669390400
transform 1 0 3360 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_50
timestamp 1669390400
transform 1 0 6944 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1669390400
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1669390400
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_105
timestamp 1669390400
transform 1 0 13104 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_121
timestamp 1669390400
transform 1 0 14896 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_160
timestamp 1669390400
transform 1 0 19264 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_164
timestamp 1669390400
transform 1 0 19712 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_222
timestamp 1669390400
transform 1 0 26208 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_226
timestamp 1669390400
transform 1 0 26656 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_230
timestamp 1669390400
transform 1 0 27104 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_236
timestamp 1669390400
transform 1 0 27776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_248
timestamp 1669390400
transform 1 0 29120 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_250
timestamp 1669390400
transform 1 0 29344 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_257
timestamp 1669390400
transform 1 0 30128 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_261
timestamp 1669390400
transform 1 0 30576 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_265
timestamp 1669390400
transform 1 0 31024 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_269
timestamp 1669390400
transform 1 0 31472 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_279
timestamp 1669390400
transform 1 0 32592 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1669390400
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_293
timestamp 1669390400
transform 1 0 34160 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_304
timestamp 1669390400
transform 1 0 35392 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_306
timestamp 1669390400
transform 1 0 35616 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_319
timestamp 1669390400
transform 1 0 37072 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_323
timestamp 1669390400
transform 1 0 37520 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_335
timestamp 1669390400
transform 1 0 38864 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_347
timestamp 1669390400
transform 1 0 40208 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_360
timestamp 1669390400
transform 1 0 41664 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_375
timestamp 1669390400
transform 1 0 43344 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_389
timestamp 1669390400
transform 1 0 44912 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_393
timestamp 1669390400
transform 1 0 45360 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_395
timestamp 1669390400
transform 1 0 45584 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_402
timestamp 1669390400
transform 1 0 46368 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_404
timestamp 1669390400
transform 1 0 46592 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_413
timestamp 1669390400
transform 1 0 47600 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1669390400
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_428
timestamp 1669390400
transform 1 0 49280 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_447
timestamp 1669390400
transform 1 0 51408 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_457
timestamp 1669390400
transform 1 0 52528 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_467
timestamp 1669390400
transform 1 0 53648 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_474
timestamp 1669390400
transform 1 0 54432 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_478
timestamp 1669390400
transform 1 0 54880 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_482
timestamp 1669390400
transform 1 0 55328 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1669390400
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_499
timestamp 1669390400
transform 1 0 57232 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_506
timestamp 1669390400
transform 1 0 58016 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_508
timestamp 1669390400
transform 1 0 58240 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_17
timestamp 1669390400
transform 1 0 3248 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_33
timestamp 1669390400
transform 1 0 5040 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1669390400
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_112
timestamp 1669390400
transform 1 0 13888 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_114
timestamp 1669390400
transform 1 0 14112 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_128
timestamp 1669390400
transform 1 0 15680 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_141
timestamp 1669390400
transform 1 0 17136 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_149
timestamp 1669390400
transform 1 0 18032 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_157
timestamp 1669390400
transform 1 0 18928 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_161
timestamp 1669390400
transform 1 0 19376 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_163
timestamp 1669390400
transform 1 0 19600 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_166
timestamp 1669390400
transform 1 0 19936 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_198
timestamp 1669390400
transform 1 0 23520 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_208
timestamp 1669390400
transform 1 0 24640 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_218
timestamp 1669390400
transform 1 0 25760 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_220
timestamp 1669390400
transform 1 0 25984 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_223
timestamp 1669390400
transform 1 0 26320 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_233
timestamp 1669390400
transform 1 0 27440 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_256
timestamp 1669390400
transform 1 0 30016 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_258
timestamp 1669390400
transform 1 0 30240 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_270
timestamp 1669390400
transform 1 0 31584 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_281
timestamp 1669390400
transform 1 0 32816 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_283
timestamp 1669390400
transform 1 0 33040 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_293
timestamp 1669390400
transform 1 0 34160 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_297
timestamp 1669390400
transform 1 0 34608 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_309
timestamp 1669390400
transform 1 0 35952 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_326
timestamp 1669390400
transform 1 0 37856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_330
timestamp 1669390400
transform 1 0 38304 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_341
timestamp 1669390400
transform 1 0 39536 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_349
timestamp 1669390400
transform 1 0 40432 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_374
timestamp 1669390400
transform 1 0 43232 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_378
timestamp 1669390400
transform 1 0 43680 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1669390400
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_394
timestamp 1669390400
transform 1 0 45472 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_435
timestamp 1669390400
transform 1 0 50064 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_439
timestamp 1669390400
transform 1 0 50512 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_449
timestamp 1669390400
transform 1 0 51632 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_453
timestamp 1669390400
transform 1 0 52080 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1669390400
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_463
timestamp 1669390400
transform 1 0 53200 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_470
timestamp 1669390400
transform 1 0 53984 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_474
timestamp 1669390400
transform 1 0 54432 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_476
timestamp 1669390400
transform 1 0 54656 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_491
timestamp 1669390400
transform 1 0 56336 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_503
timestamp 1669390400
transform 1 0 57680 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_507
timestamp 1669390400
transform 1 0 58128 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1669390400
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1669390400
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_105
timestamp 1669390400
transform 1 0 13104 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_121
timestamp 1669390400
transform 1 0 14896 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_125
timestamp 1669390400
transform 1 0 15344 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_127
timestamp 1669390400
transform 1 0 15568 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_148
timestamp 1669390400
transform 1 0 17920 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_173
timestamp 1669390400
transform 1 0 20720 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_187
timestamp 1669390400
transform 1 0 22288 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_189
timestamp 1669390400
transform 1 0 22512 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_192
timestamp 1669390400
transform 1 0 22848 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_200
timestamp 1669390400
transform 1 0 23744 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_208
timestamp 1669390400
transform 1 0 24640 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_221
timestamp 1669390400
transform 1 0 26096 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_231
timestamp 1669390400
transform 1 0 27216 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_241
timestamp 1669390400
transform 1 0 28336 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_247
timestamp 1669390400
transform 1 0 29008 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_251
timestamp 1669390400
transform 1 0 29456 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_255
timestamp 1669390400
transform 1 0 29904 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_257
timestamp 1669390400
transform 1 0 30128 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_260
timestamp 1669390400
transform 1 0 30464 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_264
timestamp 1669390400
transform 1 0 30912 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_266
timestamp 1669390400
transform 1 0 31136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_275
timestamp 1669390400
transform 1 0 32144 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_279
timestamp 1669390400
transform 1 0 32592 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_289
timestamp 1669390400
transform 1 0 33712 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_293
timestamp 1669390400
transform 1 0 34160 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_305
timestamp 1669390400
transform 1 0 35504 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_312
timestamp 1669390400
transform 1 0 36288 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_316
timestamp 1669390400
transform 1 0 36736 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_320
timestamp 1669390400
transform 1 0 37184 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_324
timestamp 1669390400
transform 1 0 37632 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_328
timestamp 1669390400
transform 1 0 38080 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_332
timestamp 1669390400
transform 1 0 38528 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_342
timestamp 1669390400
transform 1 0 39648 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_350
timestamp 1669390400
transform 1 0 40544 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_359
timestamp 1669390400
transform 1 0 41552 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_368
timestamp 1669390400
transform 1 0 42560 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_372
timestamp 1669390400
transform 1 0 43008 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_376
timestamp 1669390400
transform 1 0 43456 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_386
timestamp 1669390400
transform 1 0 44576 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_390
timestamp 1669390400
transform 1 0 45024 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_394
timestamp 1669390400
transform 1 0 45472 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_399
timestamp 1669390400
transform 1 0 46032 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_401
timestamp 1669390400
transform 1 0 46256 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_407
timestamp 1669390400
transform 1 0 46928 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_415
timestamp 1669390400
transform 1 0 47824 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1669390400
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_428
timestamp 1669390400
transform 1 0 49280 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_452
timestamp 1669390400
transform 1 0 51968 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_477
timestamp 1669390400
transform 1 0 54768 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1669390400
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_499
timestamp 1669390400
transform 1 0 57232 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_506
timestamp 1669390400
transform 1 0 58016 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_508
timestamp 1669390400
transform 1 0 58240 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1669390400
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1669390400
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_188
timestamp 1669390400
transform 1 0 22400 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_192
timestamp 1669390400
transform 1 0 22848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_196
timestamp 1669390400
transform 1 0 23296 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_199
timestamp 1669390400
transform 1 0 23632 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_213
timestamp 1669390400
transform 1 0 25200 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_223
timestamp 1669390400
transform 1 0 26320 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_227
timestamp 1669390400
transform 1 0 26768 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_233
timestamp 1669390400
transform 1 0 27440 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_241
timestamp 1669390400
transform 1 0 28336 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_243
timestamp 1669390400
transform 1 0 28560 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_246
timestamp 1669390400
transform 1 0 28896 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_254
timestamp 1669390400
transform 1 0 29792 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_262
timestamp 1669390400
transform 1 0 30688 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_265
timestamp 1669390400
transform 1 0 31024 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_275
timestamp 1669390400
transform 1 0 32144 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_279
timestamp 1669390400
transform 1 0 32592 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_283
timestamp 1669390400
transform 1 0 33040 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_290
timestamp 1669390400
transform 1 0 33824 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_294
timestamp 1669390400
transform 1 0 34272 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_301
timestamp 1669390400
transform 1 0 35056 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_308
timestamp 1669390400
transform 1 0 35840 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_312
timestamp 1669390400
transform 1 0 36288 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_316
timestamp 1669390400
transform 1 0 36736 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1669390400
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_325
timestamp 1669390400
transform 1 0 37744 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_332
timestamp 1669390400
transform 1 0 38528 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_339
timestamp 1669390400
transform 1 0 39312 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_343
timestamp 1669390400
transform 1 0 39760 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_347
timestamp 1669390400
transform 1 0 40208 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_357
timestamp 1669390400
transform 1 0 41328 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_361
timestamp 1669390400
transform 1 0 41776 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_365
timestamp 1669390400
transform 1 0 42224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_375
timestamp 1669390400
transform 1 0 43344 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_379
timestamp 1669390400
transform 1 0 43792 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_386
timestamp 1669390400
transform 1 0 44576 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_395
timestamp 1669390400
transform 1 0 45584 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_399
timestamp 1669390400
transform 1 0 46032 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_403
timestamp 1669390400
transform 1 0 46480 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_407
timestamp 1669390400
transform 1 0 46928 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_411
timestamp 1669390400
transform 1 0 47376 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_415
timestamp 1669390400
transform 1 0 47824 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_419
timestamp 1669390400
transform 1 0 48272 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_423
timestamp 1669390400
transform 1 0 48720 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_427
timestamp 1669390400
transform 1 0 49168 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_431
timestamp 1669390400
transform 1 0 49616 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_435
timestamp 1669390400
transform 1 0 50064 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_450
timestamp 1669390400
transform 1 0 51744 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_454
timestamp 1669390400
transform 1 0 52192 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_458
timestamp 1669390400
transform 1 0 52640 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1669390400
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_463
timestamp 1669390400
transform 1 0 53200 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_466
timestamp 1669390400
transform 1 0 53536 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_468
timestamp 1669390400
transform 1 0 53760 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_475
timestamp 1669390400
transform 1 0 54544 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_485
timestamp 1669390400
transform 1 0 55664 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_507
timestamp 1669390400
transform 1 0 58128 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1669390400
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1669390400
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_176
timestamp 1669390400
transform 1 0 21056 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_184
timestamp 1669390400
transform 1 0 21952 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_186
timestamp 1669390400
transform 1 0 22176 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_189
timestamp 1669390400
transform 1 0 22512 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_195
timestamp 1669390400
transform 1 0 23184 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_199
timestamp 1669390400
transform 1 0 23632 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_207
timestamp 1669390400
transform 1 0 24528 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_211
timestamp 1669390400
transform 1 0 24976 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_218
timestamp 1669390400
transform 1 0 25760 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_222
timestamp 1669390400
transform 1 0 26208 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_231
timestamp 1669390400
transform 1 0 27216 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_237
timestamp 1669390400
transform 1 0 27888 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_244
timestamp 1669390400
transform 1 0 28672 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_252
timestamp 1669390400
transform 1 0 29568 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_256
timestamp 1669390400
transform 1 0 30016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_268
timestamp 1669390400
transform 1 0 31360 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_276
timestamp 1669390400
transform 1 0 32256 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_280
timestamp 1669390400
transform 1 0 32704 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_296
timestamp 1669390400
transform 1 0 34496 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_306
timestamp 1669390400
transform 1 0 35616 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_310
timestamp 1669390400
transform 1 0 36064 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_314
timestamp 1669390400
transform 1 0 36512 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_324
timestamp 1669390400
transform 1 0 37632 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_338
timestamp 1669390400
transform 1 0 39200 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_342
timestamp 1669390400
transform 1 0 39648 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_346
timestamp 1669390400
transform 1 0 40096 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_350
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_360
timestamp 1669390400
transform 1 0 41664 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_368
timestamp 1669390400
transform 1 0 42560 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_376
timestamp 1669390400
transform 1 0 43456 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_378
timestamp 1669390400
transform 1 0 43680 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_386
timestamp 1669390400
transform 1 0 44576 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_388
timestamp 1669390400
transform 1 0 44800 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1669390400
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_428
timestamp 1669390400
transform 1 0 49280 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_431
timestamp 1669390400
transform 1 0 49616 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_435
timestamp 1669390400
transform 1 0 50064 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_437
timestamp 1669390400
transform 1 0 50288 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_448
timestamp 1669390400
transform 1 0 51520 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_458
timestamp 1669390400
transform 1 0 52640 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_466
timestamp 1669390400
transform 1 0 53536 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_470
timestamp 1669390400
transform 1 0 53984 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_489
timestamp 1669390400
transform 1 0 56112 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_493
timestamp 1669390400
transform 1 0 56560 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_499
timestamp 1669390400
transform 1 0 57232 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_506
timestamp 1669390400
transform 1 0 58016 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_508
timestamp 1669390400
transform 1 0 58240 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_6
timestamp 1669390400
transform 1 0 2016 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_14
timestamp 1669390400
transform 1 0 2912 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_18
timestamp 1669390400
transform 1 0 3360 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1669390400
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1669390400
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1669390400
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_193
timestamp 1669390400
transform 1 0 22960 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_195
timestamp 1669390400
transform 1 0 23184 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_198
timestamp 1669390400
transform 1 0 23520 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_205
timestamp 1669390400
transform 1 0 24304 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_213
timestamp 1669390400
transform 1 0 25200 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_221
timestamp 1669390400
transform 1 0 26096 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_235
timestamp 1669390400
transform 1 0 27664 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_246
timestamp 1669390400
transform 1 0 28896 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_252
timestamp 1669390400
transform 1 0 29568 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_259
timestamp 1669390400
transform 1 0 30352 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_269
timestamp 1669390400
transform 1 0 31472 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_277
timestamp 1669390400
transform 1 0 32368 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_281
timestamp 1669390400
transform 1 0 32816 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_285
timestamp 1669390400
transform 1 0 33264 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_289
timestamp 1669390400
transform 1 0 33712 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_302
timestamp 1669390400
transform 1 0 35168 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_314
timestamp 1669390400
transform 1 0 36512 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1669390400
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_337
timestamp 1669390400
transform 1 0 39088 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_341
timestamp 1669390400
transform 1 0 39536 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_345
timestamp 1669390400
transform 1 0 39984 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_349
timestamp 1669390400
transform 1 0 40432 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_351
timestamp 1669390400
transform 1 0 40656 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_360
timestamp 1669390400
transform 1 0 41664 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_364
timestamp 1669390400
transform 1 0 42112 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_373
timestamp 1669390400
transform 1 0 43120 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_385
timestamp 1669390400
transform 1 0 44464 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1669390400
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_395
timestamp 1669390400
transform 1 0 45584 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_399
timestamp 1669390400
transform 1 0 46032 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_410
timestamp 1669390400
transform 1 0 47264 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_418
timestamp 1669390400
transform 1 0 48160 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_432
timestamp 1669390400
transform 1 0 49728 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_444
timestamp 1669390400
transform 1 0 51072 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_448
timestamp 1669390400
transform 1 0 51520 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_452
timestamp 1669390400
transform 1 0 51968 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_456
timestamp 1669390400
transform 1 0 52416 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1669390400
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_463
timestamp 1669390400
transform 1 0 53200 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_474
timestamp 1669390400
transform 1 0 54432 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_478
timestamp 1669390400
transform 1 0 54880 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_506
timestamp 1669390400
transform 1 0 58016 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_508
timestamp 1669390400
transform 1 0 58240 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_66
timestamp 1669390400
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1669390400
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1669390400
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_176
timestamp 1669390400
transform 1 0 21056 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_180
timestamp 1669390400
transform 1 0 21504 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_193
timestamp 1669390400
transform 1 0 22960 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_203
timestamp 1669390400
transform 1 0 24080 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_207
timestamp 1669390400
transform 1 0 24528 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_211
timestamp 1669390400
transform 1 0 24976 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_219
timestamp 1669390400
transform 1 0 25872 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_223
timestamp 1669390400
transform 1 0 26320 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_241
timestamp 1669390400
transform 1 0 28336 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_245
timestamp 1669390400
transform 1 0 28784 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_253
timestamp 1669390400
transform 1 0 29680 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_257
timestamp 1669390400
transform 1 0 30128 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_259
timestamp 1669390400
transform 1 0 30352 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_265
timestamp 1669390400
transform 1 0 31024 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_277
timestamp 1669390400
transform 1 0 32368 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_281
timestamp 1669390400
transform 1 0 32816 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_295
timestamp 1669390400
transform 1 0 34384 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_299
timestamp 1669390400
transform 1 0 34832 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_307
timestamp 1669390400
transform 1 0 35728 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_311
timestamp 1669390400
transform 1 0 36176 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_315
timestamp 1669390400
transform 1 0 36624 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_322
timestamp 1669390400
transform 1 0 37408 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_332
timestamp 1669390400
transform 1 0 38528 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_336
timestamp 1669390400
transform 1 0 38976 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_344
timestamp 1669390400
transform 1 0 39872 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_367
timestamp 1669390400
transform 1 0 42448 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_371
timestamp 1669390400
transform 1 0 42896 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_373
timestamp 1669390400
transform 1 0 43120 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_379
timestamp 1669390400
transform 1 0 43792 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_383
timestamp 1669390400
transform 1 0 44240 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_387
timestamp 1669390400
transform 1 0 44688 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_394
timestamp 1669390400
transform 1 0 45472 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_413
timestamp 1669390400
transform 1 0 47600 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_421
timestamp 1669390400
transform 1 0 48496 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1669390400
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_428
timestamp 1669390400
transform 1 0 49280 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_437
timestamp 1669390400
transform 1 0 50288 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_445
timestamp 1669390400
transform 1 0 51184 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_449
timestamp 1669390400
transform 1 0 51632 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_453
timestamp 1669390400
transform 1 0 52080 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_457
timestamp 1669390400
transform 1 0 52528 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_461
timestamp 1669390400
transform 1 0 52976 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_465
timestamp 1669390400
transform 1 0 53424 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_469
timestamp 1669390400
transform 1 0 53872 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_473
timestamp 1669390400
transform 1 0 54320 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_481
timestamp 1669390400
transform 1 0 55216 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_491
timestamp 1669390400
transform 1 0 56336 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_495
timestamp 1669390400
transform 1 0 56784 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_499
timestamp 1669390400
transform 1 0 57232 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_506
timestamp 1669390400
transform 1 0 58016 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_508
timestamp 1669390400
transform 1 0 58240 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_17
timestamp 1669390400
transform 1 0 3248 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_33
timestamp 1669390400
transform 1 0 5040 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1669390400
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_140
timestamp 1669390400
transform 1 0 17024 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_148
timestamp 1669390400
transform 1 0 17920 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_152
timestamp 1669390400
transform 1 0 18368 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_160
timestamp 1669390400
transform 1 0 19264 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_24_166
timestamp 1669390400
transform 1 0 19936 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_174
timestamp 1669390400
transform 1 0 20832 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_183
timestamp 1669390400
transform 1 0 21840 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_190
timestamp 1669390400
transform 1 0 22624 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_192
timestamp 1669390400
transform 1 0 22848 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_198
timestamp 1669390400
transform 1 0 23520 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_202
timestamp 1669390400
transform 1 0 23968 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_206
timestamp 1669390400
transform 1 0 24416 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_210
timestamp 1669390400
transform 1 0 24864 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_214
timestamp 1669390400
transform 1 0 25312 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_224
timestamp 1669390400
transform 1 0 26432 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_228
timestamp 1669390400
transform 1 0 26880 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_236
timestamp 1669390400
transform 1 0 27776 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_240
timestamp 1669390400
transform 1 0 28224 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_244
timestamp 1669390400
transform 1 0 28672 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_257
timestamp 1669390400
transform 1 0 30128 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_261
timestamp 1669390400
transform 1 0 30576 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_264
timestamp 1669390400
transform 1 0 30912 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_266
timestamp 1669390400
transform 1 0 31136 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_273
timestamp 1669390400
transform 1 0 31920 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_277
timestamp 1669390400
transform 1 0 32368 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_281
timestamp 1669390400
transform 1 0 32816 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_283
timestamp 1669390400
transform 1 0 33040 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_286
timestamp 1669390400
transform 1 0 33376 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_296
timestamp 1669390400
transform 1 0 34496 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_300
timestamp 1669390400
transform 1 0 34944 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_304
timestamp 1669390400
transform 1 0 35392 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_308
timestamp 1669390400
transform 1 0 35840 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_312
timestamp 1669390400
transform 1 0 36288 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_316
timestamp 1669390400
transform 1 0 36736 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_323
timestamp 1669390400
transform 1 0 37520 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_331
timestamp 1669390400
transform 1 0 38416 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_340
timestamp 1669390400
transform 1 0 39424 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_342
timestamp 1669390400
transform 1 0 39648 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_351
timestamp 1669390400
transform 1 0 40656 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_358
timestamp 1669390400
transform 1 0 41440 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_362
timestamp 1669390400
transform 1 0 41888 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_366
timestamp 1669390400
transform 1 0 42336 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_370
timestamp 1669390400
transform 1 0 42784 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_374
timestamp 1669390400
transform 1 0 43232 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_378
timestamp 1669390400
transform 1 0 43680 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_386
timestamp 1669390400
transform 1 0 44576 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_395
timestamp 1669390400
transform 1 0 45584 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_397
timestamp 1669390400
transform 1 0 45808 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_403
timestamp 1669390400
transform 1 0 46480 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_415
timestamp 1669390400
transform 1 0 47824 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_428
timestamp 1669390400
transform 1 0 49280 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_432
timestamp 1669390400
transform 1 0 49728 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_436
timestamp 1669390400
transform 1 0 50176 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_440
timestamp 1669390400
transform 1 0 50624 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_444
timestamp 1669390400
transform 1 0 51072 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_448
timestamp 1669390400
transform 1 0 51520 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_452
timestamp 1669390400
transform 1 0 51968 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_454
timestamp 1669390400
transform 1 0 52192 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1669390400
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_463
timestamp 1669390400
transform 1 0 53200 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_474
timestamp 1669390400
transform 1 0 54432 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_482
timestamp 1669390400
transform 1 0 55328 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_486
timestamp 1669390400
transform 1 0 55776 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_490
timestamp 1669390400
transform 1 0 56224 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_499
timestamp 1669390400
transform 1 0 57232 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_507
timestamp 1669390400
transform 1 0 58128 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_66
timestamp 1669390400
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1669390400
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1669390400
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_150
timestamp 1669390400
transform 1 0 18144 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_164
timestamp 1669390400
transform 1 0 19712 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_170
timestamp 1669390400
transform 1 0 20384 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_174
timestamp 1669390400
transform 1 0 20832 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_201
timestamp 1669390400
transform 1 0 23856 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_205
timestamp 1669390400
transform 1 0 24304 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_228
timestamp 1669390400
transform 1 0 26880 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_235
timestamp 1669390400
transform 1 0 27664 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_252
timestamp 1669390400
transform 1 0 29568 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_262
timestamp 1669390400
transform 1 0 30688 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_270
timestamp 1669390400
transform 1 0 31584 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_274
timestamp 1669390400
transform 1 0 32032 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_276
timestamp 1669390400
transform 1 0 32256 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_279
timestamp 1669390400
transform 1 0 32592 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_289
timestamp 1669390400
transform 1 0 33712 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_293
timestamp 1669390400
transform 1 0 34160 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_295
timestamp 1669390400
transform 1 0 34384 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_304
timestamp 1669390400
transform 1 0 35392 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_312
timestamp 1669390400
transform 1 0 36288 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_316
timestamp 1669390400
transform 1 0 36736 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_320
timestamp 1669390400
transform 1 0 37184 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_324
timestamp 1669390400
transform 1 0 37632 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_328
timestamp 1669390400
transform 1 0 38080 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_332
timestamp 1669390400
transform 1 0 38528 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_336
timestamp 1669390400
transform 1 0 38976 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_340
timestamp 1669390400
transform 1 0 39424 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_343
timestamp 1669390400
transform 1 0 39760 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_360
timestamp 1669390400
transform 1 0 41664 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_364
timestamp 1669390400
transform 1 0 42112 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_372
timestamp 1669390400
transform 1 0 43008 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_376
timestamp 1669390400
transform 1 0 43456 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_380
timestamp 1669390400
transform 1 0 43904 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_384
timestamp 1669390400
transform 1 0 44352 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_388
timestamp 1669390400
transform 1 0 44800 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_392
timestamp 1669390400
transform 1 0 45248 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_396
timestamp 1669390400
transform 1 0 45696 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_400
timestamp 1669390400
transform 1 0 46144 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_404
timestamp 1669390400
transform 1 0 46592 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_408
timestamp 1669390400
transform 1 0 47040 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_412
timestamp 1669390400
transform 1 0 47488 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_416
timestamp 1669390400
transform 1 0 47936 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_420
timestamp 1669390400
transform 1 0 48384 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_424
timestamp 1669390400
transform 1 0 48832 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_428
timestamp 1669390400
transform 1 0 49280 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_437
timestamp 1669390400
transform 1 0 50288 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_441
timestamp 1669390400
transform 1 0 50736 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_445
timestamp 1669390400
transform 1 0 51184 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_447
timestamp 1669390400
transform 1 0 51408 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_456
timestamp 1669390400
transform 1 0 52416 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_476
timestamp 1669390400
transform 1 0 54656 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_486
timestamp 1669390400
transform 1 0 55776 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1669390400
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_499
timestamp 1669390400
transform 1 0 57232 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_508
timestamp 1669390400
transform 1 0 58240 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1669390400
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_140
timestamp 1669390400
transform 1 0 17024 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_186
timestamp 1669390400
transform 1 0 22176 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_190
timestamp 1669390400
transform 1 0 22624 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_200
timestamp 1669390400
transform 1 0 23744 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_227
timestamp 1669390400
transform 1 0 26768 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_235
timestamp 1669390400
transform 1 0 27664 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_239
timestamp 1669390400
transform 1 0 28112 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_243
timestamp 1669390400
transform 1 0 28560 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_259
timestamp 1669390400
transform 1 0 30352 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_263
timestamp 1669390400
transform 1 0 30800 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_267
timestamp 1669390400
transform 1 0 31248 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_286
timestamp 1669390400
transform 1 0 33376 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_290
timestamp 1669390400
transform 1 0 33824 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_295
timestamp 1669390400
transform 1 0 34384 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_306
timestamp 1669390400
transform 1 0 35616 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_314
timestamp 1669390400
transform 1 0 36512 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_328
timestamp 1669390400
transform 1 0 38080 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_341
timestamp 1669390400
transform 1 0 39536 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_351
timestamp 1669390400
transform 1 0 40656 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_358
timestamp 1669390400
transform 1 0 41440 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_360
timestamp 1669390400
transform 1 0 41664 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_371
timestamp 1669390400
transform 1 0 42896 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_375
timestamp 1669390400
transform 1 0 43344 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_386
timestamp 1669390400
transform 1 0 44576 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_395
timestamp 1669390400
transform 1 0 45584 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_399
timestamp 1669390400
transform 1 0 46032 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_411
timestamp 1669390400
transform 1 0 47376 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_415
timestamp 1669390400
transform 1 0 47824 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_419
timestamp 1669390400
transform 1 0 48272 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_421
timestamp 1669390400
transform 1 0 48496 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_427
timestamp 1669390400
transform 1 0 49168 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_435
timestamp 1669390400
transform 1 0 50064 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_445
timestamp 1669390400
transform 1 0 51184 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1669390400
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_463
timestamp 1669390400
transform 1 0 53200 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_472
timestamp 1669390400
transform 1 0 54208 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_476
timestamp 1669390400
transform 1 0 54656 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_491
timestamp 1669390400
transform 1 0 56336 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_503
timestamp 1669390400
transform 1 0 57680 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_507
timestamp 1669390400
transform 1 0 58128 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1669390400
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1669390400
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_105
timestamp 1669390400
transform 1 0 13104 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_113
timestamp 1669390400
transform 1 0 14000 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_121
timestamp 1669390400
transform 1 0 14896 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_125
timestamp 1669390400
transform 1 0 15344 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_148
timestamp 1669390400
transform 1 0 17920 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_150
timestamp 1669390400
transform 1 0 18144 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_176
timestamp 1669390400
transform 1 0 21056 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_180
timestamp 1669390400
transform 1 0 21504 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_182
timestamp 1669390400
transform 1 0 21728 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_185
timestamp 1669390400
transform 1 0 22064 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_209
timestamp 1669390400
transform 1 0 24752 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_224
timestamp 1669390400
transform 1 0 26432 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_231
timestamp 1669390400
transform 1 0 27216 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_235
timestamp 1669390400
transform 1 0 27664 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_239
timestamp 1669390400
transform 1 0 28112 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_247
timestamp 1669390400
transform 1 0 29008 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_256
timestamp 1669390400
transform 1 0 30016 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_260
timestamp 1669390400
transform 1 0 30464 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_262
timestamp 1669390400
transform 1 0 30688 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_265
timestamp 1669390400
transform 1 0 31024 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_269
timestamp 1669390400
transform 1 0 31472 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_282
timestamp 1669390400
transform 1 0 32928 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_297
timestamp 1669390400
transform 1 0 34608 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_311
timestamp 1669390400
transform 1 0 36176 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_319
timestamp 1669390400
transform 1 0 37072 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_323
timestamp 1669390400
transform 1 0 37520 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_327
timestamp 1669390400
transform 1 0 37968 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_331
timestamp 1669390400
transform 1 0 38416 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_335
timestamp 1669390400
transform 1 0 38864 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_348
timestamp 1669390400
transform 1 0 40320 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_352
timestamp 1669390400
transform 1 0 40768 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_360
timestamp 1669390400
transform 1 0 41664 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_362
timestamp 1669390400
transform 1 0 41888 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_374
timestamp 1669390400
transform 1 0 43232 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_376
timestamp 1669390400
transform 1 0 43456 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_386
timestamp 1669390400
transform 1 0 44576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_390
timestamp 1669390400
transform 1 0 45024 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_401
timestamp 1669390400
transform 1 0 46256 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_415
timestamp 1669390400
transform 1 0 47824 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_419
timestamp 1669390400
transform 1 0 48272 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_423
timestamp 1669390400
transform 1 0 48720 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1669390400
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_428
timestamp 1669390400
transform 1 0 49280 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_438
timestamp 1669390400
transform 1 0 50400 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_446
timestamp 1669390400
transform 1 0 51296 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_453
timestamp 1669390400
transform 1 0 52080 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_457
timestamp 1669390400
transform 1 0 52528 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_461
timestamp 1669390400
transform 1 0 52976 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_465
timestamp 1669390400
transform 1 0 53424 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_467
timestamp 1669390400
transform 1 0 53648 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_474
timestamp 1669390400
transform 1 0 54432 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_482
timestamp 1669390400
transform 1 0 55328 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_484
timestamp 1669390400
transform 1 0 55552 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1669390400
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_499
timestamp 1669390400
transform 1 0 57232 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_508
timestamp 1669390400
transform 1 0 58240 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1669390400
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1669390400
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1669390400
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_112
timestamp 1669390400
transform 1 0 13888 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_114
timestamp 1669390400
transform 1 0 14112 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_121
timestamp 1669390400
transform 1 0 14896 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_129
timestamp 1669390400
transform 1 0 15792 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_133
timestamp 1669390400
transform 1 0 16240 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_141
timestamp 1669390400
transform 1 0 17136 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_182
timestamp 1669390400
transform 1 0 21728 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_198
timestamp 1669390400
transform 1 0 23520 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_204
timestamp 1669390400
transform 1 0 24192 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_222
timestamp 1669390400
transform 1 0 26208 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_226
timestamp 1669390400
transform 1 0 26656 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_228
timestamp 1669390400
transform 1 0 26880 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_231
timestamp 1669390400
transform 1 0 27216 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_241
timestamp 1669390400
transform 1 0 28336 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_245
timestamp 1669390400
transform 1 0 28784 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_254
timestamp 1669390400
transform 1 0 29792 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_258
timestamp 1669390400
transform 1 0 30240 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_274
timestamp 1669390400
transform 1 0 32032 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_286
timestamp 1669390400
transform 1 0 33376 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_296
timestamp 1669390400
transform 1 0 34496 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_310
timestamp 1669390400
transform 1 0 36064 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_333
timestamp 1669390400
transform 1 0 38640 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_343
timestamp 1669390400
transform 1 0 39760 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_345
timestamp 1669390400
transform 1 0 39984 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_352
timestamp 1669390400
transform 1 0 40768 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_359
timestamp 1669390400
transform 1 0 41552 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_363
timestamp 1669390400
transform 1 0 42000 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_367
timestamp 1669390400
transform 1 0 42448 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_377
timestamp 1669390400
transform 1 0 43568 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_387
timestamp 1669390400
transform 1 0 44688 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1669390400
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_402
timestamp 1669390400
transform 1 0 46368 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_408
timestamp 1669390400
transform 1 0 47040 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_420
timestamp 1669390400
transform 1 0 48384 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_424
timestamp 1669390400
transform 1 0 48832 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_428
timestamp 1669390400
transform 1 0 49280 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_432
timestamp 1669390400
transform 1 0 49728 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_440
timestamp 1669390400
transform 1 0 50624 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_444
timestamp 1669390400
transform 1 0 51072 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_448
timestamp 1669390400
transform 1 0 51520 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_452
timestamp 1669390400
transform 1 0 51968 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_456
timestamp 1669390400
transform 1 0 52416 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1669390400
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_463
timestamp 1669390400
transform 1 0 53200 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_470
timestamp 1669390400
transform 1 0 53984 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_474
timestamp 1669390400
transform 1 0 54432 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_478
timestamp 1669390400
transform 1 0 54880 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_482
timestamp 1669390400
transform 1 0 55328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_486
timestamp 1669390400
transform 1 0 55776 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_499
timestamp 1669390400
transform 1 0 57232 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_507
timestamp 1669390400
transform 1 0 58128 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1669390400
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_105
timestamp 1669390400
transform 1 0 13104 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_154
timestamp 1669390400
transform 1 0 18592 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_168
timestamp 1669390400
transform 1 0 20160 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_172
timestamp 1669390400
transform 1 0 20608 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_176
timestamp 1669390400
transform 1 0 21056 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_218
timestamp 1669390400
transform 1 0 25760 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_226
timestamp 1669390400
transform 1 0 26656 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_262
timestamp 1669390400
transform 1 0 30688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_266
timestamp 1669390400
transform 1 0 31136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_280
timestamp 1669390400
transform 1 0 32704 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_289
timestamp 1669390400
transform 1 0 33712 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_293
timestamp 1669390400
transform 1 0 34160 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_300
timestamp 1669390400
transform 1 0 34944 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_307
timestamp 1669390400
transform 1 0 35728 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_311
timestamp 1669390400
transform 1 0 36176 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_313
timestamp 1669390400
transform 1 0 36400 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_321
timestamp 1669390400
transform 1 0 37296 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_329
timestamp 1669390400
transform 1 0 38192 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_333
timestamp 1669390400
transform 1 0 38640 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_337
timestamp 1669390400
transform 1 0 39088 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_341
timestamp 1669390400
transform 1 0 39536 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_345
timestamp 1669390400
transform 1 0 39984 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_349
timestamp 1669390400
transform 1 0 40432 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_353
timestamp 1669390400
transform 1 0 40880 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_360
timestamp 1669390400
transform 1 0 41664 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_366
timestamp 1669390400
transform 1 0 42336 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_370
timestamp 1669390400
transform 1 0 42784 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_374
timestamp 1669390400
transform 1 0 43232 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_377
timestamp 1669390400
transform 1 0 43568 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_402
timestamp 1669390400
transform 1 0 46368 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_406
timestamp 1669390400
transform 1 0 46816 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_410
timestamp 1669390400
transform 1 0 47264 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_414
timestamp 1669390400
transform 1 0 47712 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1669390400
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_428
timestamp 1669390400
transform 1 0 49280 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_431
timestamp 1669390400
transform 1 0 49616 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_435
timestamp 1669390400
transform 1 0 50064 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_445
timestamp 1669390400
transform 1 0 51184 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_455
timestamp 1669390400
transform 1 0 52304 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_457
timestamp 1669390400
transform 1 0 52528 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_472
timestamp 1669390400
transform 1 0 54208 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_476
timestamp 1669390400
transform 1 0 54656 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_480
timestamp 1669390400
transform 1 0 55104 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_484
timestamp 1669390400
transform 1 0 55552 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_486
timestamp 1669390400
transform 1 0 55776 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_493
timestamp 1669390400
transform 1 0 56560 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_499
timestamp 1669390400
transform 1 0 57232 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_502
timestamp 1669390400
transform 1 0 57568 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_506
timestamp 1669390400
transform 1 0 58016 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_508
timestamp 1669390400
transform 1 0 58240 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_8
timestamp 1669390400
transform 1 0 2240 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_24
timestamp 1669390400
transform 1 0 4032 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_32
timestamp 1669390400
transform 1 0 4928 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1669390400
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_69
timestamp 1669390400
transform 1 0 9072 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_91
timestamp 1669390400
transform 1 0 11536 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_99
timestamp 1669390400
transform 1 0 12432 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_125
timestamp 1669390400
transform 1 0 15344 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_143
timestamp 1669390400
transform 1 0 17360 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_151
timestamp 1669390400
transform 1 0 18256 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_155
timestamp 1669390400
transform 1 0 18704 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_171
timestamp 1669390400
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_175
timestamp 1669390400
transform 1 0 20944 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_186
timestamp 1669390400
transform 1 0 22176 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_202
timestamp 1669390400
transform 1 0 23968 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_212
timestamp 1669390400
transform 1 0 25088 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_219
timestamp 1669390400
transform 1 0 25872 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_223
timestamp 1669390400
transform 1 0 26320 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_227
timestamp 1669390400
transform 1 0 26768 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_235
timestamp 1669390400
transform 1 0 27664 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_241
timestamp 1669390400
transform 1 0 28336 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_245
timestamp 1669390400
transform 1 0 28784 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_254
timestamp 1669390400
transform 1 0 29792 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_257
timestamp 1669390400
transform 1 0 30128 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_261
timestamp 1669390400
transform 1 0 30576 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_263
timestamp 1669390400
transform 1 0 30800 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_266
timestamp 1669390400
transform 1 0 31136 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_270
timestamp 1669390400
transform 1 0 31584 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_276
timestamp 1669390400
transform 1 0 32256 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_282
timestamp 1669390400
transform 1 0 32928 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_286
timestamp 1669390400
transform 1 0 33376 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_310
timestamp 1669390400
transform 1 0 36064 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_314
timestamp 1669390400
transform 1 0 36512 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_330
timestamp 1669390400
transform 1 0 38304 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_340
timestamp 1669390400
transform 1 0 39424 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_344
timestamp 1669390400
transform 1 0 39872 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_348
timestamp 1669390400
transform 1 0 40320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_354
timestamp 1669390400
transform 1 0 40992 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_364
timestamp 1669390400
transform 1 0 42112 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_371
timestamp 1669390400
transform 1 0 42896 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_375
timestamp 1669390400
transform 1 0 43344 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_379
timestamp 1669390400
transform 1 0 43792 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_383
timestamp 1669390400
transform 1 0 44240 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_387
timestamp 1669390400
transform 1 0 44688 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1669390400
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_401
timestamp 1669390400
transform 1 0 46256 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_411
timestamp 1669390400
transform 1 0 47376 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_432
timestamp 1669390400
transform 1 0 49728 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_443
timestamp 1669390400
transform 1 0 50960 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_451
timestamp 1669390400
transform 1 0 51856 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_453
timestamp 1669390400
transform 1 0 52080 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1669390400
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_463
timestamp 1669390400
transform 1 0 53200 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_470
timestamp 1669390400
transform 1 0 53984 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_478
timestamp 1669390400
transform 1 0 54880 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_486
timestamp 1669390400
transform 1 0 55776 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_488
timestamp 1669390400
transform 1 0 56000 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_497
timestamp 1669390400
transform 1 0 57008 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_505
timestamp 1669390400
transform 1 0 57904 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_17
timestamp 1669390400
transform 1 0 3248 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_21
timestamp 1669390400
transform 1 0 3696 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_25
timestamp 1669390400
transform 1 0 4144 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_57
timestamp 1669390400
transform 1 0 7728 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_65
timestamp 1669390400
transform 1 0 8624 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_69
timestamp 1669390400
transform 1 0 9072 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_77
timestamp 1669390400
transform 1 0 9968 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_115
timestamp 1669390400
transform 1 0 14224 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_123
timestamp 1669390400
transform 1 0 15120 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_127
timestamp 1669390400
transform 1 0 15568 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_131
timestamp 1669390400
transform 1 0 16016 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_135
timestamp 1669390400
transform 1 0 16464 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_153
timestamp 1669390400
transform 1 0 18480 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_161
timestamp 1669390400
transform 1 0 19376 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_169
timestamp 1669390400
transform 1 0 20272 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_173
timestamp 1669390400
transform 1 0 20720 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_175
timestamp 1669390400
transform 1 0 20944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_210
timestamp 1669390400
transform 1 0 24864 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_224
timestamp 1669390400
transform 1 0 26432 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_228
timestamp 1669390400
transform 1 0 26880 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_236
timestamp 1669390400
transform 1 0 27776 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_244
timestamp 1669390400
transform 1 0 28672 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_248
timestamp 1669390400
transform 1 0 29120 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_255
timestamp 1669390400
transform 1 0 29904 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_273
timestamp 1669390400
transform 1 0 31920 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_277
timestamp 1669390400
transform 1 0 32368 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_280
timestamp 1669390400
transform 1 0 32704 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_293
timestamp 1669390400
transform 1 0 34160 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_295
timestamp 1669390400
transform 1 0 34384 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_304
timestamp 1669390400
transform 1 0 35392 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_312
timestamp 1669390400
transform 1 0 36288 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_316
timestamp 1669390400
transform 1 0 36736 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_320
timestamp 1669390400
transform 1 0 37184 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_324
timestamp 1669390400
transform 1 0 37632 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_326
timestamp 1669390400
transform 1 0 37856 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_333
timestamp 1669390400
transform 1 0 38640 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_337
timestamp 1669390400
transform 1 0 39088 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_347
timestamp 1669390400
transform 1 0 40208 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_364
timestamp 1669390400
transform 1 0 42112 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_376
timestamp 1669390400
transform 1 0 43456 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_386
timestamp 1669390400
transform 1 0 44576 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_403
timestamp 1669390400
transform 1 0 46480 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_410
timestamp 1669390400
transform 1 0 47264 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_420
timestamp 1669390400
transform 1 0 48384 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_424
timestamp 1669390400
transform 1 0 48832 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_428
timestamp 1669390400
transform 1 0 49280 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_434
timestamp 1669390400
transform 1 0 49952 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_438
timestamp 1669390400
transform 1 0 50400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_442
timestamp 1669390400
transform 1 0 50848 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_453
timestamp 1669390400
transform 1 0 52080 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_457
timestamp 1669390400
transform 1 0 52528 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_459
timestamp 1669390400
transform 1 0 52752 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_466
timestamp 1669390400
transform 1 0 53536 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_470
timestamp 1669390400
transform 1 0 53984 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_474
timestamp 1669390400
transform 1 0 54432 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_478
timestamp 1669390400
transform 1 0 54880 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_488
timestamp 1669390400
transform 1 0 56000 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1669390400
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_499
timestamp 1669390400
transform 1 0 57232 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_502
timestamp 1669390400
transform 1 0 57568 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_506
timestamp 1669390400
transform 1 0 58016 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_508
timestamp 1669390400
transform 1 0 58240 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_8
timestamp 1669390400
transform 1 0 2240 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_12
timestamp 1669390400
transform 1 0 2688 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_16
timestamp 1669390400
transform 1 0 3136 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_18
timestamp 1669390400
transform 1 0 3360 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_21
timestamp 1669390400
transform 1 0 3696 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_25
timestamp 1669390400
transform 1 0 4144 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_29
timestamp 1669390400
transform 1 0 4592 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_33
timestamp 1669390400
transform 1 0 5040 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1669390400
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_110
timestamp 1669390400
transform 1 0 13664 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_147
timestamp 1669390400
transform 1 0 17808 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_151
timestamp 1669390400
transform 1 0 18256 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_159
timestamp 1669390400
transform 1 0 19152 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_163
timestamp 1669390400
transform 1 0 19600 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_165
timestamp 1669390400
transform 1 0 19824 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_168
timestamp 1669390400
transform 1 0 20160 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_187
timestamp 1669390400
transform 1 0 22288 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_190
timestamp 1669390400
transform 1 0 22624 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_206
timestamp 1669390400
transform 1 0 24416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_210
timestamp 1669390400
transform 1 0 24864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_217
timestamp 1669390400
transform 1 0 25648 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_221
timestamp 1669390400
transform 1 0 26096 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_223
timestamp 1669390400
transform 1 0 26320 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_226
timestamp 1669390400
transform 1 0 26656 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_234
timestamp 1669390400
transform 1 0 27552 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_242
timestamp 1669390400
transform 1 0 28448 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_244
timestamp 1669390400
transform 1 0 28672 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_252
timestamp 1669390400
transform 1 0 29568 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_255
timestamp 1669390400
transform 1 0 29904 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_269
timestamp 1669390400
transform 1 0 31472 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_278
timestamp 1669390400
transform 1 0 32480 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_282
timestamp 1669390400
transform 1 0 32928 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_284
timestamp 1669390400
transform 1 0 33152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_291
timestamp 1669390400
transform 1 0 33936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_295
timestamp 1669390400
transform 1 0 34384 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_304
timestamp 1669390400
transform 1 0 35392 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_308
timestamp 1669390400
transform 1 0 35840 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_312
timestamp 1669390400
transform 1 0 36288 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_316
timestamp 1669390400
transform 1 0 36736 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1669390400
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_327
timestamp 1669390400
transform 1 0 37968 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_331
timestamp 1669390400
transform 1 0 38416 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_349
timestamp 1669390400
transform 1 0 40432 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_353
timestamp 1669390400
transform 1 0 40880 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_360
timestamp 1669390400
transform 1 0 41664 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_364
timestamp 1669390400
transform 1 0 42112 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_373
timestamp 1669390400
transform 1 0 43120 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_381
timestamp 1669390400
transform 1 0 44016 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1669390400
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_398
timestamp 1669390400
transform 1 0 45920 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_402
timestamp 1669390400
transform 1 0 46368 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_406
timestamp 1669390400
transform 1 0 46816 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_410
timestamp 1669390400
transform 1 0 47264 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_414
timestamp 1669390400
transform 1 0 47712 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_418
timestamp 1669390400
transform 1 0 48160 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_425
timestamp 1669390400
transform 1 0 48944 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_429
timestamp 1669390400
transform 1 0 49392 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_435
timestamp 1669390400
transform 1 0 50064 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_439
timestamp 1669390400
transform 1 0 50512 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_443
timestamp 1669390400
transform 1 0 50960 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_451
timestamp 1669390400
transform 1 0 51856 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_455
timestamp 1669390400
transform 1 0 52304 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_459
timestamp 1669390400
transform 1 0 52752 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_463
timestamp 1669390400
transform 1 0 53200 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_472
timestamp 1669390400
transform 1 0 54208 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_476
timestamp 1669390400
transform 1 0 54656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_480
timestamp 1669390400
transform 1 0 55104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_487
timestamp 1669390400
transform 1 0 55888 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_489
timestamp 1669390400
transform 1 0 56112 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_496
timestamp 1669390400
transform 1 0 56896 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_504
timestamp 1669390400
transform 1 0 57792 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_508
timestamp 1669390400
transform 1 0 58240 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_6
timestamp 1669390400
transform 1 0 2016 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_10
timestamp 1669390400
transform 1 0 2464 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_14
timestamp 1669390400
transform 1 0 2912 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_16
timestamp 1669390400
transform 1 0 3136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_19
timestamp 1669390400
transform 1 0 3472 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_23
timestamp 1669390400
transform 1 0 3920 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_27
timestamp 1669390400
transform 1 0 4368 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_31
timestamp 1669390400
transform 1 0 4816 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_33
timestamp 1669390400
transform 1 0 5040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_36
timestamp 1669390400
transform 1 0 5376 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_40
timestamp 1669390400
transform 1 0 5824 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_44
timestamp 1669390400
transform 1 0 6272 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_48
timestamp 1669390400
transform 1 0 6720 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_50
timestamp 1669390400
transform 1 0 6944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_53
timestamp 1669390400
transform 1 0 7280 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_57
timestamp 1669390400
transform 1 0 7728 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_63
timestamp 1669390400
transform 1 0 8400 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_67
timestamp 1669390400
transform 1 0 8848 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_76
timestamp 1669390400
transform 1 0 9856 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_82
timestamp 1669390400
transform 1 0 10528 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_96
timestamp 1669390400
transform 1 0 12096 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_104
timestamp 1669390400
transform 1 0 12992 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_108
timestamp 1669390400
transform 1 0 13440 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_122
timestamp 1669390400
transform 1 0 15008 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_130
timestamp 1669390400
transform 1 0 15904 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_134
timestamp 1669390400
transform 1 0 16352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_138
timestamp 1669390400
transform 1 0 16800 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_147
timestamp 1669390400
transform 1 0 17808 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_149
timestamp 1669390400
transform 1 0 18032 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_152
timestamp 1669390400
transform 1 0 18368 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_188
timestamp 1669390400
transform 1 0 22400 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_192
timestamp 1669390400
transform 1 0 22848 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_200
timestamp 1669390400
transform 1 0 23744 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_204
timestamp 1669390400
transform 1 0 24192 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_208
timestamp 1669390400
transform 1 0 24640 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_250
timestamp 1669390400
transform 1 0 29344 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_254
timestamp 1669390400
transform 1 0 29792 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_257
timestamp 1669390400
transform 1 0 30128 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_265
timestamp 1669390400
transform 1 0 31024 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_267
timestamp 1669390400
transform 1 0 31248 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_280
timestamp 1669390400
transform 1 0 32704 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_289
timestamp 1669390400
transform 1 0 33712 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_293
timestamp 1669390400
transform 1 0 34160 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_297
timestamp 1669390400
transform 1 0 34608 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_307
timestamp 1669390400
transform 1 0 35728 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_311
timestamp 1669390400
transform 1 0 36176 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_317
timestamp 1669390400
transform 1 0 36848 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_327
timestamp 1669390400
transform 1 0 37968 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_335
timestamp 1669390400
transform 1 0 38864 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_339
timestamp 1669390400
transform 1 0 39312 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_364
timestamp 1669390400
transform 1 0 42112 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_368
timestamp 1669390400
transform 1 0 42560 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_376
timestamp 1669390400
transform 1 0 43456 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_380
timestamp 1669390400
transform 1 0 43904 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_382
timestamp 1669390400
transform 1 0 44128 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_390
timestamp 1669390400
transform 1 0 45024 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_392
timestamp 1669390400
transform 1 0 45248 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_406
timestamp 1669390400
transform 1 0 46816 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_416
timestamp 1669390400
transform 1 0 47936 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_420
timestamp 1669390400
transform 1 0 48384 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_422
timestamp 1669390400
transform 1 0 48608 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1669390400
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_428
timestamp 1669390400
transform 1 0 49280 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_434
timestamp 1669390400
transform 1 0 49952 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_442
timestamp 1669390400
transform 1 0 50848 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_451
timestamp 1669390400
transform 1 0 51856 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_455
timestamp 1669390400
transform 1 0 52304 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_459
timestamp 1669390400
transform 1 0 52752 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_463
timestamp 1669390400
transform 1 0 53200 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_465
timestamp 1669390400
transform 1 0 53424 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_468
timestamp 1669390400
transform 1 0 53760 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_475
timestamp 1669390400
transform 1 0 54544 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_491
timestamp 1669390400
transform 1 0 56336 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_493
timestamp 1669390400
transform 1 0 56560 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1669390400
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_499
timestamp 1669390400
transform 1 0 57232 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_506
timestamp 1669390400
transform 1 0 58016 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_508
timestamp 1669390400
transform 1 0 58240 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_6
timestamp 1669390400
transform 1 0 2016 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_14
timestamp 1669390400
transform 1 0 2912 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_18
timestamp 1669390400
transform 1 0 3360 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_22
timestamp 1669390400
transform 1 0 3808 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_24
timestamp 1669390400
transform 1 0 4032 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_27
timestamp 1669390400
transform 1 0 4368 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_31
timestamp 1669390400
transform 1 0 4816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_40
timestamp 1669390400
transform 1 0 5824 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_44
timestamp 1669390400
transform 1 0 6272 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_47
timestamp 1669390400
transform 1 0 6608 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_49
timestamp 1669390400
transform 1 0 6832 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_63
timestamp 1669390400
transform 1 0 8400 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_71
timestamp 1669390400
transform 1 0 9296 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_73
timestamp 1669390400
transform 1 0 9520 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_76
timestamp 1669390400
transform 1 0 9856 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_84
timestamp 1669390400
transform 1 0 10752 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_92
timestamp 1669390400
transform 1 0 11648 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_96
timestamp 1669390400
transform 1 0 12096 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_100
timestamp 1669390400
transform 1 0 12544 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_104
timestamp 1669390400
transform 1 0 12992 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_112
timestamp 1669390400
transform 1 0 13888 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_114
timestamp 1669390400
transform 1 0 14112 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_123
timestamp 1669390400
transform 1 0 15120 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_143
timestamp 1669390400
transform 1 0 17360 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_151
timestamp 1669390400
transform 1 0 18256 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_166
timestamp 1669390400
transform 1 0 19936 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_173
timestamp 1669390400
transform 1 0 20720 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_182
timestamp 1669390400
transform 1 0 21728 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_186
timestamp 1669390400
transform 1 0 22176 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_190
timestamp 1669390400
transform 1 0 22624 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_194
timestamp 1669390400
transform 1 0 23072 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_230
timestamp 1669390400
transform 1 0 27104 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_234
timestamp 1669390400
transform 1 0 27552 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_242
timestamp 1669390400
transform 1 0 28448 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_246
timestamp 1669390400
transform 1 0 28896 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_256
timestamp 1669390400
transform 1 0 30016 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_260
timestamp 1669390400
transform 1 0 30464 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_264
timestamp 1669390400
transform 1 0 30912 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_268
timestamp 1669390400
transform 1 0 31360 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_272
timestamp 1669390400
transform 1 0 31808 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_278
timestamp 1669390400
transform 1 0 32480 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_286
timestamp 1669390400
transform 1 0 33376 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_294
timestamp 1669390400
transform 1 0 34272 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_298
timestamp 1669390400
transform 1 0 34720 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_305
timestamp 1669390400
transform 1 0 35504 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_324
timestamp 1669390400
transform 1 0 37632 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_353
timestamp 1669390400
transform 1 0 40880 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_357
timestamp 1669390400
transform 1 0 41328 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_365
timestamp 1669390400
transform 1 0 42224 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_369
timestamp 1669390400
transform 1 0 42672 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_373
timestamp 1669390400
transform 1 0 43120 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_376
timestamp 1669390400
transform 1 0 43456 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_378
timestamp 1669390400
transform 1 0 43680 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_387
timestamp 1669390400
transform 1 0 44688 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1669390400
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_395
timestamp 1669390400
transform 1 0 45584 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_407
timestamp 1669390400
transform 1 0 46928 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_415
timestamp 1669390400
transform 1 0 47824 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_423
timestamp 1669390400
transform 1 0 48720 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_433
timestamp 1669390400
transform 1 0 49840 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_443
timestamp 1669390400
transform 1 0 50960 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_451
timestamp 1669390400
transform 1 0 51856 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_459
timestamp 1669390400
transform 1 0 52752 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_463
timestamp 1669390400
transform 1 0 53200 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_470
timestamp 1669390400
transform 1 0 53984 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_480
timestamp 1669390400
transform 1 0 55104 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_486
timestamp 1669390400
transform 1 0 55776 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_494
timestamp 1669390400
transform 1 0 56672 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_502
timestamp 1669390400
transform 1 0 57568 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_506
timestamp 1669390400
transform 1 0 58016 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_508
timestamp 1669390400
transform 1 0 58240 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_4
timestamp 1669390400
transform 1 0 1792 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_7
timestamp 1669390400
transform 1 0 2128 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_11
timestamp 1669390400
transform 1 0 2576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_15
timestamp 1669390400
transform 1 0 3024 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_18
timestamp 1669390400
transform 1 0 3360 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_22
timestamp 1669390400
transform 1 0 3808 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_24
timestamp 1669390400
transform 1 0 4032 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_27
timestamp 1669390400
transform 1 0 4368 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_35
timestamp 1669390400
transform 1 0 5264 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_39
timestamp 1669390400
transform 1 0 5712 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_43
timestamp 1669390400
transform 1 0 6160 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_50
timestamp 1669390400
transform 1 0 6944 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_58
timestamp 1669390400
transform 1 0 7840 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_62
timestamp 1669390400
transform 1 0 8288 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_66
timestamp 1669390400
transform 1 0 8736 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1669390400
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_75
timestamp 1669390400
transform 1 0 9744 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_82
timestamp 1669390400
transform 1 0 10528 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_92
timestamp 1669390400
transform 1 0 11648 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_110
timestamp 1669390400
transform 1 0 13664 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_112
timestamp 1669390400
transform 1 0 13888 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_115
timestamp 1669390400
transform 1 0 14224 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_119
timestamp 1669390400
transform 1 0 14672 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_129
timestamp 1669390400
transform 1 0 15792 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_133
timestamp 1669390400
transform 1 0 16240 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_147
timestamp 1669390400
transform 1 0 17808 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_149
timestamp 1669390400
transform 1 0 18032 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_186
timestamp 1669390400
transform 1 0 22176 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_194
timestamp 1669390400
transform 1 0 23072 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_198
timestamp 1669390400
transform 1 0 23520 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_202
timestamp 1669390400
transform 1 0 23968 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_206
timestamp 1669390400
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_210
timestamp 1669390400
transform 1 0 24864 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_223
timestamp 1669390400
transform 1 0 26320 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_227
timestamp 1669390400
transform 1 0 26768 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_229
timestamp 1669390400
transform 1 0 26992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_232
timestamp 1669390400
transform 1 0 27328 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_268
timestamp 1669390400
transform 1 0 31360 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_272
timestamp 1669390400
transform 1 0 31808 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_276
timestamp 1669390400
transform 1 0 32256 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_280
timestamp 1669390400
transform 1 0 32704 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_302
timestamp 1669390400
transform 1 0 35168 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_305
timestamp 1669390400
transform 1 0 35504 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_309
timestamp 1669390400
transform 1 0 35952 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_313
timestamp 1669390400
transform 1 0 36400 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_317
timestamp 1669390400
transform 1 0 36848 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_319
timestamp 1669390400
transform 1 0 37072 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_374
timestamp 1669390400
transform 1 0 43232 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_378
timestamp 1669390400
transform 1 0 43680 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_385
timestamp 1669390400
transform 1 0 44464 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_389
timestamp 1669390400
transform 1 0 44912 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_391
timestamp 1669390400
transform 1 0 45136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_400
timestamp 1669390400
transform 1 0 46144 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_404
timestamp 1669390400
transform 1 0 46592 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_408
timestamp 1669390400
transform 1 0 47040 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_412
timestamp 1669390400
transform 1 0 47488 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_420
timestamp 1669390400
transform 1 0 48384 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_424
timestamp 1669390400
transform 1 0 48832 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_428
timestamp 1669390400
transform 1 0 49280 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_435
timestamp 1669390400
transform 1 0 50064 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_443
timestamp 1669390400
transform 1 0 50960 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_451
timestamp 1669390400
transform 1 0 51856 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_466
timestamp 1669390400
transform 1 0 53536 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_470
timestamp 1669390400
transform 1 0 53984 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_474
timestamp 1669390400
transform 1 0 54432 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_476
timestamp 1669390400
transform 1 0 54656 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_483
timestamp 1669390400
transform 1 0 55440 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_487
timestamp 1669390400
transform 1 0 55888 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_491
timestamp 1669390400
transform 1 0 56336 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_495
timestamp 1669390400
transform 1 0 56784 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_499
timestamp 1669390400
transform 1 0 57232 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_502
timestamp 1669390400
transform 1 0 57568 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_506
timestamp 1669390400
transform 1 0 58016 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_508
timestamp 1669390400
transform 1 0 58240 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_9
timestamp 1669390400
transform 1 0 2352 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_17
timestamp 1669390400
transform 1 0 3248 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_25
timestamp 1669390400
transform 1 0 4144 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_27
timestamp 1669390400
transform 1 0 4368 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1669390400
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_44
timestamp 1669390400
transform 1 0 6272 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_52
timestamp 1669390400
transform 1 0 7168 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_56
timestamp 1669390400
transform 1 0 7616 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_59
timestamp 1669390400
transform 1 0 7952 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_61
timestamp 1669390400
transform 1 0 8176 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_68
timestamp 1669390400
transform 1 0 8960 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_79
timestamp 1669390400
transform 1 0 10192 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_89
timestamp 1669390400
transform 1 0 11312 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_97
timestamp 1669390400
transform 1 0 12208 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_111
timestamp 1669390400
transform 1 0 13776 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_115
timestamp 1669390400
transform 1 0 14224 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_119
timestamp 1669390400
transform 1 0 14672 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_123
timestamp 1669390400
transform 1 0 15120 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_129
timestamp 1669390400
transform 1 0 15792 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_133
timestamp 1669390400
transform 1 0 16240 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_137
timestamp 1669390400
transform 1 0 16688 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_141
timestamp 1669390400
transform 1 0 17136 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_157
timestamp 1669390400
transform 1 0 18928 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_167
timestamp 1669390400
transform 1 0 20048 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_171
timestamp 1669390400
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_175
timestamp 1669390400
transform 1 0 20944 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_185
timestamp 1669390400
transform 1 0 22064 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_193
timestamp 1669390400
transform 1 0 22960 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_201
timestamp 1669390400
transform 1 0 23856 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_205
timestamp 1669390400
transform 1 0 24304 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_221
timestamp 1669390400
transform 1 0 26096 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_227
timestamp 1669390400
transform 1 0 26768 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_253
timestamp 1669390400
transform 1 0 29680 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_261
timestamp 1669390400
transform 1 0 30576 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_265
timestamp 1669390400
transform 1 0 31024 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_269
timestamp 1669390400
transform 1 0 31472 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_285
timestamp 1669390400
transform 1 0 33264 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_294
timestamp 1669390400
transform 1 0 34272 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_310
timestamp 1669390400
transform 1 0 36064 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_325
timestamp 1669390400
transform 1 0 37744 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_342
timestamp 1669390400
transform 1 0 39648 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_378
timestamp 1669390400
transform 1 0 43680 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_386
timestamp 1669390400
transform 1 0 44576 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_405
timestamp 1669390400
transform 1 0 46704 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_409
timestamp 1669390400
transform 1 0 47152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_415
timestamp 1669390400
transform 1 0 47824 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_423
timestamp 1669390400
transform 1 0 48720 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_427
timestamp 1669390400
transform 1 0 49168 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_437
timestamp 1669390400
transform 1 0 50288 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_439
timestamp 1669390400
transform 1 0 50512 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_442
timestamp 1669390400
transform 1 0 50848 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_450
timestamp 1669390400
transform 1 0 51744 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_458
timestamp 1669390400
transform 1 0 52640 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1669390400
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_463
timestamp 1669390400
transform 1 0 53200 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_466
timestamp 1669390400
transform 1 0 53536 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_468
timestamp 1669390400
transform 1 0 53760 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_471
timestamp 1669390400
transform 1 0 54096 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_479
timestamp 1669390400
transform 1 0 54992 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_487
timestamp 1669390400
transform 1 0 55888 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_491
timestamp 1669390400
transform 1 0 56336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_497
timestamp 1669390400
transform 1 0 57008 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_501
timestamp 1669390400
transform 1 0 57456 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_505
timestamp 1669390400
transform 1 0 57904 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_6
timestamp 1669390400
transform 1 0 2016 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_20
timestamp 1669390400
transform 1 0 3584 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_28
timestamp 1669390400
transform 1 0 4480 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_30
timestamp 1669390400
transform 1 0 4704 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_43
timestamp 1669390400
transform 1 0 6160 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_47
timestamp 1669390400
transform 1 0 6608 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_57
timestamp 1669390400
transform 1 0 7728 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_61
timestamp 1669390400
transform 1 0 8176 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_82
timestamp 1669390400
transform 1 0 10528 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_89
timestamp 1669390400
transform 1 0 11312 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_97
timestamp 1669390400
transform 1 0 12208 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_107
timestamp 1669390400
transform 1 0 13328 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_117
timestamp 1669390400
transform 1 0 14448 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_125
timestamp 1669390400
transform 1 0 15344 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1669390400
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_147
timestamp 1669390400
transform 1 0 17808 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_151
timestamp 1669390400
transform 1 0 18256 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_165
timestamp 1669390400
transform 1 0 19824 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_181
timestamp 1669390400
transform 1 0 21616 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_183
timestamp 1669390400
transform 1 0 21840 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_186
timestamp 1669390400
transform 1 0 22176 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_200
timestamp 1669390400
transform 1 0 23744 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_204
timestamp 1669390400
transform 1 0 24192 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_222
timestamp 1669390400
transform 1 0 26208 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_226
timestamp 1669390400
transform 1 0 26656 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_233
timestamp 1669390400
transform 1 0 27440 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_237
timestamp 1669390400
transform 1 0 27888 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_241
timestamp 1669390400
transform 1 0 28336 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_244
timestamp 1669390400
transform 1 0 28672 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_248
timestamp 1669390400
transform 1 0 29120 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_252
timestamp 1669390400
transform 1 0 29568 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_276
timestamp 1669390400
transform 1 0 32256 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_321
timestamp 1669390400
transform 1 0 37296 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_325
timestamp 1669390400
transform 1 0 37744 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_329
timestamp 1669390400
transform 1 0 38192 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_331
timestamp 1669390400
transform 1 0 38416 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_334
timestamp 1669390400
transform 1 0 38752 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_352
timestamp 1669390400
transform 1 0 40768 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_360
timestamp 1669390400
transform 1 0 41664 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_392
timestamp 1669390400
transform 1 0 45248 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_402
timestamp 1669390400
transform 1 0 46368 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_406
timestamp 1669390400
transform 1 0 46816 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_420
timestamp 1669390400
transform 1 0 48384 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_424
timestamp 1669390400
transform 1 0 48832 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_428
timestamp 1669390400
transform 1 0 49280 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_446
timestamp 1669390400
transform 1 0 51296 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_454
timestamp 1669390400
transform 1 0 52192 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_460
timestamp 1669390400
transform 1 0 52864 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_464
timestamp 1669390400
transform 1 0 53312 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_468
timestamp 1669390400
transform 1 0 53760 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_476
timestamp 1669390400
transform 1 0 54656 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_478
timestamp 1669390400
transform 1 0 54880 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_481
timestamp 1669390400
transform 1 0 55216 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_485
timestamp 1669390400
transform 1 0 55664 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_488
timestamp 1669390400
transform 1 0 56000 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_492
timestamp 1669390400
transform 1 0 56448 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1669390400
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_499
timestamp 1669390400
transform 1 0 57232 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_502
timestamp 1669390400
transform 1 0 57568 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_506
timestamp 1669390400
transform 1 0 58016 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_508
timestamp 1669390400
transform 1 0 58240 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_6
timestamp 1669390400
transform 1 0 2016 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_10
timestamp 1669390400
transform 1 0 2464 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_18
timestamp 1669390400
transform 1 0 3360 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_24
timestamp 1669390400
transform 1 0 4032 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_28
timestamp 1669390400
transform 1 0 4480 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_31
timestamp 1669390400
transform 1 0 4816 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_42
timestamp 1669390400
transform 1 0 6048 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_50
timestamp 1669390400
transform 1 0 6944 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_57
timestamp 1669390400
transform 1 0 7728 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_59
timestamp 1669390400
transform 1 0 7952 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_62
timestamp 1669390400
transform 1 0 8288 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_79
timestamp 1669390400
transform 1 0 10192 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_83
timestamp 1669390400
transform 1 0 10640 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_87
timestamp 1669390400
transform 1 0 11088 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_91
timestamp 1669390400
transform 1 0 11536 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_95
timestamp 1669390400
transform 1 0 11984 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_99
timestamp 1669390400
transform 1 0 12432 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_114
timestamp 1669390400
transform 1 0 14112 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_118
timestamp 1669390400
transform 1 0 14560 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_122
timestamp 1669390400
transform 1 0 15008 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_126
timestamp 1669390400
transform 1 0 15456 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_134
timestamp 1669390400
transform 1 0 16352 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_144
timestamp 1669390400
transform 1 0 17472 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_152
timestamp 1669390400
transform 1 0 18368 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_156
timestamp 1669390400
transform 1 0 18816 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_162
timestamp 1669390400
transform 1 0 19488 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_183
timestamp 1669390400
transform 1 0 21840 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_187
timestamp 1669390400
transform 1 0 22288 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_194
timestamp 1669390400
transform 1 0 23072 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_201
timestamp 1669390400
transform 1 0 23856 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_205
timestamp 1669390400
transform 1 0 24304 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_209
timestamp 1669390400
transform 1 0 24752 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_257
timestamp 1669390400
transform 1 0 30128 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_267
timestamp 1669390400
transform 1 0 31248 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_274
timestamp 1669390400
transform 1 0 32032 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_282
timestamp 1669390400
transform 1 0 32928 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_356
timestamp 1669390400
transform 1 0 41216 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_360
timestamp 1669390400
transform 1 0 41664 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1669390400
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_456
timestamp 1669390400
transform 1 0 52416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1669390400
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_463
timestamp 1669390400
transform 1 0 53200 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_495
timestamp 1669390400
transform 1 0 56784 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_503
timestamp 1669390400
transform 1 0 57680 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_507
timestamp 1669390400
transform 1 0 58128 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_17
timestamp 1669390400
transform 1 0 3248 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_25
timestamp 1669390400
transform 1 0 4144 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_29
timestamp 1669390400
transform 1 0 4592 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_33
timestamp 1669390400
transform 1 0 5040 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_37
timestamp 1669390400
transform 1 0 5488 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_41
timestamp 1669390400
transform 1 0 5936 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_51
timestamp 1669390400
transform 1 0 7056 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_61
timestamp 1669390400
transform 1 0 8176 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_65
timestamp 1669390400
transform 1 0 8624 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_69
timestamp 1669390400
transform 1 0 9072 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_77
timestamp 1669390400
transform 1 0 9968 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_81
timestamp 1669390400
transform 1 0 10416 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_83
timestamp 1669390400
transform 1 0 10640 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_86
timestamp 1669390400
transform 1 0 10976 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_90
timestamp 1669390400
transform 1 0 11424 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_94
timestamp 1669390400
transform 1 0 11872 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_98
timestamp 1669390400
transform 1 0 12320 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_102
timestamp 1669390400
transform 1 0 12768 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_106
timestamp 1669390400
transform 1 0 13216 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_115
timestamp 1669390400
transform 1 0 14224 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_123
timestamp 1669390400
transform 1 0 15120 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_129
timestamp 1669390400
transform 1 0 15792 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_137
timestamp 1669390400
transform 1 0 16688 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_150
timestamp 1669390400
transform 1 0 18144 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_162
timestamp 1669390400
transform 1 0 19488 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_166
timestamp 1669390400
transform 1 0 19936 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_170
timestamp 1669390400
transform 1 0 20384 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_178
timestamp 1669390400
transform 1 0 21280 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_186
timestamp 1669390400
transform 1 0 22176 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_196
timestamp 1669390400
transform 1 0 23296 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_211
timestamp 1669390400
transform 1 0 24976 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_218
timestamp 1669390400
transform 1 0 25760 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_222
timestamp 1669390400
transform 1 0 26208 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_230
timestamp 1669390400
transform 1 0 27104 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_234
timestamp 1669390400
transform 1 0 27552 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_238
timestamp 1669390400
transform 1 0 28000 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_242
timestamp 1669390400
transform 1 0 28448 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_246
timestamp 1669390400
transform 1 0 28896 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_250
timestamp 1669390400
transform 1 0 29344 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_260
timestamp 1669390400
transform 1 0 30464 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_264
timestamp 1669390400
transform 1 0 30912 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_267
timestamp 1669390400
transform 1 0 31248 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_273
timestamp 1669390400
transform 1 0 31920 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_277
timestamp 1669390400
transform 1 0 32368 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_315
timestamp 1669390400
transform 1 0 36624 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_333
timestamp 1669390400
transform 1 0 38640 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_349
timestamp 1669390400
transform 1 0 40432 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_353
timestamp 1669390400
transform 1 0 40880 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_421
timestamp 1669390400
transform 1 0 48496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1669390400
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1669390400
transform 1 0 49280 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1669390400
transform 1 0 56448 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1669390400
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_499
timestamp 1669390400
transform 1 0 57232 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_507
timestamp 1669390400
transform 1 0 58128 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_8
timestamp 1669390400
transform 1 0 2240 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_16
timestamp 1669390400
transform 1 0 3136 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_24
timestamp 1669390400
transform 1 0 4032 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1669390400
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_40
timestamp 1669390400
transform 1 0 5824 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_50
timestamp 1669390400
transform 1 0 6944 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_52
timestamp 1669390400
transform 1 0 7168 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_55
timestamp 1669390400
transform 1 0 7504 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_63
timestamp 1669390400
transform 1 0 8400 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_73
timestamp 1669390400
transform 1 0 9520 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_77
timestamp 1669390400
transform 1 0 9968 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_84
timestamp 1669390400
transform 1 0 10752 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_115
timestamp 1669390400
transform 1 0 14224 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_125
timestamp 1669390400
transform 1 0 15344 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_131
timestamp 1669390400
transform 1 0 16016 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_140
timestamp 1669390400
transform 1 0 17024 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_165
timestamp 1669390400
transform 1 0 19824 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_169
timestamp 1669390400
transform 1 0 20272 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_205
timestamp 1669390400
transform 1 0 24304 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_220
timestamp 1669390400
transform 1 0 25984 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_230
timestamp 1669390400
transform 1 0 27104 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_234
timestamp 1669390400
transform 1 0 27552 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_236
timestamp 1669390400
transform 1 0 27776 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_239
timestamp 1669390400
transform 1 0 28112 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_245
timestamp 1669390400
transform 1 0 28784 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_257
timestamp 1669390400
transform 1 0 30128 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_259
timestamp 1669390400
transform 1 0 30352 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_262
timestamp 1669390400
transform 1 0 30688 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_276
timestamp 1669390400
transform 1 0 32256 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_280
timestamp 1669390400
transform 1 0 32704 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_290
timestamp 1669390400
transform 1 0 33824 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_294
timestamp 1669390400
transform 1 0 34272 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_297
timestamp 1669390400
transform 1 0 34608 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_307
timestamp 1669390400
transform 1 0 35728 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_317
timestamp 1669390400
transform 1 0 36848 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_328
timestamp 1669390400
transform 1 0 38080 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_338
timestamp 1669390400
transform 1 0 39200 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_342
timestamp 1669390400
transform 1 0 39648 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_378
timestamp 1669390400
transform 1 0 43680 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_386
timestamp 1669390400
transform 1 0 44576 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_456
timestamp 1669390400
transform 1 0 52416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1669390400
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_463
timestamp 1669390400
transform 1 0 53200 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_495
timestamp 1669390400
transform 1 0 56784 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_503
timestamp 1669390400
transform 1 0 57680 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_507
timestamp 1669390400
transform 1 0 58128 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_5
timestamp 1669390400
transform 1 0 1904 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_9
timestamp 1669390400
transform 1 0 2352 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_17
timestamp 1669390400
transform 1 0 3248 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_27
timestamp 1669390400
transform 1 0 4368 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_29
timestamp 1669390400
transform 1 0 4592 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_32
timestamp 1669390400
transform 1 0 4928 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_40
timestamp 1669390400
transform 1 0 5824 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_50
timestamp 1669390400
transform 1 0 6944 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_54
timestamp 1669390400
transform 1 0 7392 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_58
timestamp 1669390400
transform 1 0 7840 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1669390400
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_77
timestamp 1669390400
transform 1 0 9968 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_92
timestamp 1669390400
transform 1 0 11648 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_96
timestamp 1669390400
transform 1 0 12096 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_115
timestamp 1669390400
transform 1 0 14224 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_123
timestamp 1669390400
transform 1 0 15120 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_129
timestamp 1669390400
transform 1 0 15792 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_133
timestamp 1669390400
transform 1 0 16240 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_168
timestamp 1669390400
transform 1 0 20160 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_170
timestamp 1669390400
transform 1 0 20384 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_177
timestamp 1669390400
transform 1 0 21168 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_185
timestamp 1669390400
transform 1 0 22064 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_193
timestamp 1669390400
transform 1 0 22960 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_197
timestamp 1669390400
transform 1 0 23408 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_205
timestamp 1669390400
transform 1 0 24304 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_211
timestamp 1669390400
transform 1 0 24976 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_218
timestamp 1669390400
transform 1 0 25760 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_222
timestamp 1669390400
transform 1 0 26208 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_226
timestamp 1669390400
transform 1 0 26656 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_228
timestamp 1669390400
transform 1 0 26880 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_235
timestamp 1669390400
transform 1 0 27664 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_239
timestamp 1669390400
transform 1 0 28112 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_241
timestamp 1669390400
transform 1 0 28336 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_254
timestamp 1669390400
transform 1 0 29792 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_258
timestamp 1669390400
transform 1 0 30240 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_264
timestamp 1669390400
transform 1 0 30912 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_272
timestamp 1669390400
transform 1 0 31808 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_276
timestamp 1669390400
transform 1 0 32256 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1669390400
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_295
timestamp 1669390400
transform 1 0 34384 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_305
timestamp 1669390400
transform 1 0 35504 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_314
timestamp 1669390400
transform 1 0 36512 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_318
timestamp 1669390400
transform 1 0 36960 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_322
timestamp 1669390400
transform 1 0 37408 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_332
timestamp 1669390400
transform 1 0 38528 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_340
timestamp 1669390400
transform 1 0 39424 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_348
timestamp 1669390400
transform 1 0 40320 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_352
timestamp 1669390400
transform 1 0 40768 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_364
timestamp 1669390400
transform 1 0 42112 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_396
timestamp 1669390400
transform 1 0 45696 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_412
timestamp 1669390400
transform 1 0 47488 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_420
timestamp 1669390400
transform 1 0 48384 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_424
timestamp 1669390400
transform 1 0 48832 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_428
timestamp 1669390400
transform 1 0 49280 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_460
timestamp 1669390400
transform 1 0 52864 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_468
timestamp 1669390400
transform 1 0 53760 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_472
timestamp 1669390400
transform 1 0 54208 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_475
timestamp 1669390400
transform 1 0 54544 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_491
timestamp 1669390400
transform 1 0 56336 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_495
timestamp 1669390400
transform 1 0 56784 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_499
timestamp 1669390400
transform 1 0 57232 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_507
timestamp 1669390400
transform 1 0 58128 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_5
timestamp 1669390400
transform 1 0 1904 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_11
timestamp 1669390400
transform 1 0 2576 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_19
timestamp 1669390400
transform 1 0 3472 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_23
timestamp 1669390400
transform 1 0 3920 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_43
timestamp 1669390400
transform 1 0 6160 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_47
timestamp 1669390400
transform 1 0 6608 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_51
timestamp 1669390400
transform 1 0 7056 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_68
timestamp 1669390400
transform 1 0 8960 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_72
timestamp 1669390400
transform 1 0 9408 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_79
timestamp 1669390400
transform 1 0 10192 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_94
timestamp 1669390400
transform 1 0 11872 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_96
timestamp 1669390400
transform 1 0 12096 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1669390400
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_108
timestamp 1669390400
transform 1 0 13440 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_110
timestamp 1669390400
transform 1 0 13664 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_119
timestamp 1669390400
transform 1 0 14672 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_123
timestamp 1669390400
transform 1 0 15120 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_147
timestamp 1669390400
transform 1 0 17808 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_155
timestamp 1669390400
transform 1 0 18704 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_157
timestamp 1669390400
transform 1 0 18928 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_160
timestamp 1669390400
transform 1 0 19264 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_168
timestamp 1669390400
transform 1 0 20160 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_175
timestamp 1669390400
transform 1 0 20944 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_179
timestamp 1669390400
transform 1 0 21392 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_185
timestamp 1669390400
transform 1 0 22064 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_187
timestamp 1669390400
transform 1 0 22288 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_193
timestamp 1669390400
transform 1 0 22960 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_201
timestamp 1669390400
transform 1 0 23856 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_209
timestamp 1669390400
transform 1 0 24752 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_213
timestamp 1669390400
transform 1 0 25200 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_217
timestamp 1669390400
transform 1 0 25648 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_223
timestamp 1669390400
transform 1 0 26320 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_238
timestamp 1669390400
transform 1 0 28000 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_240
timestamp 1669390400
transform 1 0 28224 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_250
timestamp 1669390400
transform 1 0 29344 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_264
timestamp 1669390400
transform 1 0 30912 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_270
timestamp 1669390400
transform 1 0 31584 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_274
timestamp 1669390400
transform 1 0 32032 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_282
timestamp 1669390400
transform 1 0 32928 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_285
timestamp 1669390400
transform 1 0 33264 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_292
timestamp 1669390400
transform 1 0 34048 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_318
timestamp 1669390400
transform 1 0 36960 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_321
timestamp 1669390400
transform 1 0 37296 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_329
timestamp 1669390400
transform 1 0 38192 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_354
timestamp 1669390400
transform 1 0 40992 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_361
timestamp 1669390400
transform 1 0 41776 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_375
timestamp 1669390400
transform 1 0 43344 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_383
timestamp 1669390400
transform 1 0 44240 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_387
timestamp 1669390400
transform 1 0 44688 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1669390400
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_392
timestamp 1669390400
transform 1 0 45248 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_456
timestamp 1669390400
transform 1 0 52416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_460
timestamp 1669390400
transform 1 0 52864 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_463
timestamp 1669390400
transform 1 0 53200 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_495
timestamp 1669390400
transform 1 0 56784 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_503
timestamp 1669390400
transform 1 0 57680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_507
timestamp 1669390400
transform 1 0 58128 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_9
timestamp 1669390400
transform 1 0 2352 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_19
timestamp 1669390400
transform 1 0 3472 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_23
timestamp 1669390400
transform 1 0 3920 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_33
timestamp 1669390400
transform 1 0 5040 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_37
timestamp 1669390400
transform 1 0 5488 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_46
timestamp 1669390400
transform 1 0 6496 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_59
timestamp 1669390400
transform 1 0 7952 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_63
timestamp 1669390400
transform 1 0 8400 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1669390400
transform 1 0 9184 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_73
timestamp 1669390400
transform 1 0 9520 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_75
timestamp 1669390400
transform 1 0 9744 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_78
timestamp 1669390400
transform 1 0 10080 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_120
timestamp 1669390400
transform 1 0 14784 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_130
timestamp 1669390400
transform 1 0 15904 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_134
timestamp 1669390400
transform 1 0 16352 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1669390400
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_144
timestamp 1669390400
transform 1 0 17472 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_147
timestamp 1669390400
transform 1 0 17808 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_172
timestamp 1669390400
transform 1 0 20608 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_176
timestamp 1669390400
transform 1 0 21056 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_183
timestamp 1669390400
transform 1 0 21840 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_191
timestamp 1669390400
transform 1 0 22736 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_206
timestamp 1669390400
transform 1 0 24416 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_210
timestamp 1669390400
transform 1 0 24864 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1669390400
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_215
timestamp 1669390400
transform 1 0 25424 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_219
timestamp 1669390400
transform 1 0 25872 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_223
timestamp 1669390400
transform 1 0 26320 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_233
timestamp 1669390400
transform 1 0 27440 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_241
timestamp 1669390400
transform 1 0 28336 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_245
timestamp 1669390400
transform 1 0 28784 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_258
timestamp 1669390400
transform 1 0 30240 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_268
timestamp 1669390400
transform 1 0 31360 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_270
timestamp 1669390400
transform 1 0 31584 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1669390400
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_286
timestamp 1669390400
transform 1 0 33376 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_292
timestamp 1669390400
transform 1 0 34048 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_300
timestamp 1669390400
transform 1 0 34944 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_310
timestamp 1669390400
transform 1 0 36064 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_318
timestamp 1669390400
transform 1 0 36960 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_322
timestamp 1669390400
transform 1 0 37408 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_325
timestamp 1669390400
transform 1 0 37744 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_335
timestamp 1669390400
transform 1 0 38864 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_351
timestamp 1669390400
transform 1 0 40656 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_357
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_363
timestamp 1669390400
transform 1 0 42000 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_377
timestamp 1669390400
transform 1 0 43568 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_409
timestamp 1669390400
transform 1 0 47152 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_425
timestamp 1669390400
transform 1 0 48944 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_43_428
timestamp 1669390400
transform 1 0 49280 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_492
timestamp 1669390400
transform 1 0 56448 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_496
timestamp 1669390400
transform 1 0 56896 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_499
timestamp 1669390400
transform 1 0 57232 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_507
timestamp 1669390400
transform 1 0 58128 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_6
timestamp 1669390400
transform 1 0 2016 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_10
timestamp 1669390400
transform 1 0 2464 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_20
timestamp 1669390400
transform 1 0 3584 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_28
timestamp 1669390400
transform 1 0 4480 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1669390400
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_37
timestamp 1669390400
transform 1 0 5488 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_47
timestamp 1669390400
transform 1 0 6608 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_85
timestamp 1669390400
transform 1 0 10864 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_95
timestamp 1669390400
transform 1 0 11984 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_103
timestamp 1669390400
transform 1 0 12880 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1669390400
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_108
timestamp 1669390400
transform 1 0 13440 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_125
timestamp 1669390400
transform 1 0 15344 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_129
timestamp 1669390400
transform 1 0 15792 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_133
timestamp 1669390400
transform 1 0 16240 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_137
timestamp 1669390400
transform 1 0 16688 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_141
timestamp 1669390400
transform 1 0 17136 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_149
timestamp 1669390400
transform 1 0 18032 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_157
timestamp 1669390400
transform 1 0 18928 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_165
timestamp 1669390400
transform 1 0 19824 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1669390400
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_179
timestamp 1669390400
transform 1 0 21392 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_188
timestamp 1669390400
transform 1 0 22400 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_192
timestamp 1669390400
transform 1 0 22848 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_204
timestamp 1669390400
transform 1 0 24192 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_208
timestamp 1669390400
transform 1 0 24640 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_212
timestamp 1669390400
transform 1 0 25088 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_220
timestamp 1669390400
transform 1 0 25984 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_228
timestamp 1669390400
transform 1 0 26880 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_242
timestamp 1669390400
transform 1 0 28448 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_244
timestamp 1669390400
transform 1 0 28672 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1669390400
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_250
timestamp 1669390400
transform 1 0 29344 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_254
timestamp 1669390400
transform 1 0 29792 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_258
timestamp 1669390400
transform 1 0 30240 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_270
timestamp 1669390400
transform 1 0 31584 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_278
timestamp 1669390400
transform 1 0 32480 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_285
timestamp 1669390400
transform 1 0 33264 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_289
timestamp 1669390400
transform 1 0 33712 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_293
timestamp 1669390400
transform 1 0 34160 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_297
timestamp 1669390400
transform 1 0 34608 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_299
timestamp 1669390400
transform 1 0 34832 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_302
timestamp 1669390400
transform 1 0 35168 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_310
timestamp 1669390400
transform 1 0 36064 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_314
timestamp 1669390400
transform 1 0 36512 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1669390400
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_321
timestamp 1669390400
transform 1 0 37296 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_348
timestamp 1669390400
transform 1 0 40320 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_352
timestamp 1669390400
transform 1 0 40768 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_356
timestamp 1669390400
transform 1 0 41216 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_369
timestamp 1669390400
transform 1 0 42672 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1669390400
transform 1 0 44464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1669390400
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_392
timestamp 1669390400
transform 1 0 45248 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_456
timestamp 1669390400
transform 1 0 52416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_460
timestamp 1669390400
transform 1 0 52864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_44_463
timestamp 1669390400
transform 1 0 53200 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_44_495
timestamp 1669390400
transform 1 0 56784 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_503
timestamp 1669390400
transform 1 0 57680 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_507
timestamp 1669390400
transform 1 0 58128 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_9
timestamp 1669390400
transform 1 0 2352 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_19
timestamp 1669390400
transform 1 0 3472 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_29
timestamp 1669390400
transform 1 0 4592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_35
timestamp 1669390400
transform 1 0 5264 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_52
timestamp 1669390400
transform 1 0 7168 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_61
timestamp 1669390400
transform 1 0 8176 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_63
timestamp 1669390400
transform 1 0 8400 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_66
timestamp 1669390400
transform 1 0 8736 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1669390400
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_73
timestamp 1669390400
transform 1 0 9520 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_81
timestamp 1669390400
transform 1 0 10416 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_89
timestamp 1669390400
transform 1 0 11312 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_93
timestamp 1669390400
transform 1 0 11760 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_96
timestamp 1669390400
transform 1 0 12096 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_103
timestamp 1669390400
transform 1 0 12880 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_105
timestamp 1669390400
transform 1 0 13104 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_112
timestamp 1669390400
transform 1 0 13888 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_120
timestamp 1669390400
transform 1 0 14784 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_122
timestamp 1669390400
transform 1 0 15008 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_125
timestamp 1669390400
transform 1 0 15344 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_129
timestamp 1669390400
transform 1 0 15792 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1669390400
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_144
timestamp 1669390400
transform 1 0 17472 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_188
timestamp 1669390400
transform 1 0 22400 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_192
timestamp 1669390400
transform 1 0 22848 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1669390400
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_215
timestamp 1669390400
transform 1 0 25424 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_217
timestamp 1669390400
transform 1 0 25648 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_220
timestamp 1669390400
transform 1 0 25984 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_224
timestamp 1669390400
transform 1 0 26432 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_238
timestamp 1669390400
transform 1 0 28000 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_248
timestamp 1669390400
transform 1 0 29120 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_254
timestamp 1669390400
transform 1 0 29792 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_258
timestamp 1669390400
transform 1 0 30240 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_262
timestamp 1669390400
transform 1 0 30688 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1669390400
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_286
timestamp 1669390400
transform 1 0 33376 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_313
timestamp 1669390400
transform 1 0 36400 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_315
timestamp 1669390400
transform 1 0 36624 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_321
timestamp 1669390400
transform 1 0 37296 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_325
timestamp 1669390400
transform 1 0 37744 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_337
timestamp 1669390400
transform 1 0 39088 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_343
timestamp 1669390400
transform 1 0 39760 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_347
timestamp 1669390400
transform 1 0 40208 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_351
timestamp 1669390400
transform 1 0 40656 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_357
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_363
timestamp 1669390400
transform 1 0 42000 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_365
timestamp 1669390400
transform 1 0 42224 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_371
timestamp 1669390400
transform 1 0 42896 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_403
timestamp 1669390400
transform 1 0 46480 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_419
timestamp 1669390400
transform 1 0 48272 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_423
timestamp 1669390400
transform 1 0 48720 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_425
timestamp 1669390400
transform 1 0 48944 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_45_428
timestamp 1669390400
transform 1 0 49280 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_492
timestamp 1669390400
transform 1 0 56448 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_496
timestamp 1669390400
transform 1 0 56896 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_499
timestamp 1669390400
transform 1 0 57232 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_507
timestamp 1669390400
transform 1 0 58128 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_17
timestamp 1669390400
transform 1 0 3248 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_27
timestamp 1669390400
transform 1 0 4368 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_31
timestamp 1669390400
transform 1 0 4816 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1669390400
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_37
timestamp 1669390400
transform 1 0 5488 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_43
timestamp 1669390400
transform 1 0 6160 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_51
timestamp 1669390400
transform 1 0 7056 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_53
timestamp 1669390400
transform 1 0 7280 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_56
timestamp 1669390400
transform 1 0 7616 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_64
timestamp 1669390400
transform 1 0 8512 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_74
timestamp 1669390400
transform 1 0 9632 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_84
timestamp 1669390400
transform 1 0 10752 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_94
timestamp 1669390400
transform 1 0 11872 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_98
timestamp 1669390400
transform 1 0 12320 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_101
timestamp 1669390400
transform 1 0 12656 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1669390400
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_108
timestamp 1669390400
transform 1 0 13440 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_119
timestamp 1669390400
transform 1 0 14672 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_121
timestamp 1669390400
transform 1 0 14896 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_124
timestamp 1669390400
transform 1 0 15232 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_128
timestamp 1669390400
transform 1 0 15680 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_132
timestamp 1669390400
transform 1 0 16128 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_136
timestamp 1669390400
transform 1 0 16576 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_149
timestamp 1669390400
transform 1 0 18032 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_157
timestamp 1669390400
transform 1 0 18928 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_161
timestamp 1669390400
transform 1 0 19376 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_170
timestamp 1669390400
transform 1 0 20384 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1669390400
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_179
timestamp 1669390400
transform 1 0 21392 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_190
timestamp 1669390400
transform 1 0 22624 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_197
timestamp 1669390400
transform 1 0 23408 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_207
timestamp 1669390400
transform 1 0 24528 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_213
timestamp 1669390400
transform 1 0 25200 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_217
timestamp 1669390400
transform 1 0 25648 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_221
timestamp 1669390400
transform 1 0 26096 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_239
timestamp 1669390400
transform 1 0 28112 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_243
timestamp 1669390400
transform 1 0 28560 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1669390400
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_250
timestamp 1669390400
transform 1 0 29344 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_256
timestamp 1669390400
transform 1 0 30016 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_260
timestamp 1669390400
transform 1 0 30464 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_266
timestamp 1669390400
transform 1 0 31136 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_274
timestamp 1669390400
transform 1 0 32032 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_282
timestamp 1669390400
transform 1 0 32928 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_286
timestamp 1669390400
transform 1 0 33376 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_299
timestamp 1669390400
transform 1 0 34832 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_303
timestamp 1669390400
transform 1 0 35280 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_311
timestamp 1669390400
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_315
timestamp 1669390400
transform 1 0 36624 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_318
timestamp 1669390400
transform 1 0 36960 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_321
timestamp 1669390400
transform 1 0 37296 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_326
timestamp 1669390400
transform 1 0 37856 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_330
timestamp 1669390400
transform 1 0 38304 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_342
timestamp 1669390400
transform 1 0 39648 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_346
timestamp 1669390400
transform 1 0 40096 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_371
timestamp 1669390400
transform 1 0 42896 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_375
timestamp 1669390400
transform 1 0 43344 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1669390400
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_392
timestamp 1669390400
transform 1 0 45248 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_408
timestamp 1669390400
transform 1 0 47040 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_410
timestamp 1669390400
transform 1 0 47264 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_417
timestamp 1669390400
transform 1 0 48048 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_449
timestamp 1669390400
transform 1 0 51632 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_457
timestamp 1669390400
transform 1 0 52528 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_463
timestamp 1669390400
transform 1 0 53200 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_479
timestamp 1669390400
transform 1 0 54992 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_487
timestamp 1669390400
transform 1 0 55888 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_491
timestamp 1669390400
transform 1 0 56336 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_495
timestamp 1669390400
transform 1 0 56784 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_503
timestamp 1669390400
transform 1 0 57680 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_507
timestamp 1669390400
transform 1 0 58128 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_5
timestamp 1669390400
transform 1 0 1904 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_9
timestamp 1669390400
transform 1 0 2352 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_47
timestamp 1669390400
transform 1 0 6608 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_55
timestamp 1669390400
transform 1 0 7504 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_59
timestamp 1669390400
transform 1 0 7952 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1669390400
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_73
timestamp 1669390400
transform 1 0 9520 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_80
timestamp 1669390400
transform 1 0 10304 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_84
timestamp 1669390400
transform 1 0 10752 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_94
timestamp 1669390400
transform 1 0 11872 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_96
timestamp 1669390400
transform 1 0 12096 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_99
timestamp 1669390400
transform 1 0 12432 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_106
timestamp 1669390400
transform 1 0 13216 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_114
timestamp 1669390400
transform 1 0 14112 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_116
timestamp 1669390400
transform 1 0 14336 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_119
timestamp 1669390400
transform 1 0 14672 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_131
timestamp 1669390400
transform 1 0 16016 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_137
timestamp 1669390400
transform 1 0 16688 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1669390400
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_144
timestamp 1669390400
transform 1 0 17472 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_150
timestamp 1669390400
transform 1 0 18144 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_156
timestamp 1669390400
transform 1 0 18816 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_160
timestamp 1669390400
transform 1 0 19264 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_164
timestamp 1669390400
transform 1 0 19712 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_174
timestamp 1669390400
transform 1 0 20832 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_178
timestamp 1669390400
transform 1 0 21280 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_181
timestamp 1669390400
transform 1 0 21616 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_191
timestamp 1669390400
transform 1 0 22736 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_201
timestamp 1669390400
transform 1 0 23856 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_205
timestamp 1669390400
transform 1 0 24304 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_209
timestamp 1669390400
transform 1 0 24752 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_215
timestamp 1669390400
transform 1 0 25424 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_221
timestamp 1669390400
transform 1 0 26096 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_225
timestamp 1669390400
transform 1 0 26544 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_229
timestamp 1669390400
transform 1 0 26992 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_233
timestamp 1669390400
transform 1 0 27440 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_239
timestamp 1669390400
transform 1 0 28112 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_243
timestamp 1669390400
transform 1 0 28560 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_247
timestamp 1669390400
transform 1 0 29008 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_257
timestamp 1669390400
transform 1 0 30128 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_265
timestamp 1669390400
transform 1 0 31024 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_268
timestamp 1669390400
transform 1 0 31360 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_286
timestamp 1669390400
transform 1 0 33376 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_288
timestamp 1669390400
transform 1 0 33600 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_294
timestamp 1669390400
transform 1 0 34272 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_302
timestamp 1669390400
transform 1 0 35168 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_310
timestamp 1669390400
transform 1 0 36064 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_312
timestamp 1669390400
transform 1 0 36288 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_319
timestamp 1669390400
transform 1 0 37072 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_327
timestamp 1669390400
transform 1 0 37968 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_331
timestamp 1669390400
transform 1 0 38416 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_335
timestamp 1669390400
transform 1 0 38864 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_343
timestamp 1669390400
transform 1 0 39760 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_347
timestamp 1669390400
transform 1 0 40208 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_351
timestamp 1669390400
transform 1 0 40656 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_354
timestamp 1669390400
transform 1 0 40992 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_357
timestamp 1669390400
transform 1 0 41328 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_371
timestamp 1669390400
transform 1 0 42896 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_375
timestamp 1669390400
transform 1 0 43344 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_381
timestamp 1669390400
transform 1 0 44016 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_400
timestamp 1669390400
transform 1 0 46144 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_414
timestamp 1669390400
transform 1 0 47712 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_422
timestamp 1669390400
transform 1 0 48608 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_47_428
timestamp 1669390400
transform 1 0 49280 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_492
timestamp 1669390400
transform 1 0 56448 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_496
timestamp 1669390400
transform 1 0 56896 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_499
timestamp 1669390400
transform 1 0 57232 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_507
timestamp 1669390400
transform 1 0 58128 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_2
timestamp 1669390400
transform 1 0 1568 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_12
timestamp 1669390400
transform 1 0 2688 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_20
timestamp 1669390400
transform 1 0 3584 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_26
timestamp 1669390400
transform 1 0 4256 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1669390400
transform 1 0 5152 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_37
timestamp 1669390400
transform 1 0 5488 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_43
timestamp 1669390400
transform 1 0 6160 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_71
timestamp 1669390400
transform 1 0 9296 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_91
timestamp 1669390400
transform 1 0 11536 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_98
timestamp 1669390400
transform 1 0 12320 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_102
timestamp 1669390400
transform 1 0 12768 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1669390400
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_108
timestamp 1669390400
transform 1 0 13440 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_123
timestamp 1669390400
transform 1 0 15120 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_127
timestamp 1669390400
transform 1 0 15568 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_131
timestamp 1669390400
transform 1 0 16016 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_148
timestamp 1669390400
transform 1 0 17920 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_158
timestamp 1669390400
transform 1 0 19040 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_162
timestamp 1669390400
transform 1 0 19488 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1669390400
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_179
timestamp 1669390400
transform 1 0 21392 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_188
timestamp 1669390400
transform 1 0 22400 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_190
timestamp 1669390400
transform 1 0 22624 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_207
timestamp 1669390400
transform 1 0 24528 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_211
timestamp 1669390400
transform 1 0 24976 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_220
timestamp 1669390400
transform 1 0 25984 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_224
timestamp 1669390400
transform 1 0 26432 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_228
timestamp 1669390400
transform 1 0 26880 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_231
timestamp 1669390400
transform 1 0 27216 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_237
timestamp 1669390400
transform 1 0 27888 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1669390400
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_250
timestamp 1669390400
transform 1 0 29344 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_259
timestamp 1669390400
transform 1 0 30352 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_263
timestamp 1669390400
transform 1 0 30800 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_267
timestamp 1669390400
transform 1 0 31248 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_271
timestamp 1669390400
transform 1 0 31696 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_273
timestamp 1669390400
transform 1 0 31920 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_279
timestamp 1669390400
transform 1 0 32592 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_283
timestamp 1669390400
transform 1 0 33040 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_299
timestamp 1669390400
transform 1 0 34832 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_303
timestamp 1669390400
transform 1 0 35280 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_306
timestamp 1669390400
transform 1 0 35616 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_310
timestamp 1669390400
transform 1 0 36064 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_313
timestamp 1669390400
transform 1 0 36400 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_317
timestamp 1669390400
transform 1 0 36848 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_321
timestamp 1669390400
transform 1 0 37296 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_329
timestamp 1669390400
transform 1 0 38192 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_333
timestamp 1669390400
transform 1 0 38640 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_346
timestamp 1669390400
transform 1 0 40096 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_353
timestamp 1669390400
transform 1 0 40880 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_369
timestamp 1669390400
transform 1 0 42672 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_375
timestamp 1669390400
transform 1 0 43344 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_385
timestamp 1669390400
transform 1 0 44464 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1669390400
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_392
timestamp 1669390400
transform 1 0 45248 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_401
timestamp 1669390400
transform 1 0 46256 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_433
timestamp 1669390400
transform 1 0 49840 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_449
timestamp 1669390400
transform 1 0 51632 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_457
timestamp 1669390400
transform 1 0 52528 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_463
timestamp 1669390400
transform 1 0 53200 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_471
timestamp 1669390400
transform 1 0 54096 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_475
timestamp 1669390400
transform 1 0 54544 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_491
timestamp 1669390400
transform 1 0 56336 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_507
timestamp 1669390400
transform 1 0 58128 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_2
timestamp 1669390400
transform 1 0 1568 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_6
timestamp 1669390400
transform 1 0 2016 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_10
timestamp 1669390400
transform 1 0 2464 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_18
timestamp 1669390400
transform 1 0 3360 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_20
timestamp 1669390400
transform 1 0 3584 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_27
timestamp 1669390400
transform 1 0 4368 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_46
timestamp 1669390400
transform 1 0 6496 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_56
timestamp 1669390400
transform 1 0 7616 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_60
timestamp 1669390400
transform 1 0 8064 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_67
timestamp 1669390400
transform 1 0 8848 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_73
timestamp 1669390400
transform 1 0 9520 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_75
timestamp 1669390400
transform 1 0 9744 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_78
timestamp 1669390400
transform 1 0 10080 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_88
timestamp 1669390400
transform 1 0 11200 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_92
timestamp 1669390400
transform 1 0 11648 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_100
timestamp 1669390400
transform 1 0 12544 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_108
timestamp 1669390400
transform 1 0 13440 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_118
timestamp 1669390400
transform 1 0 14560 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_122
timestamp 1669390400
transform 1 0 15008 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_125
timestamp 1669390400
transform 1 0 15344 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_129
timestamp 1669390400
transform 1 0 15792 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_133
timestamp 1669390400
transform 1 0 16240 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1669390400
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_144
timestamp 1669390400
transform 1 0 17472 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_163
timestamp 1669390400
transform 1 0 19600 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_167
timestamp 1669390400
transform 1 0 20048 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_171
timestamp 1669390400
transform 1 0 20496 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_175
timestamp 1669390400
transform 1 0 20944 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_179
timestamp 1669390400
transform 1 0 21392 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_183
timestamp 1669390400
transform 1 0 21840 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_187
timestamp 1669390400
transform 1 0 22288 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_191
timestamp 1669390400
transform 1 0 22736 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_201
timestamp 1669390400
transform 1 0 23856 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_205
timestamp 1669390400
transform 1 0 24304 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_210
timestamp 1669390400
transform 1 0 24864 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1669390400
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_215
timestamp 1669390400
transform 1 0 25424 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_221
timestamp 1669390400
transform 1 0 26096 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_231
timestamp 1669390400
transform 1 0 27216 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_239
timestamp 1669390400
transform 1 0 28112 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_253
timestamp 1669390400
transform 1 0 29680 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_261
timestamp 1669390400
transform 1 0 30576 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_267
timestamp 1669390400
transform 1 0 31248 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_279
timestamp 1669390400
transform 1 0 32592 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1669390400
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_286
timestamp 1669390400
transform 1 0 33376 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_296
timestamp 1669390400
transform 1 0 34496 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_304
timestamp 1669390400
transform 1 0 35392 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_311
timestamp 1669390400
transform 1 0 36176 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_319
timestamp 1669390400
transform 1 0 37072 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_327
timestamp 1669390400
transform 1 0 37968 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_331
timestamp 1669390400
transform 1 0 38416 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_344
timestamp 1669390400
transform 1 0 39872 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_354
timestamp 1669390400
transform 1 0 40992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_357
timestamp 1669390400
transform 1 0 41328 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_360
timestamp 1669390400
transform 1 0 41664 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_386
timestamp 1669390400
transform 1 0 44576 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_418
timestamp 1669390400
transform 1 0 48160 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_49_428
timestamp 1669390400
transform 1 0 49280 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_492
timestamp 1669390400
transform 1 0 56448 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_496
timestamp 1669390400
transform 1 0 56896 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_499
timestamp 1669390400
transform 1 0 57232 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_507
timestamp 1669390400
transform 1 0 58128 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_2
timestamp 1669390400
transform 1 0 1568 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_14
timestamp 1669390400
transform 1 0 2912 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_31
timestamp 1669390400
transform 1 0 4816 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_37
timestamp 1669390400
transform 1 0 5488 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_40
timestamp 1669390400
transform 1 0 5824 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_51
timestamp 1669390400
transform 1 0 7056 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_59
timestamp 1669390400
transform 1 0 7952 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_63
timestamp 1669390400
transform 1 0 8400 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_66
timestamp 1669390400
transform 1 0 8736 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_70
timestamp 1669390400
transform 1 0 9184 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_78
timestamp 1669390400
transform 1 0 10080 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_103
timestamp 1669390400
transform 1 0 12880 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1669390400
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_108
timestamp 1669390400
transform 1 0 13440 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_119
timestamp 1669390400
transform 1 0 14672 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_123
timestamp 1669390400
transform 1 0 15120 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_126
timestamp 1669390400
transform 1 0 15456 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_135
timestamp 1669390400
transform 1 0 16464 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_137
timestamp 1669390400
transform 1 0 16688 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_140
timestamp 1669390400
transform 1 0 17024 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_144
timestamp 1669390400
transform 1 0 17472 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_154
timestamp 1669390400
transform 1 0 18592 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_168
timestamp 1669390400
transform 1 0 20160 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_172
timestamp 1669390400
transform 1 0 20608 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1669390400
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_179
timestamp 1669390400
transform 1 0 21392 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_183
timestamp 1669390400
transform 1 0 21840 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_195
timestamp 1669390400
transform 1 0 23184 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_197
timestamp 1669390400
transform 1 0 23408 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_204
timestamp 1669390400
transform 1 0 24192 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_208
timestamp 1669390400
transform 1 0 24640 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_212
timestamp 1669390400
transform 1 0 25088 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_215
timestamp 1669390400
transform 1 0 25424 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_227
timestamp 1669390400
transform 1 0 26768 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_233
timestamp 1669390400
transform 1 0 27440 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_237
timestamp 1669390400
transform 1 0 27888 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_244
timestamp 1669390400
transform 1 0 28672 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_250
timestamp 1669390400
transform 1 0 29344 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_253
timestamp 1669390400
transform 1 0 29680 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_257
timestamp 1669390400
transform 1 0 30128 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_265
timestamp 1669390400
transform 1 0 31024 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_286
timestamp 1669390400
transform 1 0 33376 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_302
timestamp 1669390400
transform 1 0 35168 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_311
timestamp 1669390400
transform 1 0 36176 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_321
timestamp 1669390400
transform 1 0 37296 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_323
timestamp 1669390400
transform 1 0 37520 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_330
timestamp 1669390400
transform 1 0 38304 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_334
timestamp 1669390400
transform 1 0 38752 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_338
timestamp 1669390400
transform 1 0 39200 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_340
timestamp 1669390400
transform 1 0 39424 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_351
timestamp 1669390400
transform 1 0 40656 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_355
timestamp 1669390400
transform 1 0 41104 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_371
timestamp 1669390400
transform 1 0 42896 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_375
timestamp 1669390400
transform 1 0 43344 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_385
timestamp 1669390400
transform 1 0 44464 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_389
timestamp 1669390400
transform 1 0 44912 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_50_392
timestamp 1669390400
transform 1 0 45248 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_456
timestamp 1669390400
transform 1 0 52416 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_460
timestamp 1669390400
transform 1 0 52864 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_463
timestamp 1669390400
transform 1 0 53200 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_495
timestamp 1669390400
transform 1 0 56784 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_503
timestamp 1669390400
transform 1 0 57680 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_507
timestamp 1669390400
transform 1 0 58128 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_2
timestamp 1669390400
transform 1 0 1568 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_6
timestamp 1669390400
transform 1 0 2016 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_10
timestamp 1669390400
transform 1 0 2464 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_14
timestamp 1669390400
transform 1 0 2912 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_22
timestamp 1669390400
transform 1 0 3808 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_30
timestamp 1669390400
transform 1 0 4704 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_32
timestamp 1669390400
transform 1 0 4928 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_35
timestamp 1669390400
transform 1 0 5264 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_39
timestamp 1669390400
transform 1 0 5712 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_43
timestamp 1669390400
transform 1 0 6160 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_47
timestamp 1669390400
transform 1 0 6608 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_51
timestamp 1669390400
transform 1 0 7056 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_61
timestamp 1669390400
transform 1 0 8176 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_63
timestamp 1669390400
transform 1 0 8400 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_66
timestamp 1669390400
transform 1 0 8736 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1669390400
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_73
timestamp 1669390400
transform 1 0 9520 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_77
timestamp 1669390400
transform 1 0 9968 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_81
timestamp 1669390400
transform 1 0 10416 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_89
timestamp 1669390400
transform 1 0 11312 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_103
timestamp 1669390400
transform 1 0 12880 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_105
timestamp 1669390400
transform 1 0 13104 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_116
timestamp 1669390400
transform 1 0 14336 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_126
timestamp 1669390400
transform 1 0 15456 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_130
timestamp 1669390400
transform 1 0 15904 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1669390400
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_144
timestamp 1669390400
transform 1 0 17472 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_147
timestamp 1669390400
transform 1 0 17808 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_151
timestamp 1669390400
transform 1 0 18256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_155
timestamp 1669390400
transform 1 0 18704 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_158
timestamp 1669390400
transform 1 0 19040 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_170
timestamp 1669390400
transform 1 0 20384 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_174
timestamp 1669390400
transform 1 0 20832 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_178
timestamp 1669390400
transform 1 0 21280 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_182
timestamp 1669390400
transform 1 0 21728 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_186
timestamp 1669390400
transform 1 0 22176 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_206
timestamp 1669390400
transform 1 0 24416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_212
timestamp 1669390400
transform 1 0 25088 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_215
timestamp 1669390400
transform 1 0 25424 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_225
timestamp 1669390400
transform 1 0 26544 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_229
timestamp 1669390400
transform 1 0 26992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_235
timestamp 1669390400
transform 1 0 27664 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_245
timestamp 1669390400
transform 1 0 28784 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_255
timestamp 1669390400
transform 1 0 29904 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_259
timestamp 1669390400
transform 1 0 30352 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_263
timestamp 1669390400
transform 1 0 30800 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_267
timestamp 1669390400
transform 1 0 31248 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_271
timestamp 1669390400
transform 1 0 31696 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_281
timestamp 1669390400
transform 1 0 32816 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_283
timestamp 1669390400
transform 1 0 33040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_286
timestamp 1669390400
transform 1 0 33376 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_289
timestamp 1669390400
transform 1 0 33712 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_303
timestamp 1669390400
transform 1 0 35280 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_313
timestamp 1669390400
transform 1 0 36400 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_317
timestamp 1669390400
transform 1 0 36848 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_321
timestamp 1669390400
transform 1 0 37296 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_329
timestamp 1669390400
transform 1 0 38192 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_342
timestamp 1669390400
transform 1 0 39648 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_346
timestamp 1669390400
transform 1 0 40096 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_350
timestamp 1669390400
transform 1 0 40544 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1669390400
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_357
timestamp 1669390400
transform 1 0 41328 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_363
timestamp 1669390400
transform 1 0 42000 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_375
timestamp 1669390400
transform 1 0 43344 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_385
timestamp 1669390400
transform 1 0 44464 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_395
timestamp 1669390400
transform 1 0 45584 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_403
timestamp 1669390400
transform 1 0 46480 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_419
timestamp 1669390400
transform 1 0 48272 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_423
timestamp 1669390400
transform 1 0 48720 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_425
timestamp 1669390400
transform 1 0 48944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_51_428
timestamp 1669390400
transform 1 0 49280 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_492
timestamp 1669390400
transform 1 0 56448 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_496
timestamp 1669390400
transform 1 0 56896 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_499
timestamp 1669390400
transform 1 0 57232 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_507
timestamp 1669390400
transform 1 0 58128 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_2
timestamp 1669390400
transform 1 0 1568 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_4
timestamp 1669390400
transform 1 0 1792 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_7
timestamp 1669390400
transform 1 0 2128 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_11
timestamp 1669390400
transform 1 0 2576 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_19
timestamp 1669390400
transform 1 0 3472 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_27
timestamp 1669390400
transform 1 0 4368 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_31
timestamp 1669390400
transform 1 0 4816 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1669390400
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_37
timestamp 1669390400
transform 1 0 5488 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_45
timestamp 1669390400
transform 1 0 6384 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_57
timestamp 1669390400
transform 1 0 7728 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_82
timestamp 1669390400
transform 1 0 10528 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_86
timestamp 1669390400
transform 1 0 10976 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_90
timestamp 1669390400
transform 1 0 11424 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_104
timestamp 1669390400
transform 1 0 12992 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_108
timestamp 1669390400
transform 1 0 13440 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_112
timestamp 1669390400
transform 1 0 13888 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_116
timestamp 1669390400
transform 1 0 14336 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_120
timestamp 1669390400
transform 1 0 14784 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_130
timestamp 1669390400
transform 1 0 15904 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_139
timestamp 1669390400
transform 1 0 16912 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_146
timestamp 1669390400
transform 1 0 17696 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_152
timestamp 1669390400
transform 1 0 18368 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_162
timestamp 1669390400
transform 1 0 19488 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_170
timestamp 1669390400
transform 1 0 20384 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_174
timestamp 1669390400
transform 1 0 20832 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1669390400
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_179
timestamp 1669390400
transform 1 0 21392 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_191
timestamp 1669390400
transform 1 0 22736 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_201
timestamp 1669390400
transform 1 0 23856 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_205
timestamp 1669390400
transform 1 0 24304 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_209
timestamp 1669390400
transform 1 0 24752 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_213
timestamp 1669390400
transform 1 0 25200 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_216
timestamp 1669390400
transform 1 0 25536 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_220
timestamp 1669390400
transform 1 0 25984 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_224
timestamp 1669390400
transform 1 0 26432 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_228
timestamp 1669390400
transform 1 0 26880 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_232
timestamp 1669390400
transform 1 0 27328 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1669390400
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_250
timestamp 1669390400
transform 1 0 29344 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_256
timestamp 1669390400
transform 1 0 30016 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_260
timestamp 1669390400
transform 1 0 30464 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_264
timestamp 1669390400
transform 1 0 30912 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_268
timestamp 1669390400
transform 1 0 31360 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_285
timestamp 1669390400
transform 1 0 33264 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_289
timestamp 1669390400
transform 1 0 33712 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_297
timestamp 1669390400
transform 1 0 34608 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_301
timestamp 1669390400
transform 1 0 35056 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_303
timestamp 1669390400
transform 1 0 35280 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_312
timestamp 1669390400
transform 1 0 36288 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_318
timestamp 1669390400
transform 1 0 36960 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_321
timestamp 1669390400
transform 1 0 37296 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_337
timestamp 1669390400
transform 1 0 39088 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_363
timestamp 1669390400
transform 1 0 42000 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_365
timestamp 1669390400
transform 1 0 42224 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_368
timestamp 1669390400
transform 1 0 42560 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_377
timestamp 1669390400
transform 1 0 43568 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_389
timestamp 1669390400
transform 1 0 44912 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_392
timestamp 1669390400
transform 1 0 45248 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_399
timestamp 1669390400
transform 1 0 46032 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_431
timestamp 1669390400
transform 1 0 49616 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_447
timestamp 1669390400
transform 1 0 51408 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_455
timestamp 1669390400
transform 1 0 52304 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_459
timestamp 1669390400
transform 1 0 52752 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_463
timestamp 1669390400
transform 1 0 53200 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_495
timestamp 1669390400
transform 1 0 56784 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_503
timestamp 1669390400
transform 1 0 57680 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_507
timestamp 1669390400
transform 1 0 58128 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_2
timestamp 1669390400
transform 1 0 1568 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_17
timestamp 1669390400
transform 1 0 3248 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_21
timestamp 1669390400
transform 1 0 3696 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_28
timestamp 1669390400
transform 1 0 4480 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_32
timestamp 1669390400
transform 1 0 4928 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_40
timestamp 1669390400
transform 1 0 5824 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_42
timestamp 1669390400
transform 1 0 6048 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_45
timestamp 1669390400
transform 1 0 6384 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_57
timestamp 1669390400
transform 1 0 7728 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_59
timestamp 1669390400
transform 1 0 7952 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_69
timestamp 1669390400
transform 1 0 9072 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_73
timestamp 1669390400
transform 1 0 9520 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_87
timestamp 1669390400
transform 1 0 11088 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_97
timestamp 1669390400
transform 1 0 12208 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_99
timestamp 1669390400
transform 1 0 12432 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_102
timestamp 1669390400
transform 1 0 12768 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_111
timestamp 1669390400
transform 1 0 13776 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_118
timestamp 1669390400
transform 1 0 14560 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_122
timestamp 1669390400
transform 1 0 15008 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_125
timestamp 1669390400
transform 1 0 15344 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_129
timestamp 1669390400
transform 1 0 15792 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_133
timestamp 1669390400
transform 1 0 16240 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_137
timestamp 1669390400
transform 1 0 16688 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1669390400
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_144
timestamp 1669390400
transform 1 0 17472 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_150
timestamp 1669390400
transform 1 0 18144 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_154
timestamp 1669390400
transform 1 0 18592 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_160
timestamp 1669390400
transform 1 0 19264 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_175
timestamp 1669390400
transform 1 0 20944 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_186
timestamp 1669390400
transform 1 0 22176 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_196
timestamp 1669390400
transform 1 0 23296 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_198
timestamp 1669390400
transform 1 0 23520 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_201
timestamp 1669390400
transform 1 0 23856 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_211
timestamp 1669390400
transform 1 0 24976 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_215
timestamp 1669390400
transform 1 0 25424 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_224
timestamp 1669390400
transform 1 0 26432 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_234
timestamp 1669390400
transform 1 0 27552 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_244
timestamp 1669390400
transform 1 0 28672 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_248
timestamp 1669390400
transform 1 0 29120 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_262
timestamp 1669390400
transform 1 0 30688 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1669390400
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_286
timestamp 1669390400
transform 1 0 33376 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_290
timestamp 1669390400
transform 1 0 33824 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_302
timestamp 1669390400
transform 1 0 35168 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_312
timestamp 1669390400
transform 1 0 36288 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_314
timestamp 1669390400
transform 1 0 36512 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_322
timestamp 1669390400
transform 1 0 37408 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_326
timestamp 1669390400
transform 1 0 37856 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_330
timestamp 1669390400
transform 1 0 38304 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_338
timestamp 1669390400
transform 1 0 39200 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_347
timestamp 1669390400
transform 1 0 40208 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_351
timestamp 1669390400
transform 1 0 40656 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_357
timestamp 1669390400
transform 1 0 41328 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_365
timestamp 1669390400
transform 1 0 42224 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_367
timestamp 1669390400
transform 1 0 42448 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_374
timestamp 1669390400
transform 1 0 43232 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_378
timestamp 1669390400
transform 1 0 43680 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_387
timestamp 1669390400
transform 1 0 44688 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_419
timestamp 1669390400
transform 1 0 48272 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_423
timestamp 1669390400
transform 1 0 48720 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_425
timestamp 1669390400
transform 1 0 48944 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_53_428
timestamp 1669390400
transform 1 0 49280 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_492
timestamp 1669390400
transform 1 0 56448 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_496
timestamp 1669390400
transform 1 0 56896 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_499
timestamp 1669390400
transform 1 0 57232 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_507
timestamp 1669390400
transform 1 0 58128 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_2
timestamp 1669390400
transform 1 0 1568 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_6
timestamp 1669390400
transform 1 0 2016 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_14
timestamp 1669390400
transform 1 0 2912 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_24
timestamp 1669390400
transform 1 0 4032 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1669390400
transform 1 0 5152 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_37
timestamp 1669390400
transform 1 0 5488 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_39
timestamp 1669390400
transform 1 0 5712 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_42
timestamp 1669390400
transform 1 0 6048 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_52
timestamp 1669390400
transform 1 0 7168 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_56
timestamp 1669390400
transform 1 0 7616 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_81
timestamp 1669390400
transform 1 0 10416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_85
timestamp 1669390400
transform 1 0 10864 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_91
timestamp 1669390400
transform 1 0 11536 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_95
timestamp 1669390400
transform 1 0 11984 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_98
timestamp 1669390400
transform 1 0 12320 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1669390400
transform 1 0 13104 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_108
timestamp 1669390400
transform 1 0 13440 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_119
timestamp 1669390400
transform 1 0 14672 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_121
timestamp 1669390400
transform 1 0 14896 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_124
timestamp 1669390400
transform 1 0 15232 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_134
timestamp 1669390400
transform 1 0 16352 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_142
timestamp 1669390400
transform 1 0 17248 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_146
timestamp 1669390400
transform 1 0 17696 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_150
timestamp 1669390400
transform 1 0 18144 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_154
timestamp 1669390400
transform 1 0 18592 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_158
timestamp 1669390400
transform 1 0 19040 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_160
timestamp 1669390400
transform 1 0 19264 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_167
timestamp 1669390400
transform 1 0 20048 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_175
timestamp 1669390400
transform 1 0 20944 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_179
timestamp 1669390400
transform 1 0 21392 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_185
timestamp 1669390400
transform 1 0 22064 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_193
timestamp 1669390400
transform 1 0 22960 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_232
timestamp 1669390400
transform 1 0 27328 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_236
timestamp 1669390400
transform 1 0 27776 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_242
timestamp 1669390400
transform 1 0 28448 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_246
timestamp 1669390400
transform 1 0 28896 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_250
timestamp 1669390400
transform 1 0 29344 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_253
timestamp 1669390400
transform 1 0 29680 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_257
timestamp 1669390400
transform 1 0 30128 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_260
timestamp 1669390400
transform 1 0 30464 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_264
timestamp 1669390400
transform 1 0 30912 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_274
timestamp 1669390400
transform 1 0 32032 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_278
timestamp 1669390400
transform 1 0 32480 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_284
timestamp 1669390400
transform 1 0 33152 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_291
timestamp 1669390400
transform 1 0 33936 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_301
timestamp 1669390400
transform 1 0 35056 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_305
timestamp 1669390400
transform 1 0 35504 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_309
timestamp 1669390400
transform 1 0 35952 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_311
timestamp 1669390400
transform 1 0 36176 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_317
timestamp 1669390400
transform 1 0 36848 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_321
timestamp 1669390400
transform 1 0 37296 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_324
timestamp 1669390400
transform 1 0 37632 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_328
timestamp 1669390400
transform 1 0 38080 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_332
timestamp 1669390400
transform 1 0 38528 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_338
timestamp 1669390400
transform 1 0 39200 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_348
timestamp 1669390400
transform 1 0 40320 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_386
timestamp 1669390400
transform 1 0 44576 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_54_392
timestamp 1669390400
transform 1 0 45248 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_456
timestamp 1669390400
transform 1 0 52416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_460
timestamp 1669390400
transform 1 0 52864 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_463
timestamp 1669390400
transform 1 0 53200 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_479
timestamp 1669390400
transform 1 0 54992 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_487
timestamp 1669390400
transform 1 0 55888 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_491
timestamp 1669390400
transform 1 0 56336 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_495
timestamp 1669390400
transform 1 0 56784 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_503
timestamp 1669390400
transform 1 0 57680 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_507
timestamp 1669390400
transform 1 0 58128 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_2
timestamp 1669390400
transform 1 0 1568 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_10
timestamp 1669390400
transform 1 0 2464 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_18
timestamp 1669390400
transform 1 0 3360 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_28
timestamp 1669390400
transform 1 0 4480 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_34
timestamp 1669390400
transform 1 0 5152 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_38
timestamp 1669390400
transform 1 0 5600 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_42
timestamp 1669390400
transform 1 0 6048 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_49
timestamp 1669390400
transform 1 0 6832 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_53
timestamp 1669390400
transform 1 0 7280 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_56
timestamp 1669390400
transform 1 0 7616 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_63
timestamp 1669390400
transform 1 0 8400 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_70
timestamp 1669390400
transform 1 0 9184 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_73
timestamp 1669390400
transform 1 0 9520 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_81
timestamp 1669390400
transform 1 0 10416 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_85
timestamp 1669390400
transform 1 0 10864 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_89
timestamp 1669390400
transform 1 0 11312 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_93
timestamp 1669390400
transform 1 0 11760 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_97
timestamp 1669390400
transform 1 0 12208 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_101
timestamp 1669390400
transform 1 0 12656 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_105
timestamp 1669390400
transform 1 0 13104 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_114
timestamp 1669390400
transform 1 0 14112 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_116
timestamp 1669390400
transform 1 0 14336 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_119
timestamp 1669390400
transform 1 0 14672 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_123
timestamp 1669390400
transform 1 0 15120 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_127
timestamp 1669390400
transform 1 0 15568 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_131
timestamp 1669390400
transform 1 0 16016 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_141
timestamp 1669390400
transform 1 0 17136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_144
timestamp 1669390400
transform 1 0 17472 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_156
timestamp 1669390400
transform 1 0 18816 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_160
timestamp 1669390400
transform 1 0 19264 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_172
timestamp 1669390400
transform 1 0 20608 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_174
timestamp 1669390400
transform 1 0 20832 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_177
timestamp 1669390400
transform 1 0 21168 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_181
timestamp 1669390400
transform 1 0 21616 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_187
timestamp 1669390400
transform 1 0 22288 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_191
timestamp 1669390400
transform 1 0 22736 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_199
timestamp 1669390400
transform 1 0 23632 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_203
timestamp 1669390400
transform 1 0 24080 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_207
timestamp 1669390400
transform 1 0 24528 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_211
timestamp 1669390400
transform 1 0 24976 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_215
timestamp 1669390400
transform 1 0 25424 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_219
timestamp 1669390400
transform 1 0 25872 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_223
timestamp 1669390400
transform 1 0 26320 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_235
timestamp 1669390400
transform 1 0 27664 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_245
timestamp 1669390400
transform 1 0 28784 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_260
timestamp 1669390400
transform 1 0 30464 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_264
timestamp 1669390400
transform 1 0 30912 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_268
timestamp 1669390400
transform 1 0 31360 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_272
timestamp 1669390400
transform 1 0 31808 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_276
timestamp 1669390400
transform 1 0 32256 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_280
timestamp 1669390400
transform 1 0 32704 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_286
timestamp 1669390400
transform 1 0 33376 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_289
timestamp 1669390400
transform 1 0 33712 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_293
timestamp 1669390400
transform 1 0 34160 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_297
timestamp 1669390400
transform 1 0 34608 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_301
timestamp 1669390400
transform 1 0 35056 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_305
timestamp 1669390400
transform 1 0 35504 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_309
timestamp 1669390400
transform 1 0 35952 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_313
timestamp 1669390400
transform 1 0 36400 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_316
timestamp 1669390400
transform 1 0 36736 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_329
timestamp 1669390400
transform 1 0 38192 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_337
timestamp 1669390400
transform 1 0 39088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_340
timestamp 1669390400
transform 1 0 39424 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_352
timestamp 1669390400
transform 1 0 40768 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1669390400
transform 1 0 40992 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_357
timestamp 1669390400
transform 1 0 41328 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_373
timestamp 1669390400
transform 1 0 43120 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_389
timestamp 1669390400
transform 1 0 44912 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_421
timestamp 1669390400
transform 1 0 48496 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_425
timestamp 1669390400
transform 1 0 48944 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_55_428
timestamp 1669390400
transform 1 0 49280 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_460
timestamp 1669390400
transform 1 0 52864 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_476
timestamp 1669390400
transform 1 0 54656 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_491
timestamp 1669390400
transform 1 0 56336 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_495
timestamp 1669390400
transform 1 0 56784 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_499
timestamp 1669390400
transform 1 0 57232 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_507
timestamp 1669390400
transform 1 0 58128 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_2
timestamp 1669390400
transform 1 0 1568 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_4
timestamp 1669390400
transform 1 0 1792 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_11
timestamp 1669390400
transform 1 0 2576 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_23
timestamp 1669390400
transform 1 0 3920 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_27
timestamp 1669390400
transform 1 0 4368 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_30
timestamp 1669390400
transform 1 0 4704 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1669390400
transform 1 0 5152 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_37
timestamp 1669390400
transform 1 0 5488 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_40
timestamp 1669390400
transform 1 0 5824 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_44
timestamp 1669390400
transform 1 0 6272 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_52
timestamp 1669390400
transform 1 0 7168 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_56
timestamp 1669390400
transform 1 0 7616 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_59
timestamp 1669390400
transform 1 0 7952 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_63
timestamp 1669390400
transform 1 0 8400 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_73
timestamp 1669390400
transform 1 0 9520 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_75
timestamp 1669390400
transform 1 0 9744 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_78
timestamp 1669390400
transform 1 0 10080 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_82
timestamp 1669390400
transform 1 0 10528 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_90
timestamp 1669390400
transform 1 0 11424 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_94
timestamp 1669390400
transform 1 0 11872 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_97
timestamp 1669390400
transform 1 0 12208 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1669390400
transform 1 0 13104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_108
timestamp 1669390400
transform 1 0 13440 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_110
timestamp 1669390400
transform 1 0 13664 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_119
timestamp 1669390400
transform 1 0 14672 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_126
timestamp 1669390400
transform 1 0 15456 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_128
timestamp 1669390400
transform 1 0 15680 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_152
timestamp 1669390400
transform 1 0 18368 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_156
timestamp 1669390400
transform 1 0 18816 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_159
timestamp 1669390400
transform 1 0 19152 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_173
timestamp 1669390400
transform 1 0 20720 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_179
timestamp 1669390400
transform 1 0 21392 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_186
timestamp 1669390400
transform 1 0 22176 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_200
timestamp 1669390400
transform 1 0 23744 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_208
timestamp 1669390400
transform 1 0 24640 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_210
timestamp 1669390400
transform 1 0 24864 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_213
timestamp 1669390400
transform 1 0 25200 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_217
timestamp 1669390400
transform 1 0 25648 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_237
timestamp 1669390400
transform 1 0 27888 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_246
timestamp 1669390400
transform 1 0 28896 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_250
timestamp 1669390400
transform 1 0 29344 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_267
timestamp 1669390400
transform 1 0 31248 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_271
timestamp 1669390400
transform 1 0 31696 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_275
timestamp 1669390400
transform 1 0 32144 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_279
timestamp 1669390400
transform 1 0 32592 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_286
timestamp 1669390400
transform 1 0 33376 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_296
timestamp 1669390400
transform 1 0 34496 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_298
timestamp 1669390400
transform 1 0 34720 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_307
timestamp 1669390400
transform 1 0 35728 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_315
timestamp 1669390400
transform 1 0 36624 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_321
timestamp 1669390400
transform 1 0 37296 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_334
timestamp 1669390400
transform 1 0 38752 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_338
timestamp 1669390400
transform 1 0 39200 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_344
timestamp 1669390400
transform 1 0 39872 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_364
timestamp 1669390400
transform 1 0 42112 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_372
timestamp 1669390400
transform 1 0 43008 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_386
timestamp 1669390400
transform 1 0 44576 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_392
timestamp 1669390400
transform 1 0 45248 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_401
timestamp 1669390400
transform 1 0 46256 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_433
timestamp 1669390400
transform 1 0 49840 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_449
timestamp 1669390400
transform 1 0 51632 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_457
timestamp 1669390400
transform 1 0 52528 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_463
timestamp 1669390400
transform 1 0 53200 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_495
timestamp 1669390400
transform 1 0 56784 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_503
timestamp 1669390400
transform 1 0 57680 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_507
timestamp 1669390400
transform 1 0 58128 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_2
timestamp 1669390400
transform 1 0 1568 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_6
timestamp 1669390400
transform 1 0 2016 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_10
timestamp 1669390400
transform 1 0 2464 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_18
timestamp 1669390400
transform 1 0 3360 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_28
timestamp 1669390400
transform 1 0 4480 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_38
timestamp 1669390400
transform 1 0 5600 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_42
timestamp 1669390400
transform 1 0 6048 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_51
timestamp 1669390400
transform 1 0 7056 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_59
timestamp 1669390400
transform 1 0 7952 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_63
timestamp 1669390400
transform 1 0 8400 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_70
timestamp 1669390400
transform 1 0 9184 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_73
timestamp 1669390400
transform 1 0 9520 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_75
timestamp 1669390400
transform 1 0 9744 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_82
timestamp 1669390400
transform 1 0 10528 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_94
timestamp 1669390400
transform 1 0 11872 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_98
timestamp 1669390400
transform 1 0 12320 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_108
timestamp 1669390400
transform 1 0 13440 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_133
timestamp 1669390400
transform 1 0 16240 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_141
timestamp 1669390400
transform 1 0 17136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_144
timestamp 1669390400
transform 1 0 17472 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_162
timestamp 1669390400
transform 1 0 19488 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_170
timestamp 1669390400
transform 1 0 20384 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_174
timestamp 1669390400
transform 1 0 20832 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_180
timestamp 1669390400
transform 1 0 21504 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_184
timestamp 1669390400
transform 1 0 21952 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_188
timestamp 1669390400
transform 1 0 22400 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_204
timestamp 1669390400
transform 1 0 24192 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1669390400
transform 1 0 25088 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_215
timestamp 1669390400
transform 1 0 25424 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_218
timestamp 1669390400
transform 1 0 25760 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_222
timestamp 1669390400
transform 1 0 26208 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_234
timestamp 1669390400
transform 1 0 27552 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_238
timestamp 1669390400
transform 1 0 28000 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_242
timestamp 1669390400
transform 1 0 28448 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_245
timestamp 1669390400
transform 1 0 28784 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_249
timestamp 1669390400
transform 1 0 29232 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_251
timestamp 1669390400
transform 1 0 29456 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_260
timestamp 1669390400
transform 1 0 30464 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_264
timestamp 1669390400
transform 1 0 30912 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_268
timestamp 1669390400
transform 1 0 31360 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_270
timestamp 1669390400
transform 1 0 31584 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_273
timestamp 1669390400
transform 1 0 31920 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_283
timestamp 1669390400
transform 1 0 33040 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_286
timestamp 1669390400
transform 1 0 33376 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_297
timestamp 1669390400
transform 1 0 34608 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_301
timestamp 1669390400
transform 1 0 35056 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_305
timestamp 1669390400
transform 1 0 35504 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_307
timestamp 1669390400
transform 1 0 35728 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_310
timestamp 1669390400
transform 1 0 36064 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_320
timestamp 1669390400
transform 1 0 37184 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_333
timestamp 1669390400
transform 1 0 38640 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_337
timestamp 1669390400
transform 1 0 39088 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_341
timestamp 1669390400
transform 1 0 39536 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_350
timestamp 1669390400
transform 1 0 40544 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_354
timestamp 1669390400
transform 1 0 40992 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_357
timestamp 1669390400
transform 1 0 41328 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_366
timestamp 1669390400
transform 1 0 42336 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_380
timestamp 1669390400
transform 1 0 43904 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_388
timestamp 1669390400
transform 1 0 44800 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_396
timestamp 1669390400
transform 1 0 45696 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_412
timestamp 1669390400
transform 1 0 47488 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_420
timestamp 1669390400
transform 1 0 48384 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_424
timestamp 1669390400
transform 1 0 48832 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_57_428
timestamp 1669390400
transform 1 0 49280 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_492
timestamp 1669390400
transform 1 0 56448 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_496
timestamp 1669390400
transform 1 0 56896 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_499
timestamp 1669390400
transform 1 0 57232 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_507
timestamp 1669390400
transform 1 0 58128 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_2
timestamp 1669390400
transform 1 0 1568 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_9
timestamp 1669390400
transform 1 0 2352 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_17
timestamp 1669390400
transform 1 0 3248 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_27
timestamp 1669390400
transform 1 0 4368 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1669390400
transform 1 0 5152 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_37
timestamp 1669390400
transform 1 0 5488 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_43
timestamp 1669390400
transform 1 0 6160 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_64
timestamp 1669390400
transform 1 0 8512 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_66
timestamp 1669390400
transform 1 0 8736 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_69
timestamp 1669390400
transform 1 0 9072 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_77
timestamp 1669390400
transform 1 0 9968 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_87
timestamp 1669390400
transform 1 0 11088 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_94
timestamp 1669390400
transform 1 0 11872 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_98
timestamp 1669390400
transform 1 0 12320 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_102
timestamp 1669390400
transform 1 0 12768 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1669390400
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_108
timestamp 1669390400
transform 1 0 13440 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_117
timestamp 1669390400
transform 1 0 14448 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_121
timestamp 1669390400
transform 1 0 14896 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_124
timestamp 1669390400
transform 1 0 15232 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_128
timestamp 1669390400
transform 1 0 15680 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_130
timestamp 1669390400
transform 1 0 15904 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_148
timestamp 1669390400
transform 1 0 17920 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_160
timestamp 1669390400
transform 1 0 19264 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_162
timestamp 1669390400
transform 1 0 19488 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_171
timestamp 1669390400
transform 1 0 20496 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_175
timestamp 1669390400
transform 1 0 20944 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_179
timestamp 1669390400
transform 1 0 21392 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_183
timestamp 1669390400
transform 1 0 21840 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_187
timestamp 1669390400
transform 1 0 22288 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_191
timestamp 1669390400
transform 1 0 22736 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_201
timestamp 1669390400
transform 1 0 23856 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_205
timestamp 1669390400
transform 1 0 24304 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_209
timestamp 1669390400
transform 1 0 24752 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_213
timestamp 1669390400
transform 1 0 25200 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_217
timestamp 1669390400
transform 1 0 25648 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_221
timestamp 1669390400
transform 1 0 26096 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_225
timestamp 1669390400
transform 1 0 26544 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_233
timestamp 1669390400
transform 1 0 27440 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_237
timestamp 1669390400
transform 1 0 27888 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_239
timestamp 1669390400
transform 1 0 28112 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_242
timestamp 1669390400
transform 1 0 28448 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_244
timestamp 1669390400
transform 1 0 28672 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_247
timestamp 1669390400
transform 1 0 29008 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_250
timestamp 1669390400
transform 1 0 29344 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_267
timestamp 1669390400
transform 1 0 31248 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_271
timestamp 1669390400
transform 1 0 31696 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_280
timestamp 1669390400
transform 1 0 32704 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_299
timestamp 1669390400
transform 1 0 34832 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_303
timestamp 1669390400
transform 1 0 35280 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_307
timestamp 1669390400
transform 1 0 35728 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_311
timestamp 1669390400
transform 1 0 36176 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_314
timestamp 1669390400
transform 1 0 36512 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_318
timestamp 1669390400
transform 1 0 36960 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_321
timestamp 1669390400
transform 1 0 37296 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_331
timestamp 1669390400
transform 1 0 38416 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_335
timestamp 1669390400
transform 1 0 38864 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_343
timestamp 1669390400
transform 1 0 39760 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_345
timestamp 1669390400
transform 1 0 39984 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_356
timestamp 1669390400
transform 1 0 41216 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_362
timestamp 1669390400
transform 1 0 41888 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_366
timestamp 1669390400
transform 1 0 42336 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_373
timestamp 1669390400
transform 1 0 43120 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_383
timestamp 1669390400
transform 1 0 44240 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_387
timestamp 1669390400
transform 1 0 44688 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_389
timestamp 1669390400
transform 1 0 44912 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_392
timestamp 1669390400
transform 1 0 45248 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_398
timestamp 1669390400
transform 1 0 45920 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_413
timestamp 1669390400
transform 1 0 47600 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_445
timestamp 1669390400
transform 1 0 51184 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_463
timestamp 1669390400
transform 1 0 53200 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_495
timestamp 1669390400
transform 1 0 56784 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_503
timestamp 1669390400
transform 1 0 57680 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_507
timestamp 1669390400
transform 1 0 58128 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_2
timestamp 1669390400
transform 1 0 1568 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_6
timestamp 1669390400
transform 1 0 2016 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_10
timestamp 1669390400
transform 1 0 2464 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_18
timestamp 1669390400
transform 1 0 3360 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_20
timestamp 1669390400
transform 1 0 3584 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_29
timestamp 1669390400
transform 1 0 4592 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_31
timestamp 1669390400
transform 1 0 4816 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_34
timestamp 1669390400
transform 1 0 5152 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_38
timestamp 1669390400
transform 1 0 5600 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_42
timestamp 1669390400
transform 1 0 6048 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_67
timestamp 1669390400
transform 1 0 8848 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_73
timestamp 1669390400
transform 1 0 9520 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_75
timestamp 1669390400
transform 1 0 9744 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_78
timestamp 1669390400
transform 1 0 10080 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_88
timestamp 1669390400
transform 1 0 11200 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_96
timestamp 1669390400
transform 1 0 12096 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_100
timestamp 1669390400
transform 1 0 12544 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_108
timestamp 1669390400
transform 1 0 13440 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_114
timestamp 1669390400
transform 1 0 14112 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_118
timestamp 1669390400
transform 1 0 14560 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_122
timestamp 1669390400
transform 1 0 15008 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_124
timestamp 1669390400
transform 1 0 15232 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_132
timestamp 1669390400
transform 1 0 16128 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_141
timestamp 1669390400
transform 1 0 17136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_144
timestamp 1669390400
transform 1 0 17472 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_147
timestamp 1669390400
transform 1 0 17808 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_153
timestamp 1669390400
transform 1 0 18480 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_155
timestamp 1669390400
transform 1 0 18704 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_158
timestamp 1669390400
transform 1 0 19040 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_170
timestamp 1669390400
transform 1 0 20384 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_176
timestamp 1669390400
transform 1 0 21056 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_184
timestamp 1669390400
transform 1 0 21952 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_192
timestamp 1669390400
transform 1 0 22848 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_199
timestamp 1669390400
transform 1 0 23632 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_208
timestamp 1669390400
transform 1 0 24640 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1669390400
transform 1 0 25088 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_215
timestamp 1669390400
transform 1 0 25424 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_218
timestamp 1669390400
transform 1 0 25760 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_222
timestamp 1669390400
transform 1 0 26208 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_224
timestamp 1669390400
transform 1 0 26432 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_233
timestamp 1669390400
transform 1 0 27440 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_244
timestamp 1669390400
transform 1 0 28672 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_248
timestamp 1669390400
transform 1 0 29120 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_252
timestamp 1669390400
transform 1 0 29568 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_256
timestamp 1669390400
transform 1 0 30016 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_260
timestamp 1669390400
transform 1 0 30464 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_264
timestamp 1669390400
transform 1 0 30912 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_266
timestamp 1669390400
transform 1 0 31136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_269
timestamp 1669390400
transform 1 0 31472 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_277
timestamp 1669390400
transform 1 0 32368 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_281
timestamp 1669390400
transform 1 0 32816 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_283
timestamp 1669390400
transform 1 0 33040 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_286
timestamp 1669390400
transform 1 0 33376 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_289
timestamp 1669390400
transform 1 0 33712 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_293
timestamp 1669390400
transform 1 0 34160 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_297
timestamp 1669390400
transform 1 0 34608 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_300
timestamp 1669390400
transform 1 0 34944 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_304
timestamp 1669390400
transform 1 0 35392 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_308
timestamp 1669390400
transform 1 0 35840 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_312
timestamp 1669390400
transform 1 0 36288 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_319
timestamp 1669390400
transform 1 0 37072 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_323
timestamp 1669390400
transform 1 0 37520 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_327
timestamp 1669390400
transform 1 0 37968 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_331
timestamp 1669390400
transform 1 0 38416 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_335
timestamp 1669390400
transform 1 0 38864 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_339
timestamp 1669390400
transform 1 0 39312 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_343
timestamp 1669390400
transform 1 0 39760 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_353
timestamp 1669390400
transform 1 0 40880 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_357
timestamp 1669390400
transform 1 0 41328 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_359
timestamp 1669390400
transform 1 0 41552 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_365
timestamp 1669390400
transform 1 0 42224 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_369
timestamp 1669390400
transform 1 0 42672 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_373
timestamp 1669390400
transform 1 0 43120 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_379
timestamp 1669390400
transform 1 0 43792 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_395
timestamp 1669390400
transform 1 0 45584 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_411
timestamp 1669390400
transform 1 0 47376 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_419
timestamp 1669390400
transform 1 0 48272 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_423
timestamp 1669390400
transform 1 0 48720 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_425
timestamp 1669390400
transform 1 0 48944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_428
timestamp 1669390400
transform 1 0 49280 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_492
timestamp 1669390400
transform 1 0 56448 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_496
timestamp 1669390400
transform 1 0 56896 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_499
timestamp 1669390400
transform 1 0 57232 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_507
timestamp 1669390400
transform 1 0 58128 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_2
timestamp 1669390400
transform 1 0 1568 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_17
timestamp 1669390400
transform 1 0 3248 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_21
timestamp 1669390400
transform 1 0 3696 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_24
timestamp 1669390400
transform 1 0 4032 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1669390400
transform 1 0 5152 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_37
timestamp 1669390400
transform 1 0 5488 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_43
timestamp 1669390400
transform 1 0 6160 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_53
timestamp 1669390400
transform 1 0 7280 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_59
timestamp 1669390400
transform 1 0 7952 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_63
timestamp 1669390400
transform 1 0 8400 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_67
timestamp 1669390400
transform 1 0 8848 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_71
timestamp 1669390400
transform 1 0 9296 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_79
timestamp 1669390400
transform 1 0 10192 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_81
timestamp 1669390400
transform 1 0 10416 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_105
timestamp 1669390400
transform 1 0 13104 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_108
timestamp 1669390400
transform 1 0 13440 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_118
timestamp 1669390400
transform 1 0 14560 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_122
timestamp 1669390400
transform 1 0 15008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_125
timestamp 1669390400
transform 1 0 15344 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_139
timestamp 1669390400
transform 1 0 16912 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_141
timestamp 1669390400
transform 1 0 17136 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_144
timestamp 1669390400
transform 1 0 17472 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_148
timestamp 1669390400
transform 1 0 17920 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_152
timestamp 1669390400
transform 1 0 18368 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_156
timestamp 1669390400
transform 1 0 18816 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_164
timestamp 1669390400
transform 1 0 19712 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_171
timestamp 1669390400
transform 1 0 20496 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_175
timestamp 1669390400
transform 1 0 20944 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_179
timestamp 1669390400
transform 1 0 21392 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_185
timestamp 1669390400
transform 1 0 22064 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_189
timestamp 1669390400
transform 1 0 22512 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_197
timestamp 1669390400
transform 1 0 23408 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_204
timestamp 1669390400
transform 1 0 24192 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_208
timestamp 1669390400
transform 1 0 24640 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_212
timestamp 1669390400
transform 1 0 25088 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_216
timestamp 1669390400
transform 1 0 25536 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_219
timestamp 1669390400
transform 1 0 25872 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_227
timestamp 1669390400
transform 1 0 26768 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_240
timestamp 1669390400
transform 1 0 28224 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_244
timestamp 1669390400
transform 1 0 28672 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_250
timestamp 1669390400
transform 1 0 29344 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_264
timestamp 1669390400
transform 1 0 30912 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_268
timestamp 1669390400
transform 1 0 31360 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_272
timestamp 1669390400
transform 1 0 31808 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_281
timestamp 1669390400
transform 1 0 32816 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_285
timestamp 1669390400
transform 1 0 33264 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_288
timestamp 1669390400
transform 1 0 33600 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_298
timestamp 1669390400
transform 1 0 34720 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1669390400
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_321
timestamp 1669390400
transform 1 0 37296 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_324
timestamp 1669390400
transform 1 0 37632 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_349
timestamp 1669390400
transform 1 0 40432 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_351
timestamp 1669390400
transform 1 0 40656 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_354
timestamp 1669390400
transform 1 0 40992 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_369
timestamp 1669390400
transform 1 0 42672 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_377
timestamp 1669390400
transform 1 0 43568 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_383
timestamp 1669390400
transform 1 0 44240 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_387
timestamp 1669390400
transform 1 0 44688 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1669390400
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_392
timestamp 1669390400
transform 1 0 45248 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_406
timestamp 1669390400
transform 1 0 46816 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_438
timestamp 1669390400
transform 1 0 50400 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_454
timestamp 1669390400
transform 1 0 52192 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_458
timestamp 1669390400
transform 1 0 52640 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_460
timestamp 1669390400
transform 1 0 52864 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_463
timestamp 1669390400
transform 1 0 53200 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_495
timestamp 1669390400
transform 1 0 56784 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_503
timestamp 1669390400
transform 1 0 57680 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_507
timestamp 1669390400
transform 1 0 58128 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_2
timestamp 1669390400
transform 1 0 1568 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_5
timestamp 1669390400
transform 1 0 1904 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_9
timestamp 1669390400
transform 1 0 2352 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_13
timestamp 1669390400
transform 1 0 2800 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_17
timestamp 1669390400
transform 1 0 3248 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_21
timestamp 1669390400
transform 1 0 3696 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_25
timestamp 1669390400
transform 1 0 4144 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_33
timestamp 1669390400
transform 1 0 5040 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_41
timestamp 1669390400
transform 1 0 5936 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_51
timestamp 1669390400
transform 1 0 7056 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_55
timestamp 1669390400
transform 1 0 7504 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_66
timestamp 1669390400
transform 1 0 8736 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_70
timestamp 1669390400
transform 1 0 9184 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_73
timestamp 1669390400
transform 1 0 9520 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_83
timestamp 1669390400
transform 1 0 10640 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_93
timestamp 1669390400
transform 1 0 11760 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_100
timestamp 1669390400
transform 1 0 12544 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_104
timestamp 1669390400
transform 1 0 12992 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_118
timestamp 1669390400
transform 1 0 14560 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_126
timestamp 1669390400
transform 1 0 15456 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_130
timestamp 1669390400
transform 1 0 15904 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1669390400
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_144
timestamp 1669390400
transform 1 0 17472 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_152
timestamp 1669390400
transform 1 0 18368 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_156
timestamp 1669390400
transform 1 0 18816 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_165
timestamp 1669390400
transform 1 0 19824 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_173
timestamp 1669390400
transform 1 0 20720 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_177
timestamp 1669390400
transform 1 0 21168 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_180
timestamp 1669390400
transform 1 0 21504 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_194
timestamp 1669390400
transform 1 0 23072 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_205
timestamp 1669390400
transform 1 0 24304 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_212
timestamp 1669390400
transform 1 0 25088 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_215
timestamp 1669390400
transform 1 0 25424 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_218
timestamp 1669390400
transform 1 0 25760 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_220
timestamp 1669390400
transform 1 0 25984 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_227
timestamp 1669390400
transform 1 0 26768 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_231
timestamp 1669390400
transform 1 0 27216 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_248
timestamp 1669390400
transform 1 0 29120 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_252
timestamp 1669390400
transform 1 0 29568 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_254
timestamp 1669390400
transform 1 0 29792 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_261
timestamp 1669390400
transform 1 0 30576 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_263
timestamp 1669390400
transform 1 0 30800 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_266
timestamp 1669390400
transform 1 0 31136 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1669390400
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_286
timestamp 1669390400
transform 1 0 33376 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_301
timestamp 1669390400
transform 1 0 35056 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_311
timestamp 1669390400
transform 1 0 36176 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_319
timestamp 1669390400
transform 1 0 37072 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_323
timestamp 1669390400
transform 1 0 37520 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_331
timestamp 1669390400
transform 1 0 38416 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_346
timestamp 1669390400
transform 1 0 40096 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_350
timestamp 1669390400
transform 1 0 40544 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_354
timestamp 1669390400
transform 1 0 40992 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_357
timestamp 1669390400
transform 1 0 41328 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_359
timestamp 1669390400
transform 1 0 41552 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_362
timestamp 1669390400
transform 1 0 41888 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_379
timestamp 1669390400
transform 1 0 43792 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_402
timestamp 1669390400
transform 1 0 46368 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_410
timestamp 1669390400
transform 1 0 47264 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_414
timestamp 1669390400
transform 1 0 47712 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_417
timestamp 1669390400
transform 1 0 48048 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_425
timestamp 1669390400
transform 1 0 48944 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_428
timestamp 1669390400
transform 1 0 49280 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_492
timestamp 1669390400
transform 1 0 56448 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_496
timestamp 1669390400
transform 1 0 56896 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_499
timestamp 1669390400
transform 1 0 57232 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_507
timestamp 1669390400
transform 1 0 58128 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_2
timestamp 1669390400
transform 1 0 1568 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_6
timestamp 1669390400
transform 1 0 2016 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_10
timestamp 1669390400
transform 1 0 2464 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_14
timestamp 1669390400
transform 1 0 2912 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_18
timestamp 1669390400
transform 1 0 3360 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_22
timestamp 1669390400
transform 1 0 3808 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_26
timestamp 1669390400
transform 1 0 4256 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_30
timestamp 1669390400
transform 1 0 4704 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_34
timestamp 1669390400
transform 1 0 5152 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_37
timestamp 1669390400
transform 1 0 5488 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_39
timestamp 1669390400
transform 1 0 5712 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_42
timestamp 1669390400
transform 1 0 6048 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_56
timestamp 1669390400
transform 1 0 7616 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_81
timestamp 1669390400
transform 1 0 10416 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_85
timestamp 1669390400
transform 1 0 10864 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_91
timestamp 1669390400
transform 1 0 11536 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1669390400
transform 1 0 13104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_108
timestamp 1669390400
transform 1 0 13440 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_119
timestamp 1669390400
transform 1 0 14672 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_127
timestamp 1669390400
transform 1 0 15568 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_131
timestamp 1669390400
transform 1 0 16016 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_140
timestamp 1669390400
transform 1 0 17024 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_146
timestamp 1669390400
transform 1 0 17696 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_156
timestamp 1669390400
transform 1 0 18816 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_168
timestamp 1669390400
transform 1 0 20160 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_175
timestamp 1669390400
transform 1 0 20944 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_179
timestamp 1669390400
transform 1 0 21392 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_181
timestamp 1669390400
transform 1 0 21616 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_184
timestamp 1669390400
transform 1 0 21952 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_193
timestamp 1669390400
transform 1 0 22960 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_205
timestamp 1669390400
transform 1 0 24304 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_214
timestamp 1669390400
transform 1 0 25312 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_218
timestamp 1669390400
transform 1 0 25760 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_238
timestamp 1669390400
transform 1 0 28000 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_240
timestamp 1669390400
transform 1 0 28224 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_247
timestamp 1669390400
transform 1 0 29008 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_250
timestamp 1669390400
transform 1 0 29344 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_264
timestamp 1669390400
transform 1 0 30912 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_266
timestamp 1669390400
transform 1 0 31136 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_269
timestamp 1669390400
transform 1 0 31472 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_279
timestamp 1669390400
transform 1 0 32592 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_286
timestamp 1669390400
transform 1 0 33376 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_293
timestamp 1669390400
transform 1 0 34160 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_297
timestamp 1669390400
transform 1 0 34608 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_314
timestamp 1669390400
transform 1 0 36512 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1669390400
transform 1 0 36960 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_321
timestamp 1669390400
transform 1 0 37296 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_326
timestamp 1669390400
transform 1 0 37856 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_335
timestamp 1669390400
transform 1 0 38864 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_339
timestamp 1669390400
transform 1 0 39312 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_343
timestamp 1669390400
transform 1 0 39760 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_347
timestamp 1669390400
transform 1 0 40208 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_351
timestamp 1669390400
transform 1 0 40656 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_355
timestamp 1669390400
transform 1 0 41104 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_361
timestamp 1669390400
transform 1 0 41776 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_376
timestamp 1669390400
transform 1 0 43456 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_380
timestamp 1669390400
transform 1 0 43904 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_382
timestamp 1669390400
transform 1 0 44128 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_389
timestamp 1669390400
transform 1 0 44912 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_392
timestamp 1669390400
transform 1 0 45248 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_401
timestamp 1669390400
transform 1 0 46256 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_433
timestamp 1669390400
transform 1 0 49840 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_449
timestamp 1669390400
transform 1 0 51632 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_457
timestamp 1669390400
transform 1 0 52528 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_463
timestamp 1669390400
transform 1 0 53200 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_471
timestamp 1669390400
transform 1 0 54096 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_475
timestamp 1669390400
transform 1 0 54544 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_491
timestamp 1669390400
transform 1 0 56336 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_507
timestamp 1669390400
transform 1 0 58128 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_2
timestamp 1669390400
transform 1 0 1568 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_8
timestamp 1669390400
transform 1 0 2240 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_12
timestamp 1669390400
transform 1 0 2688 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_16
timestamp 1669390400
transform 1 0 3136 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_20
timestamp 1669390400
transform 1 0 3584 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_24
timestamp 1669390400
transform 1 0 4032 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_28
timestamp 1669390400
transform 1 0 4480 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_32
timestamp 1669390400
transform 1 0 4928 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_36
timestamp 1669390400
transform 1 0 5376 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_40
timestamp 1669390400
transform 1 0 5824 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_44
timestamp 1669390400
transform 1 0 6272 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_48
timestamp 1669390400
transform 1 0 6720 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_50
timestamp 1669390400
transform 1 0 6944 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_56
timestamp 1669390400
transform 1 0 7616 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_62
timestamp 1669390400
transform 1 0 8288 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_66
timestamp 1669390400
transform 1 0 8736 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_70
timestamp 1669390400
transform 1 0 9184 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_73
timestamp 1669390400
transform 1 0 9520 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_77
timestamp 1669390400
transform 1 0 9968 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_81
timestamp 1669390400
transform 1 0 10416 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_88
timestamp 1669390400
transform 1 0 11200 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_113
timestamp 1669390400
transform 1 0 14000 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_117
timestamp 1669390400
transform 1 0 14448 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_121
timestamp 1669390400
transform 1 0 14896 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_125
timestamp 1669390400
transform 1 0 15344 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_129
timestamp 1669390400
transform 1 0 15792 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_133
timestamp 1669390400
transform 1 0 16240 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_137
timestamp 1669390400
transform 1 0 16688 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1669390400
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_144
timestamp 1669390400
transform 1 0 17472 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_147
timestamp 1669390400
transform 1 0 17808 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_151
timestamp 1669390400
transform 1 0 18256 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_154
timestamp 1669390400
transform 1 0 18592 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_158
timestamp 1669390400
transform 1 0 19040 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_162
timestamp 1669390400
transform 1 0 19488 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_166
timestamp 1669390400
transform 1 0 19936 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_169
timestamp 1669390400
transform 1 0 20272 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_173
timestamp 1669390400
transform 1 0 20720 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_181
timestamp 1669390400
transform 1 0 21616 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_191
timestamp 1669390400
transform 1 0 22736 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_193
timestamp 1669390400
transform 1 0 22960 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_196
timestamp 1669390400
transform 1 0 23296 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_200
timestamp 1669390400
transform 1 0 23744 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_204
timestamp 1669390400
transform 1 0 24192 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_207
timestamp 1669390400
transform 1 0 24528 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_211
timestamp 1669390400
transform 1 0 24976 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_215
timestamp 1669390400
transform 1 0 25424 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_217
timestamp 1669390400
transform 1 0 25648 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_223
timestamp 1669390400
transform 1 0 26320 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_233
timestamp 1669390400
transform 1 0 27440 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_240
timestamp 1669390400
transform 1 0 28224 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_244
timestamp 1669390400
transform 1 0 28672 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_248
timestamp 1669390400
transform 1 0 29120 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_252
timestamp 1669390400
transform 1 0 29568 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_256
timestamp 1669390400
transform 1 0 30016 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_260
timestamp 1669390400
transform 1 0 30464 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_268
timestamp 1669390400
transform 1 0 31360 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_272
timestamp 1669390400
transform 1 0 31808 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_276
timestamp 1669390400
transform 1 0 32256 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_278
timestamp 1669390400
transform 1 0 32480 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_281
timestamp 1669390400
transform 1 0 32816 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1669390400
transform 1 0 33040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_286
timestamp 1669390400
transform 1 0 33376 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_293
timestamp 1669390400
transform 1 0 34160 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_297
timestamp 1669390400
transform 1 0 34608 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_303
timestamp 1669390400
transform 1 0 35280 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_310
timestamp 1669390400
transform 1 0 36064 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_317
timestamp 1669390400
transform 1 0 36848 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_327
timestamp 1669390400
transform 1 0 37968 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_331
timestamp 1669390400
transform 1 0 38416 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_335
timestamp 1669390400
transform 1 0 38864 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_339
timestamp 1669390400
transform 1 0 39312 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_343
timestamp 1669390400
transform 1 0 39760 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_347
timestamp 1669390400
transform 1 0 40208 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_351
timestamp 1669390400
transform 1 0 40656 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1669390400
transform 1 0 40992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_357
timestamp 1669390400
transform 1 0 41328 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_370
timestamp 1669390400
transform 1 0 42784 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_374
timestamp 1669390400
transform 1 0 43232 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_381
timestamp 1669390400
transform 1 0 44016 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_63_407
timestamp 1669390400
transform 1 0 46928 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_423
timestamp 1669390400
transform 1 0 48720 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_425
timestamp 1669390400
transform 1 0 48944 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_428
timestamp 1669390400
transform 1 0 49280 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_492
timestamp 1669390400
transform 1 0 56448 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_496
timestamp 1669390400
transform 1 0 56896 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_499
timestamp 1669390400
transform 1 0 57232 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_507
timestamp 1669390400
transform 1 0 58128 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_2
timestamp 1669390400
transform 1 0 1568 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_5
timestamp 1669390400
transform 1 0 1904 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_9
timestamp 1669390400
transform 1 0 2352 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_13
timestamp 1669390400
transform 1 0 2800 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_17
timestamp 1669390400
transform 1 0 3248 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_21
timestamp 1669390400
transform 1 0 3696 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_25
timestamp 1669390400
transform 1 0 4144 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_29
timestamp 1669390400
transform 1 0 4592 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_31
timestamp 1669390400
transform 1 0 4816 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1669390400
transform 1 0 5152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_37
timestamp 1669390400
transform 1 0 5488 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_41
timestamp 1669390400
transform 1 0 5936 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_45
timestamp 1669390400
transform 1 0 6384 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_53
timestamp 1669390400
transform 1 0 7280 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_60
timestamp 1669390400
transform 1 0 8064 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_66
timestamp 1669390400
transform 1 0 8736 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_74
timestamp 1669390400
transform 1 0 9632 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_81
timestamp 1669390400
transform 1 0 10416 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_91
timestamp 1669390400
transform 1 0 11536 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_95
timestamp 1669390400
transform 1 0 11984 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_101
timestamp 1669390400
transform 1 0 12656 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1669390400
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_108
timestamp 1669390400
transform 1 0 13440 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_116
timestamp 1669390400
transform 1 0 14336 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_123
timestamp 1669390400
transform 1 0 15120 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_129
timestamp 1669390400
transform 1 0 15792 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_133
timestamp 1669390400
transform 1 0 16240 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_140
timestamp 1669390400
transform 1 0 17024 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_144
timestamp 1669390400
transform 1 0 17472 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_153
timestamp 1669390400
transform 1 0 18480 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_160
timestamp 1669390400
transform 1 0 19264 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_164
timestamp 1669390400
transform 1 0 19712 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_173
timestamp 1669390400
transform 1 0 20720 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_179
timestamp 1669390400
transform 1 0 21392 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_187
timestamp 1669390400
transform 1 0 22288 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_205
timestamp 1669390400
transform 1 0 24304 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_209
timestamp 1669390400
transform 1 0 24752 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_213
timestamp 1669390400
transform 1 0 25200 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_217
timestamp 1669390400
transform 1 0 25648 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_219
timestamp 1669390400
transform 1 0 25872 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_222
timestamp 1669390400
transform 1 0 26208 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_226
timestamp 1669390400
transform 1 0 26656 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_234
timestamp 1669390400
transform 1 0 27552 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_236
timestamp 1669390400
transform 1 0 27776 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1669390400
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_250
timestamp 1669390400
transform 1 0 29344 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_261
timestamp 1669390400
transform 1 0 30576 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_265
timestamp 1669390400
transform 1 0 31024 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_282
timestamp 1669390400
transform 1 0 32928 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_295
timestamp 1669390400
transform 1 0 34384 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_299
timestamp 1669390400
transform 1 0 34832 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_303
timestamp 1669390400
transform 1 0 35280 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_313
timestamp 1669390400
transform 1 0 36400 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_315
timestamp 1669390400
transform 1 0 36624 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1669390400
transform 1 0 36960 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_321
timestamp 1669390400
transform 1 0 37296 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_334
timestamp 1669390400
transform 1 0 38752 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_346
timestamp 1669390400
transform 1 0 40096 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_350
timestamp 1669390400
transform 1 0 40544 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_360
timestamp 1669390400
transform 1 0 41664 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_364
timestamp 1669390400
transform 1 0 42112 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_366
timestamp 1669390400
transform 1 0 42336 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_375
timestamp 1669390400
transform 1 0 43344 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_379
timestamp 1669390400
transform 1 0 43792 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_383
timestamp 1669390400
transform 1 0 44240 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_387
timestamp 1669390400
transform 1 0 44688 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1669390400
transform 1 0 44912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_392
timestamp 1669390400
transform 1 0 45248 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_402
timestamp 1669390400
transform 1 0 46368 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_434
timestamp 1669390400
transform 1 0 49952 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_450
timestamp 1669390400
transform 1 0 51744 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_458
timestamp 1669390400
transform 1 0 52640 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_460
timestamp 1669390400
transform 1 0 52864 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_463
timestamp 1669390400
transform 1 0 53200 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_495
timestamp 1669390400
transform 1 0 56784 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_503
timestamp 1669390400
transform 1 0 57680 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_507
timestamp 1669390400
transform 1 0 58128 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_2
timestamp 1669390400
transform 1 0 1568 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_4
timestamp 1669390400
transform 1 0 1792 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_7
timestamp 1669390400
transform 1 0 2128 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_11
timestamp 1669390400
transform 1 0 2576 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_15
timestamp 1669390400
transform 1 0 3024 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_19
timestamp 1669390400
transform 1 0 3472 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_23
timestamp 1669390400
transform 1 0 3920 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_27
timestamp 1669390400
transform 1 0 4368 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_31
timestamp 1669390400
transform 1 0 4816 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_35
timestamp 1669390400
transform 1 0 5264 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_39
timestamp 1669390400
transform 1 0 5712 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_43
timestamp 1669390400
transform 1 0 6160 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_47
timestamp 1669390400
transform 1 0 6608 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_51
timestamp 1669390400
transform 1 0 7056 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_55
timestamp 1669390400
transform 1 0 7504 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_57
timestamp 1669390400
transform 1 0 7728 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_60
timestamp 1669390400
transform 1 0 8064 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_70
timestamp 1669390400
transform 1 0 9184 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_73
timestamp 1669390400
transform 1 0 9520 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_83
timestamp 1669390400
transform 1 0 10640 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_108
timestamp 1669390400
transform 1 0 13440 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_125
timestamp 1669390400
transform 1 0 15344 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_138
timestamp 1669390400
transform 1 0 16800 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_144
timestamp 1669390400
transform 1 0 17472 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_160
timestamp 1669390400
transform 1 0 19264 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_166
timestamp 1669390400
transform 1 0 19936 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_178
timestamp 1669390400
transform 1 0 21280 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_188
timestamp 1669390400
transform 1 0 22400 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_190
timestamp 1669390400
transform 1 0 22624 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_193
timestamp 1669390400
transform 1 0 22960 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_195
timestamp 1669390400
transform 1 0 23184 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_202
timestamp 1669390400
transform 1 0 23968 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_204
timestamp 1669390400
transform 1 0 24192 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_210
timestamp 1669390400
transform 1 0 24864 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1669390400
transform 1 0 25088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_215
timestamp 1669390400
transform 1 0 25424 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_217
timestamp 1669390400
transform 1 0 25648 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_220
timestamp 1669390400
transform 1 0 25984 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_232
timestamp 1669390400
transform 1 0 27328 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_252
timestamp 1669390400
transform 1 0 29568 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_256
timestamp 1669390400
transform 1 0 30016 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_258
timestamp 1669390400
transform 1 0 30240 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_268
timestamp 1669390400
transform 1 0 31360 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1669390400
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_286
timestamp 1669390400
transform 1 0 33376 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_289
timestamp 1669390400
transform 1 0 33712 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_314
timestamp 1669390400
transform 1 0 36512 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_321
timestamp 1669390400
transform 1 0 37296 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_327
timestamp 1669390400
transform 1 0 37968 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_341
timestamp 1669390400
transform 1 0 39536 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_353
timestamp 1669390400
transform 1 0 40880 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_357
timestamp 1669390400
transform 1 0 41328 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_359
timestamp 1669390400
transform 1 0 41552 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_373
timestamp 1669390400
transform 1 0 43120 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_380
timestamp 1669390400
transform 1 0 43904 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_384
timestamp 1669390400
transform 1 0 44352 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_392
timestamp 1669390400
transform 1 0 45248 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_65_402
timestamp 1669390400
transform 1 0 46368 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_418
timestamp 1669390400
transform 1 0 48160 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_428
timestamp 1669390400
transform 1 0 49280 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_492
timestamp 1669390400
transform 1 0 56448 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_496
timestamp 1669390400
transform 1 0 56896 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_499
timestamp 1669390400
transform 1 0 57232 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_507
timestamp 1669390400
transform 1 0 58128 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_2
timestamp 1669390400
transform 1 0 1568 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_17
timestamp 1669390400
transform 1 0 3248 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_19
timestamp 1669390400
transform 1 0 3472 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_22
timestamp 1669390400
transform 1 0 3808 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_26
timestamp 1669390400
transform 1 0 4256 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_30
timestamp 1669390400
transform 1 0 4704 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_34
timestamp 1669390400
transform 1 0 5152 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_37
timestamp 1669390400
transform 1 0 5488 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_41
timestamp 1669390400
transform 1 0 5936 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_45
timestamp 1669390400
transform 1 0 6384 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_49
timestamp 1669390400
transform 1 0 6832 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_57
timestamp 1669390400
transform 1 0 7728 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_61
timestamp 1669390400
transform 1 0 8176 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_65
timestamp 1669390400
transform 1 0 8624 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_69
timestamp 1669390400
transform 1 0 9072 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_77
timestamp 1669390400
transform 1 0 9968 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_81
timestamp 1669390400
transform 1 0 10416 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_88
timestamp 1669390400
transform 1 0 11200 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_90
timestamp 1669390400
transform 1 0 11424 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_93
timestamp 1669390400
transform 1 0 11760 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_97
timestamp 1669390400
transform 1 0 12208 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_101
timestamp 1669390400
transform 1 0 12656 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_105
timestamp 1669390400
transform 1 0 13104 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_108
timestamp 1669390400
transform 1 0 13440 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_111
timestamp 1669390400
transform 1 0 13776 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_113
timestamp 1669390400
transform 1 0 14000 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_116
timestamp 1669390400
transform 1 0 14336 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_128
timestamp 1669390400
transform 1 0 15680 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_138
timestamp 1669390400
transform 1 0 16800 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_145
timestamp 1669390400
transform 1 0 17584 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_155
timestamp 1669390400
transform 1 0 18704 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_163
timestamp 1669390400
transform 1 0 19600 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_167
timestamp 1669390400
transform 1 0 20048 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_171
timestamp 1669390400
transform 1 0 20496 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_173
timestamp 1669390400
transform 1 0 20720 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_176
timestamp 1669390400
transform 1 0 21056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_179
timestamp 1669390400
transform 1 0 21392 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_189
timestamp 1669390400
transform 1 0 22512 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_199
timestamp 1669390400
transform 1 0 23632 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_207
timestamp 1669390400
transform 1 0 24528 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_214
timestamp 1669390400
transform 1 0 25312 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_220
timestamp 1669390400
transform 1 0 25984 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_224
timestamp 1669390400
transform 1 0 26432 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_228
timestamp 1669390400
transform 1 0 26880 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_232
timestamp 1669390400
transform 1 0 27328 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_236
timestamp 1669390400
transform 1 0 27776 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_247
timestamp 1669390400
transform 1 0 29008 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_250
timestamp 1669390400
transform 1 0 29344 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_259
timestamp 1669390400
transform 1 0 30352 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_263
timestamp 1669390400
transform 1 0 30800 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_272
timestamp 1669390400
transform 1 0 31808 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_276
timestamp 1669390400
transform 1 0 32256 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_280
timestamp 1669390400
transform 1 0 32704 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_284
timestamp 1669390400
transform 1 0 33152 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_288
timestamp 1669390400
transform 1 0 33600 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_292
timestamp 1669390400
transform 1 0 34048 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_296
timestamp 1669390400
transform 1 0 34496 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_304
timestamp 1669390400
transform 1 0 35392 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_312
timestamp 1669390400
transform 1 0 36288 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_316
timestamp 1669390400
transform 1 0 36736 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1669390400
transform 1 0 36960 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_321
timestamp 1669390400
transform 1 0 37296 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_324
timestamp 1669390400
transform 1 0 37632 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_328
timestamp 1669390400
transform 1 0 38080 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_330
timestamp 1669390400
transform 1 0 38304 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_337
timestamp 1669390400
transform 1 0 39088 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_347
timestamp 1669390400
transform 1 0 40208 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_351
timestamp 1669390400
transform 1 0 40656 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_353
timestamp 1669390400
transform 1 0 40880 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_359
timestamp 1669390400
transform 1 0 41552 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_363
timestamp 1669390400
transform 1 0 42000 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_365
timestamp 1669390400
transform 1 0 42224 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_378
timestamp 1669390400
transform 1 0 43680 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_380
timestamp 1669390400
transform 1 0 43904 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_389
timestamp 1669390400
transform 1 0 44912 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_392
timestamp 1669390400
transform 1 0 45248 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_406
timestamp 1669390400
transform 1 0 46816 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_414
timestamp 1669390400
transform 1 0 47712 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_446
timestamp 1669390400
transform 1 0 51296 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_454
timestamp 1669390400
transform 1 0 52192 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_458
timestamp 1669390400
transform 1 0 52640 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_460
timestamp 1669390400
transform 1 0 52864 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_463
timestamp 1669390400
transform 1 0 53200 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_467
timestamp 1669390400
transform 1 0 53648 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_471
timestamp 1669390400
transform 1 0 54096 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_475
timestamp 1669390400
transform 1 0 54544 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_491
timestamp 1669390400
transform 1 0 56336 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_507
timestamp 1669390400
transform 1 0 58128 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_2
timestamp 1669390400
transform 1 0 1568 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_19
timestamp 1669390400
transform 1 0 3472 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_23
timestamp 1669390400
transform 1 0 3920 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_26
timestamp 1669390400
transform 1 0 4256 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_30
timestamp 1669390400
transform 1 0 4704 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_34
timestamp 1669390400
transform 1 0 5152 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_37
timestamp 1669390400
transform 1 0 5488 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_43
timestamp 1669390400
transform 1 0 6160 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_47
timestamp 1669390400
transform 1 0 6608 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_63
timestamp 1669390400
transform 1 0 8400 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_69
timestamp 1669390400
transform 1 0 9072 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_72
timestamp 1669390400
transform 1 0 9408 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_76
timestamp 1669390400
transform 1 0 9856 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_80
timestamp 1669390400
transform 1 0 10304 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_84
timestamp 1669390400
transform 1 0 10752 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_88
timestamp 1669390400
transform 1 0 11200 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_104
timestamp 1669390400
transform 1 0 12992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_107
timestamp 1669390400
transform 1 0 13328 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_111
timestamp 1669390400
transform 1 0 13776 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_115
timestamp 1669390400
transform 1 0 14224 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_119
timestamp 1669390400
transform 1 0 14672 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_123
timestamp 1669390400
transform 1 0 15120 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_127
timestamp 1669390400
transform 1 0 15568 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_131
timestamp 1669390400
transform 1 0 16016 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_135
timestamp 1669390400
transform 1 0 16464 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_139
timestamp 1669390400
transform 1 0 16912 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_142
timestamp 1669390400
transform 1 0 17248 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_145
timestamp 1669390400
transform 1 0 17584 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_149
timestamp 1669390400
transform 1 0 18032 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_165
timestamp 1669390400
transform 1 0 19824 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_169
timestamp 1669390400
transform 1 0 20272 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_171
timestamp 1669390400
transform 1 0 20496 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_174
timestamp 1669390400
transform 1 0 20832 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_177
timestamp 1669390400
transform 1 0 21168 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_180
timestamp 1669390400
transform 1 0 21504 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_186
timestamp 1669390400
transform 1 0 22176 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_193
timestamp 1669390400
transform 1 0 22960 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_209
timestamp 1669390400
transform 1 0 24752 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_212
timestamp 1669390400
transform 1 0 25088 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_215
timestamp 1669390400
transform 1 0 25424 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_219
timestamp 1669390400
transform 1 0 25872 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_223
timestamp 1669390400
transform 1 0 26320 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_227
timestamp 1669390400
transform 1 0 26768 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_231
timestamp 1669390400
transform 1 0 27216 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_234
timestamp 1669390400
transform 1 0 27552 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_244
timestamp 1669390400
transform 1 0 28672 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_247
timestamp 1669390400
transform 1 0 29008 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_264
timestamp 1669390400
transform 1 0 30912 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_268
timestamp 1669390400
transform 1 0 31360 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_272
timestamp 1669390400
transform 1 0 31808 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_276
timestamp 1669390400
transform 1 0 32256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_282
timestamp 1669390400
transform 1 0 32928 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_285
timestamp 1669390400
transform 1 0 33264 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_289
timestamp 1669390400
transform 1 0 33712 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_293
timestamp 1669390400
transform 1 0 34160 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_297
timestamp 1669390400
transform 1 0 34608 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_299
timestamp 1669390400
transform 1 0 34832 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_314
timestamp 1669390400
transform 1 0 36512 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_317
timestamp 1669390400
transform 1 0 36848 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_320
timestamp 1669390400
transform 1 0 37184 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_324
timestamp 1669390400
transform 1 0 37632 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_328
timestamp 1669390400
transform 1 0 38080 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_332
timestamp 1669390400
transform 1 0 38528 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_336
timestamp 1669390400
transform 1 0 38976 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_338
timestamp 1669390400
transform 1 0 39200 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_345
timestamp 1669390400
transform 1 0 39984 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_349
timestamp 1669390400
transform 1 0 40432 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_352
timestamp 1669390400
transform 1 0 40768 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_367
timestamp 1669390400
transform 1 0 42448 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_371
timestamp 1669390400
transform 1 0 42896 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_375
timestamp 1669390400
transform 1 0 43344 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_379
timestamp 1669390400
transform 1 0 43792 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_383
timestamp 1669390400
transform 1 0 44240 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_387
timestamp 1669390400
transform 1 0 44688 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_395
timestamp 1669390400
transform 1 0 45584 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_401
timestamp 1669390400
transform 1 0 46256 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_417
timestamp 1669390400
transform 1 0 48048 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_419
timestamp 1669390400
transform 1 0 48272 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_422
timestamp 1669390400
transform 1 0 48608 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_454
timestamp 1669390400
transform 1 0 52192 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_457
timestamp 1669390400
transform 1 0 52528 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_472
timestamp 1669390400
transform 1 0 54208 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_474
timestamp 1669390400
transform 1 0 54432 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_489
timestamp 1669390400
transform 1 0 56112 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_492
timestamp 1669390400
transform 1 0 56448 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_508
timestamp 1669390400
transform 1 0 58240 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1669390400
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1669390400
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1669390400
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1669390400
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1669390400
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1669390400
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1669390400
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1669390400
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1669390400
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1669390400
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1669390400
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1669390400
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1669390400
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1669390400
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1669390400
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1669390400
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1669390400
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1669390400
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1669390400
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1669390400
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1669390400
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1669390400
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1669390400
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1669390400
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1669390400
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1669390400
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1669390400
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1669390400
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1669390400
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1669390400
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1669390400
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1669390400
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1669390400
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1669390400
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1669390400
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1669390400
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1669390400
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1669390400
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1669390400
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1669390400
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1669390400
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1669390400
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1669390400
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1669390400
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1669390400
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1669390400
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1669390400
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1669390400
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1669390400
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1669390400
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1669390400
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1669390400
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1669390400
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1669390400
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1669390400
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1669390400
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1669390400
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1669390400
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1669390400
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1669390400
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1669390400
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1669390400
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1669390400
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1669390400
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1669390400
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1669390400
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1669390400
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1669390400
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1669390400
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1669390400
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1669390400
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1669390400
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1669390400
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1669390400
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1669390400
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1669390400
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1669390400
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1669390400
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1669390400
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1669390400
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1669390400
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1669390400
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1669390400
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1669390400
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1669390400
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1669390400
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1669390400
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1669390400
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1669390400
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1669390400
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1669390400
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1669390400
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1669390400
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1669390400
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1669390400
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1669390400
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1669390400
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1669390400
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1669390400
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1669390400
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1669390400
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1669390400
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1669390400
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1669390400
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1669390400
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1669390400
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1669390400
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1669390400
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1669390400
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1669390400
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1669390400
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1669390400
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1669390400
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1669390400
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1669390400
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1669390400
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1669390400
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1669390400
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1669390400
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1669390400
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1669390400
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1669390400
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1669390400
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1669390400
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1669390400
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1669390400
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1669390400
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1669390400
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1669390400
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1669390400
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1669390400
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1669390400
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1669390400
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1669390400
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1669390400
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1669390400
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1669390400
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1669390400
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1669390400
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1669390400
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1669390400
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1669390400
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1669390400
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1669390400
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1669390400
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1669390400
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1669390400
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1669390400
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1669390400
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1669390400
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1669390400
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1669390400
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1669390400
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1669390400
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1669390400
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1669390400
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1669390400
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1669390400
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1669390400
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1669390400
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1669390400
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1669390400
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1669390400
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1669390400
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1669390400
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1669390400
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1669390400
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1669390400
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1669390400
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1669390400
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1669390400
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1669390400
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1669390400
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1669390400
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1669390400
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1669390400
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1669390400
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1669390400
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1669390400
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1669390400
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1669390400
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1669390400
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1669390400
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1669390400
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1669390400
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1669390400
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1669390400
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1669390400
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1669390400
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1669390400
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1669390400
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1669390400
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1669390400
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1669390400
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1669390400
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1669390400
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1669390400
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1669390400
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1669390400
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1669390400
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1669390400
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1669390400
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1669390400
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1669390400
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1669390400
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1669390400
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1669390400
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1669390400
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1669390400
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1669390400
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1669390400
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1669390400
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1669390400
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1669390400
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1669390400
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1669390400
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1669390400
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1669390400
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1669390400
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1669390400
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1669390400
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1669390400
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1669390400
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1669390400
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1669390400
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1669390400
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1669390400
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1669390400
transform 1 0 5264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1669390400
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1669390400
transform 1 0 13104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1669390400
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1669390400
transform 1 0 20944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1669390400
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1669390400
transform 1 0 28784 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1669390400
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1669390400
transform 1 0 36624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1669390400
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1669390400
transform 1 0 44464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1669390400
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1669390400
transform 1 0 52304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1669390400
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1346_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 57904 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1347_
timestamp 1669390400
transform 1 0 56896 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1348_
timestamp 1669390400
transform 1 0 57344 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1349_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 57008 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1350_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 55552 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1351_
timestamp 1669390400
transform 1 0 56224 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1352_
timestamp 1669390400
transform -1 0 54992 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1353_
timestamp 1669390400
transform -1 0 53984 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1354_
timestamp 1669390400
transform -1 0 52192 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1355_
timestamp 1669390400
transform -1 0 52752 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1356_
timestamp 1669390400
transform -1 0 56896 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1357_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 51856 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1358_
timestamp 1669390400
transform -1 0 31472 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1359_
timestamp 1669390400
transform -1 0 51632 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1360_
timestamp 1669390400
transform -1 0 54432 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1361_
timestamp 1669390400
transform -1 0 51968 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1362_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 50736 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1363_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 30464 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1364_
timestamp 1669390400
transform 1 0 50512 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1365_
timestamp 1669390400
transform 1 0 55216 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1366_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 58016 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1367_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 55664 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1368_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 51408 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1369_
timestamp 1669390400
transform 1 0 57344 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1370_
timestamp 1669390400
transform -1 0 58240 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1371_
timestamp 1669390400
transform -1 0 57904 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1372_
timestamp 1669390400
transform 1 0 55216 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1373_
timestamp 1669390400
transform -1 0 57792 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1374_
timestamp 1669390400
transform 1 0 57456 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1375_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 56896 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1376_
timestamp 1669390400
transform -1 0 33040 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1377_
timestamp 1669390400
transform -1 0 28672 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1378_
timestamp 1669390400
transform -1 0 50848 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1379_
timestamp 1669390400
transform -1 0 44912 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1380_
timestamp 1669390400
transform -1 0 55440 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1381_
timestamp 1669390400
transform 1 0 53312 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1382_
timestamp 1669390400
transform -1 0 52864 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1383_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 57344 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1384_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 52640 0 -1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1385_
timestamp 1669390400
transform -1 0 35728 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1386_
timestamp 1669390400
transform -1 0 27776 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1387_
timestamp 1669390400
transform -1 0 27664 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1388_
timestamp 1669390400
transform 1 0 21504 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1389_
timestamp 1669390400
transform -1 0 9296 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1390_
timestamp 1669390400
transform -1 0 8960 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1391_
timestamp 1669390400
transform -1 0 8176 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1392_
timestamp 1669390400
transform -1 0 10752 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1393_
timestamp 1669390400
transform -1 0 5264 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1394_
timestamp 1669390400
transform 1 0 4480 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1395_
timestamp 1669390400
transform -1 0 6944 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1396_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 9632 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1397_
timestamp 1669390400
transform -1 0 22176 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1398_
timestamp 1669390400
transform 1 0 5600 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1399_
timestamp 1669390400
transform -1 0 7168 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1400_
timestamp 1669390400
transform 1 0 9408 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1401_
timestamp 1669390400
transform 1 0 13552 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1402_
timestamp 1669390400
transform 1 0 20608 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1403_
timestamp 1669390400
transform -1 0 2352 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1404_
timestamp 1669390400
transform -1 0 7840 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1405_
timestamp 1669390400
transform -1 0 7056 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1406_
timestamp 1669390400
transform 1 0 21392 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1407_
timestamp 1669390400
transform 1 0 23296 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1408_
timestamp 1669390400
transform 1 0 24528 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1409_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 22400 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1410_
timestamp 1669390400
transform 1 0 10976 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1411_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 10752 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1412_
timestamp 1669390400
transform 1 0 13440 0 -1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1413_
timestamp 1669390400
transform 1 0 26208 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1414_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 25984 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1415_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 23520 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1416_
timestamp 1669390400
transform 1 0 31472 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1417_
timestamp 1669390400
transform -1 0 32928 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1418_
timestamp 1669390400
transform -1 0 25984 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1419_
timestamp 1669390400
transform -1 0 25872 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1420_
timestamp 1669390400
transform -1 0 24528 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1421_
timestamp 1669390400
transform 1 0 23072 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1422_
timestamp 1669390400
transform -1 0 26432 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1423_
timestamp 1669390400
transform 1 0 24976 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1424_
timestamp 1669390400
transform 1 0 38192 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1425_
timestamp 1669390400
transform -1 0 30688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1426_
timestamp 1669390400
transform -1 0 28560 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1427_
timestamp 1669390400
transform -1 0 27440 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1428_
timestamp 1669390400
transform -1 0 26096 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1429_
timestamp 1669390400
transform -1 0 25200 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1430_
timestamp 1669390400
transform -1 0 27216 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1431_
timestamp 1669390400
transform 1 0 25536 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1432_
timestamp 1669390400
transform -1 0 25088 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1433_
timestamp 1669390400
transform 1 0 22848 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1434_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 30688 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1435_
timestamp 1669390400
transform -1 0 32928 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1436_
timestamp 1669390400
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1437_
timestamp 1669390400
transform -1 0 30128 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1438_
timestamp 1669390400
transform -1 0 32032 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1439_
timestamp 1669390400
transform 1 0 29568 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1440_
timestamp 1669390400
transform 1 0 29568 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1441_
timestamp 1669390400
transform -1 0 31248 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1442_
timestamp 1669390400
transform 1 0 17584 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1443_
timestamp 1669390400
transform 1 0 18704 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1444_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 20160 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1445_
timestamp 1669390400
transform -1 0 18592 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1446_
timestamp 1669390400
transform -1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1447_
timestamp 1669390400
transform 1 0 25984 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1448_
timestamp 1669390400
transform -1 0 27664 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1449_
timestamp 1669390400
transform -1 0 30576 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1450_
timestamp 1669390400
transform 1 0 29232 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1451_
timestamp 1669390400
transform 1 0 36400 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1452_
timestamp 1669390400
transform -1 0 21168 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1453_
timestamp 1669390400
transform -1 0 19824 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1454_
timestamp 1669390400
transform -1 0 10528 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1455_
timestamp 1669390400
transform 1 0 10416 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1456_
timestamp 1669390400
transform -1 0 12208 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1457_
timestamp 1669390400
transform -1 0 6272 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1458_
timestamp 1669390400
transform -1 0 24752 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1459_
timestamp 1669390400
transform 1 0 19488 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1460_
timestamp 1669390400
transform -1 0 2576 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1461_
timestamp 1669390400
transform 1 0 1680 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1462_
timestamp 1669390400
transform 1 0 8176 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1463_
timestamp 1669390400
transform -1 0 20832 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1464_
timestamp 1669390400
transform -1 0 4480 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1465_
timestamp 1669390400
transform -1 0 4032 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1466_
timestamp 1669390400
transform 1 0 3472 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1467_
timestamp 1669390400
transform -1 0 2464 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1468_
timestamp 1669390400
transform 1 0 1680 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1469_
timestamp 1669390400
transform 1 0 3696 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1470_
timestamp 1669390400
transform -1 0 6944 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1471_
timestamp 1669390400
transform -1 0 5824 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1472_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4592 0 -1 42336
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1473_
timestamp 1669390400
transform 1 0 14672 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1474_
timestamp 1669390400
transform -1 0 16688 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1475_
timestamp 1669390400
transform 1 0 7168 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1476_
timestamp 1669390400
transform 1 0 17696 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1477_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 18368 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1478_
timestamp 1669390400
transform -1 0 16016 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1479_
timestamp 1669390400
transform -1 0 15120 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1480_
timestamp 1669390400
transform 1 0 14112 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1481_
timestamp 1669390400
transform 1 0 3472 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1482_
timestamp 1669390400
transform -1 0 3472 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1483_
timestamp 1669390400
transform 1 0 2576 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1484_
timestamp 1669390400
transform -1 0 3472 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1485_
timestamp 1669390400
transform 1 0 2464 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1486_
timestamp 1669390400
transform 1 0 3696 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1487_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2576 0 -1 40768
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1488_
timestamp 1669390400
transform 1 0 21504 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1489_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 19712 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1490_
timestamp 1669390400
transform 1 0 6048 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1491_
timestamp 1669390400
transform 1 0 15680 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1492_
timestamp 1669390400
transform -1 0 22960 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1493_
timestamp 1669390400
transform 1 0 21840 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1494_
timestamp 1669390400
transform 1 0 22960 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1495_
timestamp 1669390400
transform 1 0 24416 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1496_
timestamp 1669390400
transform 1 0 25088 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1497_
timestamp 1669390400
transform 1 0 28112 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1498_
timestamp 1669390400
transform -1 0 23856 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1499_
timestamp 1669390400
transform 1 0 17360 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1500_
timestamp 1669390400
transform 1 0 16576 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1501_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6944 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1502_
timestamp 1669390400
transform 1 0 6048 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1503_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7280 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1504_
timestamp 1669390400
transform 1 0 7728 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1505_
timestamp 1669390400
transform 1 0 10752 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1506_
timestamp 1669390400
transform 1 0 4480 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1507_
timestamp 1669390400
transform 1 0 10192 0 -1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1508_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 19824 0 1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1509_
timestamp 1669390400
transform 1 0 10080 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1510_
timestamp 1669390400
transform 1 0 2688 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1511_
timestamp 1669390400
transform -1 0 9520 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1512_
timestamp 1669390400
transform 1 0 8288 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1513_
timestamp 1669390400
transform 1 0 12432 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1514_
timestamp 1669390400
transform 1 0 12320 0 -1 36064
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1515_
timestamp 1669390400
transform 1 0 4816 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1516_
timestamp 1669390400
transform 1 0 20384 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1517_
timestamp 1669390400
transform 1 0 21504 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1518_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 6608 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1519_
timestamp 1669390400
transform -1 0 7728 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1520_
timestamp 1669390400
transform 1 0 4480 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1521_
timestamp 1669390400
transform 1 0 2688 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _1522_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6384 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1523_
timestamp 1669390400
transform -1 0 7168 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1524_
timestamp 1669390400
transform 1 0 7392 0 -1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1525_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 18032 0 -1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1526_
timestamp 1669390400
transform 1 0 37408 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1527_
timestamp 1669390400
transform -1 0 37856 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1528_
timestamp 1669390400
transform 1 0 37296 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1529_
timestamp 1669390400
transform 1 0 30464 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1530_
timestamp 1669390400
transform -1 0 31584 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1531_
timestamp 1669390400
transform 1 0 23632 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1532_
timestamp 1669390400
transform 1 0 16464 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1533_
timestamp 1669390400
transform 1 0 2800 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1534_
timestamp 1669390400
transform -1 0 4480 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1535_
timestamp 1669390400
transform 1 0 13776 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1536_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 10192 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1537_
timestamp 1669390400
transform 1 0 12208 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1538_
timestamp 1669390400
transform -1 0 12208 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1539_
timestamp 1669390400
transform 1 0 14672 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1540_
timestamp 1669390400
transform 1 0 4144 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1541_
timestamp 1669390400
transform 1 0 15008 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1542_
timestamp 1669390400
transform -1 0 17808 0 1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1543_
timestamp 1669390400
transform 1 0 7280 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1544_
timestamp 1669390400
transform 1 0 2240 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1545_
timestamp 1669390400
transform -1 0 9184 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1546_
timestamp 1669390400
transform -1 0 8176 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1547_
timestamp 1669390400
transform 1 0 5600 0 1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1548_
timestamp 1669390400
transform -1 0 21056 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1549_
timestamp 1669390400
transform -1 0 24304 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1550_
timestamp 1669390400
transform -1 0 18928 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1551_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 20384 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1552_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 23072 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1553_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 23072 0 -1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1554_
timestamp 1669390400
transform 1 0 25312 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1555_
timestamp 1669390400
transform 1 0 28896 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1556_
timestamp 1669390400
transform -1 0 29792 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1557_
timestamp 1669390400
transform -1 0 2912 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1558_
timestamp 1669390400
transform 1 0 28336 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1559_
timestamp 1669390400
transform -1 0 30912 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1560_
timestamp 1669390400
transform -1 0 37072 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1561_
timestamp 1669390400
transform 1 0 31360 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1562_
timestamp 1669390400
transform -1 0 33264 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1563_
timestamp 1669390400
transform 1 0 22400 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1564_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2800 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1565_
timestamp 1669390400
transform 1 0 9632 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1566_
timestamp 1669390400
transform 1 0 16464 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _1567_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17584 0 -1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1568_
timestamp 1669390400
transform 1 0 22064 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1569_
timestamp 1669390400
transform -1 0 24416 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1570_
timestamp 1669390400
transform 1 0 2576 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1571_
timestamp 1669390400
transform -1 0 2688 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1572_
timestamp 1669390400
transform -1 0 4032 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1573_
timestamp 1669390400
transform -1 0 2912 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1574_
timestamp 1669390400
transform -1 0 4816 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1575_
timestamp 1669390400
transform -1 0 4368 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1576_
timestamp 1669390400
transform -1 0 11872 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1577_
timestamp 1669390400
transform -1 0 15344 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1578_
timestamp 1669390400
transform 1 0 11088 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1579_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 14784 0 -1 37632
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1580_
timestamp 1669390400
transform -1 0 32480 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1581_
timestamp 1669390400
transform 1 0 31696 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1582_
timestamp 1669390400
transform 1 0 33488 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1583_
timestamp 1669390400
transform 1 0 2576 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1584_
timestamp 1669390400
transform 1 0 1680 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1585_
timestamp 1669390400
transform -1 0 2912 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1586_
timestamp 1669390400
transform 1 0 2688 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1587_
timestamp 1669390400
transform 1 0 3584 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1588_
timestamp 1669390400
transform 1 0 15008 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1589_
timestamp 1669390400
transform 1 0 2688 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1590_
timestamp 1669390400
transform -1 0 12544 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1591_
timestamp 1669390400
transform 1 0 9632 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1592_
timestamp 1669390400
transform -1 0 11200 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1593_
timestamp 1669390400
transform 1 0 13552 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1594_
timestamp 1669390400
transform -1 0 15456 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1595_
timestamp 1669390400
transform 1 0 13216 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1596_
timestamp 1669390400
transform -1 0 11312 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1597_
timestamp 1669390400
transform 1 0 18704 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1598_
timestamp 1669390400
transform 1 0 2912 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1599_
timestamp 1669390400
transform 1 0 12656 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1600_
timestamp 1669390400
transform -1 0 21840 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1601_
timestamp 1669390400
transform 1 0 22624 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1602_
timestamp 1669390400
transform 1 0 22064 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1603_
timestamp 1669390400
transform -1 0 24416 0 -1 43904
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1604_
timestamp 1669390400
transform -1 0 27664 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1605_
timestamp 1669390400
transform 1 0 26544 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1606_
timestamp 1669390400
transform -1 0 27888 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1607_
timestamp 1669390400
transform 1 0 28112 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1608_
timestamp 1669390400
transform -1 0 20160 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1609_
timestamp 1669390400
transform 1 0 22960 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1610_
timestamp 1669390400
transform 1 0 4592 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1611_
timestamp 1669390400
transform 1 0 4368 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1612_
timestamp 1669390400
transform 1 0 11424 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1613_
timestamp 1669390400
transform 1 0 18592 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1614_
timestamp 1669390400
transform 1 0 9296 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1615_
timestamp 1669390400
transform 1 0 19040 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1616_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 19264 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1617_
timestamp 1669390400
transform 1 0 6160 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1618_
timestamp 1669390400
transform 1 0 7280 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1619_
timestamp 1669390400
transform -1 0 11312 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1620_
timestamp 1669390400
transform 1 0 10416 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1621_
timestamp 1669390400
transform 1 0 14896 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1622_
timestamp 1669390400
transform -1 0 16352 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1623_
timestamp 1669390400
transform 1 0 18368 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1624_
timestamp 1669390400
transform 1 0 19376 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1625_
timestamp 1669390400
transform 1 0 21504 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1626_
timestamp 1669390400
transform 1 0 18256 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1627_
timestamp 1669390400
transform 1 0 17696 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1628_
timestamp 1669390400
transform 1 0 19712 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1629_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 21168 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1630_
timestamp 1669390400
transform 1 0 28336 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1631_
timestamp 1669390400
transform 1 0 35616 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1632_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 34272 0 1 36064
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1633_
timestamp 1669390400
transform -1 0 39424 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1634_
timestamp 1669390400
transform -1 0 34944 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1635_
timestamp 1669390400
transform -1 0 35504 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1636_
timestamp 1669390400
transform -1 0 36512 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1637_
timestamp 1669390400
transform -1 0 36064 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1638_
timestamp 1669390400
transform 1 0 30912 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1639_
timestamp 1669390400
transform 1 0 33488 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1640_
timestamp 1669390400
transform -1 0 24192 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1641_
timestamp 1669390400
transform -1 0 13888 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1642_
timestamp 1669390400
transform 1 0 8512 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1643_
timestamp 1669390400
transform -1 0 12880 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1644_
timestamp 1669390400
transform 1 0 13552 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1645_
timestamp 1669390400
transform -1 0 14112 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1646_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13552 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1647_
timestamp 1669390400
transform 1 0 2800 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1648_
timestamp 1669390400
transform 1 0 15792 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1649_
timestamp 1669390400
transform -1 0 21056 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1650_
timestamp 1669390400
transform 1 0 16800 0 1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1651_
timestamp 1669390400
transform -1 0 5152 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1652_
timestamp 1669390400
transform 1 0 6720 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1653_
timestamp 1669390400
transform 1 0 21504 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1654_
timestamp 1669390400
transform 1 0 22848 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1655_
timestamp 1669390400
transform -1 0 23856 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1656_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 33040 0 -1 39200
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1657_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 33824 0 -1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1658_
timestamp 1669390400
transform 1 0 36736 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1659_
timestamp 1669390400
transform 1 0 16016 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1660_
timestamp 1669390400
transform -1 0 6496 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1661_
timestamp 1669390400
transform -1 0 10864 0 1 37632
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1662_
timestamp 1669390400
transform -1 0 11872 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1663_
timestamp 1669390400
transform -1 0 17136 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1664_
timestamp 1669390400
transform 1 0 3472 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1665_
timestamp 1669390400
transform -1 0 10752 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1666_
timestamp 1669390400
transform 1 0 10976 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1667_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17584 0 -1 39200
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1668_
timestamp 1669390400
transform 1 0 26544 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1669_
timestamp 1669390400
transform -1 0 26880 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1670_
timestamp 1669390400
transform 1 0 27104 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1671_
timestamp 1669390400
transform 1 0 25536 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1672_
timestamp 1669390400
transform -1 0 28112 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1673_
timestamp 1669390400
transform -1 0 27216 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1674_
timestamp 1669390400
transform -1 0 18144 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1675_
timestamp 1669390400
transform -1 0 17920 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1676_
timestamp 1669390400
transform 1 0 9408 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1677_
timestamp 1669390400
transform -1 0 12320 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1678_
timestamp 1669390400
transform -1 0 7616 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1679_
timestamp 1669390400
transform 1 0 9744 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1680_
timestamp 1669390400
transform -1 0 7280 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _1681_
timestamp 1669390400
transform 1 0 10304 0 1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1682_
timestamp 1669390400
transform 1 0 6384 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1683_
timestamp 1669390400
transform 1 0 15680 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1684_
timestamp 1669390400
transform -1 0 16912 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1685_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 16128 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1686_
timestamp 1669390400
transform -1 0 19600 0 -1 42336
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1687_
timestamp 1669390400
transform 1 0 29456 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1688_
timestamp 1669390400
transform 1 0 29232 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1689_
timestamp 1669390400
transform 1 0 37744 0 1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1690_
timestamp 1669390400
transform 1 0 38416 0 1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1691_
timestamp 1669390400
transform -1 0 39984 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1692_
timestamp 1669390400
transform 1 0 41440 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1693_
timestamp 1669390400
transform 1 0 41216 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1694_
timestamp 1669390400
transform 1 0 41440 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1695_
timestamp 1669390400
transform 1 0 37968 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1696_
timestamp 1669390400
transform -1 0 39760 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1697_
timestamp 1669390400
transform 1 0 38192 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1698_
timestamp 1669390400
transform -1 0 39648 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1699_
timestamp 1669390400
transform 1 0 1904 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1700_
timestamp 1669390400
transform -1 0 4480 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1701_
timestamp 1669390400
transform 1 0 6608 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1702_
timestamp 1669390400
transform 1 0 11648 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1703_
timestamp 1669390400
transform 1 0 11760 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1704_
timestamp 1669390400
transform 1 0 12992 0 -1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1705_
timestamp 1669390400
transform 1 0 2688 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1706_
timestamp 1669390400
transform -1 0 18256 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1707_
timestamp 1669390400
transform -1 0 14448 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1708_
timestamp 1669390400
transform 1 0 12544 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1709_
timestamp 1669390400
transform 1 0 6608 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1710_
timestamp 1669390400
transform -1 0 14560 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1711_
timestamp 1669390400
transform -1 0 5824 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1712_
timestamp 1669390400
transform 1 0 4256 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1713_
timestamp 1669390400
transform 1 0 3696 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1714_
timestamp 1669390400
transform 1 0 3808 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1715_
timestamp 1669390400
transform 1 0 2688 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1716_
timestamp 1669390400
transform 1 0 3136 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1717_
timestamp 1669390400
transform -1 0 12880 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1718_
timestamp 1669390400
transform 1 0 3472 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1719_
timestamp 1669390400
transform 1 0 3696 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1720_
timestamp 1669390400
transform 1 0 4704 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1721_
timestamp 1669390400
transform 1 0 13552 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1722_
timestamp 1669390400
transform 1 0 12768 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1723_
timestamp 1669390400
transform 1 0 13664 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1724_
timestamp 1669390400
transform -1 0 7056 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1725_
timestamp 1669390400
transform 1 0 18816 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1726_
timestamp 1669390400
transform 1 0 25648 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1727_
timestamp 1669390400
transform 1 0 27104 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1728_
timestamp 1669390400
transform 1 0 27888 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1729_
timestamp 1669390400
transform -1 0 29008 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1730_
timestamp 1669390400
transform 1 0 37520 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1731_
timestamp 1669390400
transform 1 0 4032 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1732_
timestamp 1669390400
transform 1 0 7840 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1733_
timestamp 1669390400
transform 1 0 6272 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1734_
timestamp 1669390400
transform -1 0 13104 0 1 34496
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _1735_
timestamp 1669390400
transform 1 0 7952 0 1 43904
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1736_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 22736 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1737_
timestamp 1669390400
transform 1 0 30464 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1738_
timestamp 1669390400
transform -1 0 17696 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1739_
timestamp 1669390400
transform -1 0 11872 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1740_
timestamp 1669390400
transform 1 0 16352 0 -1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1741_
timestamp 1669390400
transform 1 0 21616 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1742_
timestamp 1669390400
transform -1 0 10416 0 -1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1743_
timestamp 1669390400
transform -1 0 9520 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1744_
timestamp 1669390400
transform 1 0 8624 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _1745_
timestamp 1669390400
transform -1 0 10416 0 1 45472
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1746_
timestamp 1669390400
transform -1 0 11088 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1747_
timestamp 1669390400
transform 1 0 30352 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1748_
timestamp 1669390400
transform 1 0 31472 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1749_
timestamp 1669390400
transform 1 0 31920 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1750_
timestamp 1669390400
transform 1 0 32032 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1751_
timestamp 1669390400
transform -1 0 36176 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1752_
timestamp 1669390400
transform 1 0 32480 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1753_
timestamp 1669390400
transform -1 0 34496 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1754_
timestamp 1669390400
transform 1 0 37296 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1755_
timestamp 1669390400
transform 1 0 34496 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1756_
timestamp 1669390400
transform 1 0 35952 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1757_
timestamp 1669390400
transform -1 0 35392 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1758_
timestamp 1669390400
transform -1 0 35168 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1759_
timestamp 1669390400
transform 1 0 34160 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1760_
timestamp 1669390400
transform 1 0 35504 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1761_
timestamp 1669390400
transform -1 0 28336 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1762_
timestamp 1669390400
transform 1 0 28224 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1763_
timestamp 1669390400
transform -1 0 7504 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _1764_
timestamp 1669390400
transform -1 0 8848 0 -1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1765_
timestamp 1669390400
transform 1 0 7840 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1766_
timestamp 1669390400
transform 1 0 8064 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1767_
timestamp 1669390400
transform -1 0 4032 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1768_
timestamp 1669390400
transform 1 0 8736 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1769_
timestamp 1669390400
transform -1 0 9184 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1770_
timestamp 1669390400
transform -1 0 11536 0 1 40768
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1771_
timestamp 1669390400
transform 1 0 26656 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1772_
timestamp 1669390400
transform 1 0 38528 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1773_
timestamp 1669390400
transform 1 0 37632 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1774_
timestamp 1669390400
transform 1 0 38864 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1775_
timestamp 1669390400
transform 1 0 40320 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1776_
timestamp 1669390400
transform 1 0 40208 0 1 39200
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1777_
timestamp 1669390400
transform -1 0 43568 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1778_
timestamp 1669390400
transform -1 0 2912 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1779_
timestamp 1669390400
transform 1 0 25648 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1780_
timestamp 1669390400
transform 1 0 26768 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1781_
timestamp 1669390400
transform -1 0 26432 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1782_
timestamp 1669390400
transform -1 0 23632 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1783_
timestamp 1669390400
transform 1 0 9856 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1784_
timestamp 1669390400
transform -1 0 13440 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1785_
timestamp 1669390400
transform 1 0 13776 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1786_
timestamp 1669390400
transform 1 0 14448 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1787_
timestamp 1669390400
transform 1 0 14896 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1788_
timestamp 1669390400
transform 1 0 16464 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1789_
timestamp 1669390400
transform -1 0 22176 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1790_
timestamp 1669390400
transform 1 0 16016 0 1 48608
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1791_
timestamp 1669390400
transform -1 0 7168 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1792_
timestamp 1669390400
transform 1 0 16576 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1793_
timestamp 1669390400
transform 1 0 16240 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1794_
timestamp 1669390400
transform -1 0 18368 0 1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1795_
timestamp 1669390400
transform 1 0 27776 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1796_
timestamp 1669390400
transform 1 0 26656 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1797_
timestamp 1669390400
transform 1 0 31248 0 1 42336
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1798_
timestamp 1669390400
transform 1 0 32704 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1799_
timestamp 1669390400
transform -1 0 20720 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1800_
timestamp 1669390400
transform -1 0 15456 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1801_
timestamp 1669390400
transform 1 0 12768 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1802_
timestamp 1669390400
transform 1 0 13552 0 1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1803_
timestamp 1669390400
transform 1 0 13664 0 -1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1804_
timestamp 1669390400
transform -1 0 11200 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1805_
timestamp 1669390400
transform -1 0 11536 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1806_
timestamp 1669390400
transform 1 0 10528 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1807_
timestamp 1669390400
transform -1 0 9184 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1808_
timestamp 1669390400
transform 1 0 9296 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1809_
timestamp 1669390400
transform -1 0 7056 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1810_
timestamp 1669390400
transform 1 0 5264 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1811_
timestamp 1669390400
transform -1 0 10640 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1812_
timestamp 1669390400
transform 1 0 10864 0 -1 54880
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1813_
timestamp 1669390400
transform 1 0 11424 0 -1 53312
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1814_
timestamp 1669390400
transform 1 0 34160 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1815_
timestamp 1669390400
transform 1 0 34048 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1816_
timestamp 1669390400
transform 1 0 35392 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1817_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 26320 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1818_
timestamp 1669390400
transform 1 0 29456 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1819_
timestamp 1669390400
transform -1 0 17136 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1820_
timestamp 1669390400
transform -1 0 11760 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1821_
timestamp 1669390400
transform -1 0 11536 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1822_
timestamp 1669390400
transform 1 0 10304 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1823_
timestamp 1669390400
transform -1 0 6160 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1824_
timestamp 1669390400
transform 1 0 7056 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1825_
timestamp 1669390400
transform 1 0 9520 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1826_
timestamp 1669390400
transform -1 0 10640 0 -1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1827_
timestamp 1669390400
transform 1 0 10528 0 1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1828_
timestamp 1669390400
transform 1 0 29344 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1829_
timestamp 1669390400
transform 1 0 37744 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1830_
timestamp 1669390400
transform 1 0 37520 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1831_
timestamp 1669390400
transform -1 0 39648 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1832_
timestamp 1669390400
transform 1 0 42224 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1833_
timestamp 1669390400
transform 1 0 42560 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1834_
timestamp 1669390400
transform 1 0 43568 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1835_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 39536 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1836_
timestamp 1669390400
transform -1 0 40992 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1837_
timestamp 1669390400
transform -1 0 44576 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1838_
timestamp 1669390400
transform 1 0 43568 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1839_
timestamp 1669390400
transform 1 0 42784 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1840_
timestamp 1669390400
transform -1 0 42896 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1841_
timestamp 1669390400
transform 1 0 41440 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1842_
timestamp 1669390400
transform 1 0 42336 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1843_
timestamp 1669390400
transform 1 0 43456 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1844_
timestamp 1669390400
transform -1 0 44912 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1845_
timestamp 1669390400
transform -1 0 2912 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1846_
timestamp 1669390400
transform 1 0 42784 0 1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1847_
timestamp 1669390400
transform 1 0 35392 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1848_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6384 0 1 48608
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1849_
timestamp 1669390400
transform 1 0 18032 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1850_
timestamp 1669390400
transform -1 0 20944 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1851_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 27328 0 1 45472
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1852_
timestamp 1669390400
transform -1 0 12208 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1853_
timestamp 1669390400
transform 1 0 22288 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1854_
timestamp 1669390400
transform 1 0 24080 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1855_
timestamp 1669390400
transform -1 0 32032 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1856_
timestamp 1669390400
transform -1 0 33264 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1857_
timestamp 1669390400
transform 1 0 33376 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1858_
timestamp 1669390400
transform 1 0 36624 0 -1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1859_
timestamp 1669390400
transform 1 0 6496 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1860_
timestamp 1669390400
transform -1 0 19264 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1861_
timestamp 1669390400
transform -1 0 11424 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1862_
timestamp 1669390400
transform 1 0 19712 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1863_
timestamp 1669390400
transform 1 0 10752 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1864_
timestamp 1669390400
transform -1 0 20720 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1865_
timestamp 1669390400
transform 1 0 29568 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1866_
timestamp 1669390400
transform 1 0 29792 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1867_
timestamp 1669390400
transform 1 0 21280 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1868_
timestamp 1669390400
transform -1 0 22848 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1869_
timestamp 1669390400
transform 1 0 19936 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1870_
timestamp 1669390400
transform 1 0 23072 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1871_
timestamp 1669390400
transform 1 0 23968 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1872_
timestamp 1669390400
transform 1 0 22736 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1873_
timestamp 1669390400
transform 1 0 17584 0 -1 48608
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1874_
timestamp 1669390400
transform 1 0 13664 0 -1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1875_
timestamp 1669390400
transform 1 0 22960 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1876_
timestamp 1669390400
transform 1 0 24416 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1877_
timestamp 1669390400
transform 1 0 13328 0 -1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1878_
timestamp 1669390400
transform -1 0 28784 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1879_
timestamp 1669390400
transform 1 0 26544 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1880_
timestamp 1669390400
transform -1 0 27552 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1881_
timestamp 1669390400
transform 1 0 28112 0 1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _1882_
timestamp 1669390400
transform 1 0 39312 0 1 43904
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1883_
timestamp 1669390400
transform -1 0 44688 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1884_
timestamp 1669390400
transform 1 0 43792 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1885_
timestamp 1669390400
transform 1 0 44688 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1886_
timestamp 1669390400
transform 1 0 43568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1887_
timestamp 1669390400
transform 1 0 45360 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1888_
timestamp 1669390400
transform 1 0 46368 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1889_
timestamp 1669390400
transform 1 0 47376 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1890_
timestamp 1669390400
transform -1 0 33040 0 -1 45472
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1891_
timestamp 1669390400
transform 1 0 4256 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1892_
timestamp 1669390400
transform 1 0 15344 0 -1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1893_
timestamp 1669390400
transform -1 0 16912 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1894_
timestamp 1669390400
transform 1 0 13552 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1895_
timestamp 1669390400
transform -1 0 15456 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1896_
timestamp 1669390400
transform -1 0 18368 0 -1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1897_
timestamp 1669390400
transform 1 0 16016 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1898_
timestamp 1669390400
transform 1 0 33600 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1899_
timestamp 1669390400
transform 1 0 33488 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1900_
timestamp 1669390400
transform 1 0 34832 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1901_
timestamp 1669390400
transform -1 0 30464 0 -1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1902_
timestamp 1669390400
transform 1 0 29904 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1903_
timestamp 1669390400
transform 1 0 12432 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1904_
timestamp 1669390400
transform 1 0 13552 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1905_
timestamp 1669390400
transform 1 0 22400 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1906_
timestamp 1669390400
transform -1 0 31248 0 1 48608
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1907_
timestamp 1669390400
transform -1 0 38752 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1908_
timestamp 1669390400
transform -1 0 38192 0 -1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1909_
timestamp 1669390400
transform 1 0 13664 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1910_
timestamp 1669390400
transform 1 0 16128 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1911_
timestamp 1669390400
transform 1 0 17920 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1912_
timestamp 1669390400
transform 1 0 11984 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1913_
timestamp 1669390400
transform 1 0 13552 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1914_
timestamp 1669390400
transform 1 0 13216 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1915_
timestamp 1669390400
transform 1 0 21728 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1916_
timestamp 1669390400
transform 1 0 22848 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1917_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 25872 0 1 47040
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1918_
timestamp 1669390400
transform 1 0 26544 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1919_
timestamp 1669390400
transform 1 0 29456 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1920_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 37408 0 -1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1921_
timestamp 1669390400
transform 1 0 37408 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1922_
timestamp 1669390400
transform 1 0 39648 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1923_
timestamp 1669390400
transform 1 0 38528 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1924_
timestamp 1669390400
transform 1 0 39424 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1925_
timestamp 1669390400
transform 1 0 39424 0 -1 45472
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1926_
timestamp 1669390400
transform -1 0 40768 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1927_
timestamp 1669390400
transform 1 0 40768 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1928_
timestamp 1669390400
transform 1 0 44240 0 -1 40768
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1929_
timestamp 1669390400
transform 1 0 45808 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1930_
timestamp 1669390400
transform -1 0 46032 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1931_
timestamp 1669390400
transform -1 0 44576 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1932_
timestamp 1669390400
transform -1 0 44912 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1933_
timestamp 1669390400
transform -1 0 7728 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1934_
timestamp 1669390400
transform 1 0 36288 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1935_
timestamp 1669390400
transform -1 0 37072 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1936_
timestamp 1669390400
transform 1 0 36288 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1937_
timestamp 1669390400
transform 1 0 32144 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1938_
timestamp 1669390400
transform -1 0 10416 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1939_
timestamp 1669390400
transform 1 0 8288 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1940_
timestamp 1669390400
transform -1 0 7280 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1941_
timestamp 1669390400
transform 1 0 7504 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1942_
timestamp 1669390400
transform 1 0 6272 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1943_
timestamp 1669390400
transform 1 0 7616 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1944_
timestamp 1669390400
transform -1 0 10416 0 1 51744
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1945_
timestamp 1669390400
transform -1 0 33040 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1946_
timestamp 1669390400
transform -1 0 34832 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1947_
timestamp 1669390400
transform 1 0 33712 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1948_
timestamp 1669390400
transform -1 0 36960 0 1 50176
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1949_
timestamp 1669390400
transform 1 0 10976 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1950_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 11760 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1951_
timestamp 1669390400
transform 1 0 20384 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1952_
timestamp 1669390400
transform -1 0 25088 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1953_
timestamp 1669390400
transform 1 0 23184 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1954_
timestamp 1669390400
transform 1 0 29568 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1955_
timestamp 1669390400
transform 1 0 37408 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1956_
timestamp 1669390400
transform -1 0 29008 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1957_
timestamp 1669390400
transform -1 0 24528 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1958_
timestamp 1669390400
transform 1 0 18928 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1959_
timestamp 1669390400
transform 1 0 17024 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai33_1  _1960_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 17584 0 -1 54880
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1961_
timestamp 1669390400
transform 1 0 24304 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1962_
timestamp 1669390400
transform -1 0 28224 0 1 50176
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1963_
timestamp 1669390400
transform 1 0 27664 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1964_
timestamp 1669390400
transform 1 0 37856 0 1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1965_
timestamp 1669390400
transform 1 0 39984 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1966_
timestamp 1669390400
transform 1 0 40096 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1967_
timestamp 1669390400
transform 1 0 42560 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1968_
timestamp 1669390400
transform -1 0 41888 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1969_
timestamp 1669390400
transform 1 0 41440 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1970_
timestamp 1669390400
transform 1 0 45024 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1971_
timestamp 1669390400
transform -1 0 43904 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1972_
timestamp 1669390400
transform -1 0 44576 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1973_
timestamp 1669390400
transform -1 0 2912 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1974_
timestamp 1669390400
transform -1 0 20944 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1975_
timestamp 1669390400
transform 1 0 19488 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1976_
timestamp 1669390400
transform 1 0 19824 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1977_
timestamp 1669390400
transform 1 0 14560 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1978_
timestamp 1669390400
transform 1 0 8960 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1979_
timestamp 1669390400
transform 1 0 14560 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1980_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 15568 0 -1 54880
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1981_
timestamp 1669390400
transform -1 0 21280 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1982_
timestamp 1669390400
transform 1 0 32816 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1983_
timestamp 1669390400
transform 1 0 31696 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1984_
timestamp 1669390400
transform 1 0 34048 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1985_
timestamp 1669390400
transform 1 0 36400 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1986_
timestamp 1669390400
transform 1 0 18928 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1987_
timestamp 1669390400
transform 1 0 19040 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1988_
timestamp 1669390400
transform 1 0 26096 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1989_
timestamp 1669390400
transform -1 0 26768 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1990_
timestamp 1669390400
transform 1 0 27664 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1991_
timestamp 1669390400
transform 1 0 41216 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1992_
timestamp 1669390400
transform -1 0 27552 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1993_
timestamp 1669390400
transform 1 0 19600 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1994_
timestamp 1669390400
transform 1 0 21504 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1995_
timestamp 1669390400
transform 1 0 21504 0 1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1996_
timestamp 1669390400
transform 1 0 26208 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1997_
timestamp 1669390400
transform 1 0 27552 0 -1 54880
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1998_
timestamp 1669390400
transform 1 0 42000 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1999_
timestamp 1669390400
transform 1 0 38304 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2000_
timestamp 1669390400
transform 1 0 37744 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2001_
timestamp 1669390400
transform -1 0 40096 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2002_
timestamp 1669390400
transform 1 0 45360 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2003_
timestamp 1669390400
transform 1 0 44128 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2004_
timestamp 1669390400
transform 1 0 45360 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2005_
timestamp 1669390400
transform 1 0 43344 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2006_
timestamp 1669390400
transform 1 0 43344 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2007_
timestamp 1669390400
transform 1 0 45360 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2008_
timestamp 1669390400
transform 1 0 46144 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2009_
timestamp 1669390400
transform 1 0 48048 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2010_
timestamp 1669390400
transform 1 0 41664 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2011_
timestamp 1669390400
transform 1 0 42112 0 -1 51744
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2012_
timestamp 1669390400
transform 1 0 20944 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2013_
timestamp 1669390400
transform -1 0 18816 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2014_
timestamp 1669390400
transform 1 0 18032 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2015_
timestamp 1669390400
transform 1 0 18704 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2016_
timestamp 1669390400
transform 1 0 21840 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2017_
timestamp 1669390400
transform 1 0 22512 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2018_
timestamp 1669390400
transform -1 0 33040 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2019_
timestamp 1669390400
transform 1 0 32928 0 1 48608
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2020_
timestamp 1669390400
transform 1 0 33488 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2021_
timestamp 1669390400
transform 1 0 22176 0 1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2022_
timestamp 1669390400
transform 1 0 24528 0 1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2023_
timestamp 1669390400
transform 1 0 27664 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2024_
timestamp 1669390400
transform 1 0 26544 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2025_
timestamp 1669390400
transform -1 0 33040 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2026_
timestamp 1669390400
transform 1 0 30688 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2027_
timestamp 1669390400
transform 1 0 21840 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2028_
timestamp 1669390400
transform 1 0 22400 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2029_
timestamp 1669390400
transform 1 0 24752 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2030_
timestamp 1669390400
transform 1 0 16464 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2031_
timestamp 1669390400
transform 1 0 17584 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2032_
timestamp 1669390400
transform 1 0 22960 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2033_
timestamp 1669390400
transform -1 0 30352 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2034_
timestamp 1669390400
transform 1 0 27888 0 1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2035_
timestamp 1669390400
transform 1 0 31024 0 1 54880
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2036_
timestamp 1669390400
transform 1 0 31472 0 1 53312
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2037_
timestamp 1669390400
transform 1 0 44240 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2038_
timestamp 1669390400
transform 1 0 44688 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2039_
timestamp 1669390400
transform 1 0 45696 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2040_
timestamp 1669390400
transform 1 0 44240 0 -1 53312
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2041_
timestamp 1669390400
transform -1 0 46368 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2042_
timestamp 1669390400
transform 1 0 33600 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2043_
timestamp 1669390400
transform 1 0 35280 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2044_
timestamp 1669390400
transform 1 0 16128 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2045_
timestamp 1669390400
transform 1 0 23296 0 -1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2046_
timestamp 1669390400
transform 1 0 35056 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2047_
timestamp 1669390400
transform 1 0 36288 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2048_
timestamp 1669390400
transform -1 0 26320 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2049_
timestamp 1669390400
transform -1 0 28000 0 1 51744
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2050_
timestamp 1669390400
transform -1 0 38752 0 1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2051_
timestamp 1669390400
transform 1 0 37520 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2052_
timestamp 1669390400
transform 1 0 23296 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2053_
timestamp 1669390400
transform -1 0 28672 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2054_
timestamp 1669390400
transform 1 0 27888 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2055_
timestamp 1669390400
transform 1 0 29792 0 1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2056_
timestamp 1669390400
transform 1 0 34720 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2057_
timestamp 1669390400
transform 1 0 38192 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2058_
timestamp 1669390400
transform 1 0 30352 0 -1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2059_
timestamp 1669390400
transform -1 0 34384 0 1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2060_
timestamp 1669390400
transform 1 0 41664 0 -1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2061_
timestamp 1669390400
transform 1 0 43456 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2062_
timestamp 1669390400
transform -1 0 46256 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2063_
timestamp 1669390400
transform -1 0 46368 0 -1 51744
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2064_
timestamp 1669390400
transform -1 0 43680 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2065_
timestamp 1669390400
transform -1 0 36288 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2066_
timestamp 1669390400
transform 1 0 37296 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2067_
timestamp 1669390400
transform 1 0 38416 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2068_
timestamp 1669390400
transform 1 0 23632 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2069_
timestamp 1669390400
transform 1 0 24080 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2070_
timestamp 1669390400
transform 1 0 31696 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2071_
timestamp 1669390400
transform -1 0 32816 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2072_
timestamp 1669390400
transform -1 0 35056 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2073_
timestamp 1669390400
transform 1 0 33936 0 -1 54880
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2074_
timestamp 1669390400
transform -1 0 40208 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2075_
timestamp 1669390400
transform 1 0 39760 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2076_
timestamp 1669390400
transform 1 0 40992 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2077_
timestamp 1669390400
transform -1 0 43904 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2078_
timestamp 1669390400
transform -1 0 44912 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2079_
timestamp 1669390400
transform 1 0 45360 0 1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2080_
timestamp 1669390400
transform 1 0 47040 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2081_
timestamp 1669390400
transform -1 0 43344 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2082_
timestamp 1669390400
transform 1 0 39200 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2083_
timestamp 1669390400
transform 1 0 40768 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2084_
timestamp 1669390400
transform 1 0 36736 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2085_
timestamp 1669390400
transform 1 0 35504 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2086_
timestamp 1669390400
transform 1 0 35504 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2087_
timestamp 1669390400
transform 1 0 41440 0 -1 53312
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2088_
timestamp 1669390400
transform 1 0 42000 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2089_
timestamp 1669390400
transform 1 0 48272 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2090_
timestamp 1669390400
transform 1 0 47040 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2091_
timestamp 1669390400
transform 1 0 48048 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2092_
timestamp 1669390400
transform -1 0 47376 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2093_
timestamp 1669390400
transform -1 0 53536 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2094_
timestamp 1669390400
transform -1 0 51856 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2095_
timestamp 1669390400
transform -1 0 56672 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2096_
timestamp 1669390400
transform -1 0 49952 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2097_
timestamp 1669390400
transform -1 0 50960 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2098_
timestamp 1669390400
transform -1 0 49840 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2099_
timestamp 1669390400
transform -1 0 52864 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2100_
timestamp 1669390400
transform -1 0 51744 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2101_
timestamp 1669390400
transform 1 0 43792 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2102_
timestamp 1669390400
transform 1 0 47712 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2103_
timestamp 1669390400
transform -1 0 44688 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2104_
timestamp 1669390400
transform -1 0 55776 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2105_
timestamp 1669390400
transform -1 0 55104 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2106_
timestamp 1669390400
transform 1 0 43344 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2107_
timestamp 1669390400
transform -1 0 58128 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2108_
timestamp 1669390400
transform -1 0 56896 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2109_
timestamp 1669390400
transform -1 0 55776 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2110_
timestamp 1669390400
transform -1 0 58016 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2111_
timestamp 1669390400
transform 1 0 43680 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2112_
timestamp 1669390400
transform -1 0 54656 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2113_
timestamp 1669390400
transform 1 0 52864 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2114_
timestamp 1669390400
transform 1 0 43792 0 -1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2115_
timestamp 1669390400
transform -1 0 57232 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2116_
timestamp 1669390400
transform -1 0 55216 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2117_
timestamp 1669390400
transform -1 0 54544 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2118_
timestamp 1669390400
transform -1 0 53984 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2119_
timestamp 1669390400
transform 1 0 50624 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2120_
timestamp 1669390400
transform -1 0 54544 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2121_
timestamp 1669390400
transform 1 0 54656 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2122_
timestamp 1669390400
transform -1 0 51184 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2123_
timestamp 1669390400
transform 1 0 50400 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2124_
timestamp 1669390400
transform 1 0 54880 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2125_
timestamp 1669390400
transform -1 0 53648 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2126_
timestamp 1669390400
transform 1 0 51632 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2127_
timestamp 1669390400
transform 1 0 56560 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2128_
timestamp 1669390400
transform 1 0 54880 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2129_
timestamp 1669390400
transform -1 0 50288 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2130_
timestamp 1669390400
transform 1 0 40208 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2131_
timestamp 1669390400
transform -1 0 56560 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2132_
timestamp 1669390400
transform -1 0 46032 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2133_
timestamp 1669390400
transform -1 0 57232 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2134_
timestamp 1669390400
transform -1 0 56000 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2135_
timestamp 1669390400
transform -1 0 51856 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2136_
timestamp 1669390400
transform -1 0 43344 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2137_
timestamp 1669390400
transform 1 0 43344 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2138_
timestamp 1669390400
transform -1 0 44688 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2139_
timestamp 1669390400
transform -1 0 46368 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2140_
timestamp 1669390400
transform 1 0 42448 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2141_
timestamp 1669390400
transform 1 0 43904 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2142_
timestamp 1669390400
transform 1 0 45360 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2143_
timestamp 1669390400
transform 1 0 52304 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2144_
timestamp 1669390400
transform 1 0 54656 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2145_
timestamp 1669390400
transform -1 0 52864 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2146_
timestamp 1669390400
transform 1 0 54208 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2147_
timestamp 1669390400
transform -1 0 55664 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _2148_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 58016 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2149_
timestamp 1669390400
transform -1 0 57568 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2150_
timestamp 1669390400
transform -1 0 55776 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2151_
timestamp 1669390400
transform 1 0 53312 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2152_
timestamp 1669390400
transform -1 0 53872 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2153_
timestamp 1669390400
transform -1 0 54992 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2154_
timestamp 1669390400
transform 1 0 53312 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2155_
timestamp 1669390400
transform 1 0 53312 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2156_
timestamp 1669390400
transform -1 0 52864 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2157_
timestamp 1669390400
transform -1 0 53648 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2158_
timestamp 1669390400
transform 1 0 57344 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2159_
timestamp 1669390400
transform 1 0 54432 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2160_
timestamp 1669390400
transform -1 0 52640 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2161_
timestamp 1669390400
transform -1 0 54208 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2162_
timestamp 1669390400
transform -1 0 54432 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2163_
timestamp 1669390400
transform 1 0 51520 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _2164_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 58128 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2165_
timestamp 1669390400
transform -1 0 57008 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2166_
timestamp 1669390400
transform 1 0 52192 0 -1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2167_
timestamp 1669390400
transform -1 0 53760 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2168_
timestamp 1669390400
transform -1 0 53088 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2169_
timestamp 1669390400
transform 1 0 44240 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2170_
timestamp 1669390400
transform -1 0 50064 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2171_
timestamp 1669390400
transform -1 0 50624 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2172_
timestamp 1669390400
transform -1 0 54432 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2173_
timestamp 1669390400
transform -1 0 54432 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2174_
timestamp 1669390400
transform 1 0 51184 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2175_
timestamp 1669390400
transform -1 0 48496 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2176_
timestamp 1669390400
transform 1 0 49392 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2177_
timestamp 1669390400
transform -1 0 50064 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2178_
timestamp 1669390400
transform -1 0 58016 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2179_
timestamp 1669390400
transform -1 0 49280 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2180_
timestamp 1669390400
transform -1 0 56896 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2181_
timestamp 1669390400
transform 1 0 48048 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2182_
timestamp 1669390400
transform -1 0 49728 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2183_
timestamp 1669390400
transform -1 0 47824 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2184_
timestamp 1669390400
transform 1 0 47600 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2185_
timestamp 1669390400
transform 1 0 52416 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2186_
timestamp 1669390400
transform 1 0 53984 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2187_
timestamp 1669390400
transform 1 0 55776 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2188_
timestamp 1669390400
transform 1 0 52304 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2189_
timestamp 1669390400
transform 1 0 54992 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2190_
timestamp 1669390400
transform 1 0 46704 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2191_
timestamp 1669390400
transform -1 0 47824 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2192_
timestamp 1669390400
transform 1 0 54544 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2193_
timestamp 1669390400
transform 1 0 46816 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2194_
timestamp 1669390400
transform -1 0 47488 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2195_
timestamp 1669390400
transform 1 0 47488 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2196_
timestamp 1669390400
transform 1 0 46368 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2197_
timestamp 1669390400
transform 1 0 46704 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2198_
timestamp 1669390400
transform 1 0 47040 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2199_
timestamp 1669390400
transform -1 0 47936 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2200_
timestamp 1669390400
transform -1 0 47824 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2201_
timestamp 1669390400
transform -1 0 45024 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2202_
timestamp 1669390400
transform 1 0 51408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2203_
timestamp 1669390400
transform -1 0 44576 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2204_
timestamp 1669390400
transform -1 0 47264 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2205_
timestamp 1669390400
transform -1 0 44912 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2206_
timestamp 1669390400
transform -1 0 45920 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2207_
timestamp 1669390400
transform -1 0 51184 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2208_
timestamp 1669390400
transform 1 0 43792 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2209_
timestamp 1669390400
transform 1 0 43792 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2210_
timestamp 1669390400
transform 1 0 44800 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2211_
timestamp 1669390400
transform -1 0 44912 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2212_
timestamp 1669390400
transform 1 0 44464 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2213_
timestamp 1669390400
transform -1 0 45696 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2214_
timestamp 1669390400
transform -1 0 44016 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2215_
timestamp 1669390400
transform 1 0 43344 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2216_
timestamp 1669390400
transform -1 0 56112 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2217_
timestamp 1669390400
transform 1 0 48048 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2218_
timestamp 1669390400
transform 1 0 48272 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2219_
timestamp 1669390400
transform -1 0 52080 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2220_
timestamp 1669390400
transform -1 0 48944 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2221_
timestamp 1669390400
transform -1 0 49952 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2222_
timestamp 1669390400
transform -1 0 49728 0 1 26656
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2223_
timestamp 1669390400
transform 1 0 52640 0 -1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2224_
timestamp 1669390400
transform 1 0 53536 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2225_
timestamp 1669390400
transform 1 0 53312 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2226_
timestamp 1669390400
transform -1 0 52416 0 1 12544
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2227_
timestamp 1669390400
transform 1 0 46480 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2228_
timestamp 1669390400
transform 1 0 43904 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2229_
timestamp 1669390400
transform -1 0 47376 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2230_
timestamp 1669390400
transform 1 0 47824 0 -1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2231_
timestamp 1669390400
transform -1 0 54432 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2232_
timestamp 1669390400
transform -1 0 53312 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2233_
timestamp 1669390400
transform -1 0 52752 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2234_
timestamp 1669390400
transform -1 0 50960 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2235_
timestamp 1669390400
transform 1 0 49616 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2236_
timestamp 1669390400
transform -1 0 52864 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2237_
timestamp 1669390400
transform -1 0 51632 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2238_
timestamp 1669390400
transform -1 0 51968 0 -1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2239_
timestamp 1669390400
transform 1 0 53312 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2240_
timestamp 1669390400
transform -1 0 51744 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2241_
timestamp 1669390400
transform -1 0 51072 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2242_
timestamp 1669390400
transform 1 0 48944 0 1 6272
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2243_
timestamp 1669390400
transform -1 0 53984 0 -1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2244_
timestamp 1669390400
transform -1 0 49952 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2245_
timestamp 1669390400
transform -1 0 50064 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2246_
timestamp 1669390400
transform 1 0 47824 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2247_
timestamp 1669390400
transform -1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2248_
timestamp 1669390400
transform -1 0 27664 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2249_
timestamp 1669390400
transform -1 0 26880 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2250_
timestamp 1669390400
transform 1 0 27104 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2251_
timestamp 1669390400
transform -1 0 46704 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2252_
timestamp 1669390400
transform -1 0 53536 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2253_
timestamp 1669390400
transform -1 0 41664 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2254_
timestamp 1669390400
transform -1 0 48720 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2255_
timestamp 1669390400
transform 1 0 47488 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2256_
timestamp 1669390400
transform -1 0 43456 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2257_
timestamp 1669390400
transform 1 0 42336 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2258_
timestamp 1669390400
transform 1 0 41216 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2259_
timestamp 1669390400
transform -1 0 51856 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2260_
timestamp 1669390400
transform 1 0 42896 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2261_
timestamp 1669390400
transform -1 0 46816 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2262_
timestamp 1669390400
transform -1 0 46480 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2263_
timestamp 1669390400
transform 1 0 43456 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2264_
timestamp 1669390400
transform 1 0 42224 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2265_
timestamp 1669390400
transform 1 0 43792 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2266_
timestamp 1669390400
transform -1 0 51184 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2267_
timestamp 1669390400
transform -1 0 43232 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2268_
timestamp 1669390400
transform 1 0 41776 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2269_
timestamp 1669390400
transform 1 0 44016 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2270_
timestamp 1669390400
transform 1 0 44240 0 -1 12544
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2271_
timestamp 1669390400
transform 1 0 30912 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2272_
timestamp 1669390400
transform 1 0 29344 0 -1 9408
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2273_
timestamp 1669390400
transform -1 0 31024 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2274_
timestamp 1669390400
transform 1 0 50400 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2275_
timestamp 1669390400
transform -1 0 56896 0 -1 18816
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2276_
timestamp 1669390400
transform -1 0 52864 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2277_
timestamp 1669390400
transform -1 0 49168 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2278_
timestamp 1669390400
transform 1 0 48160 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2279_
timestamp 1669390400
transform 1 0 49392 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2280_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 58016 0 1 20384
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2281_
timestamp 1669390400
transform -1 0 57680 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2282_
timestamp 1669390400
transform -1 0 51968 0 -1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2283_
timestamp 1669390400
transform -1 0 51408 0 -1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2284_
timestamp 1669390400
transform -1 0 46256 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2285_
timestamp 1669390400
transform -1 0 47264 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2286_
timestamp 1669390400
transform -1 0 50736 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2287_
timestamp 1669390400
transform 1 0 56000 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2288_
timestamp 1669390400
transform 1 0 55440 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2289_
timestamp 1669390400
transform 1 0 46704 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2290_
timestamp 1669390400
transform 1 0 49952 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2291_
timestamp 1669390400
transform -1 0 52080 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2292_
timestamp 1669390400
transform 1 0 50512 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2293_
timestamp 1669390400
transform 1 0 51744 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2294_
timestamp 1669390400
transform 1 0 41552 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2295_
timestamp 1669390400
transform -1 0 42896 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2296_
timestamp 1669390400
transform 1 0 49392 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2297_
timestamp 1669390400
transform 1 0 50960 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2298_
timestamp 1669390400
transform -1 0 50848 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2299_
timestamp 1669390400
transform -1 0 36400 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2300_
timestamp 1669390400
transform -1 0 36736 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2301_
timestamp 1669390400
transform 1 0 34944 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2302_
timestamp 1669390400
transform -1 0 34384 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2303_
timestamp 1669390400
transform 1 0 30464 0 -1 6272
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2304_
timestamp 1669390400
transform -1 0 33040 0 -1 4704
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2305_
timestamp 1669390400
transform -1 0 26880 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2306_
timestamp 1669390400
transform 1 0 31248 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2307_
timestamp 1669390400
transform 1 0 27104 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2308_
timestamp 1669390400
transform -1 0 32368 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2309_
timestamp 1669390400
transform 1 0 32704 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2310_
timestamp 1669390400
transform -1 0 33376 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2311_
timestamp 1669390400
transform -1 0 35840 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2312_
timestamp 1669390400
transform -1 0 31696 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2313_
timestamp 1669390400
transform -1 0 32592 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2314_
timestamp 1669390400
transform -1 0 40880 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2315_
timestamp 1669390400
transform -1 0 40096 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2316_
timestamp 1669390400
transform 1 0 39200 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2317_
timestamp 1669390400
transform -1 0 42560 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2318_
timestamp 1669390400
transform 1 0 40096 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2319_
timestamp 1669390400
transform -1 0 43232 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2320_
timestamp 1669390400
transform -1 0 40208 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2321_
timestamp 1669390400
transform 1 0 38864 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2322_
timestamp 1669390400
transform -1 0 38752 0 -1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2323_
timestamp 1669390400
transform -1 0 34160 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2324_
timestamp 1669390400
transform -1 0 38080 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2325_
timestamp 1669390400
transform 1 0 31808 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2326_
timestamp 1669390400
transform -1 0 42112 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2327_
timestamp 1669390400
transform 1 0 40992 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2328_
timestamp 1669390400
transform 1 0 41888 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2329_
timestamp 1669390400
transform 1 0 41552 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2330_
timestamp 1669390400
transform -1 0 43120 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2331_
timestamp 1669390400
transform 1 0 42336 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2332_
timestamp 1669390400
transform -1 0 43568 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2333_
timestamp 1669390400
transform 1 0 42448 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2334_
timestamp 1669390400
transform -1 0 33376 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2335_
timestamp 1669390400
transform 1 0 32256 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2336_
timestamp 1669390400
transform 1 0 30912 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2337_
timestamp 1669390400
transform -1 0 26432 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2338_
timestamp 1669390400
transform 1 0 24976 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2339_
timestamp 1669390400
transform -1 0 26768 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2340_
timestamp 1669390400
transform 1 0 25760 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2341_
timestamp 1669390400
transform 1 0 26544 0 1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2342_
timestamp 1669390400
transform -1 0 48272 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2343_
timestamp 1669390400
transform -1 0 44016 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2344_
timestamp 1669390400
transform -1 0 31584 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2345_
timestamp 1669390400
transform -1 0 50960 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2346_
timestamp 1669390400
transform -1 0 47824 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2347_
timestamp 1669390400
transform -1 0 46144 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2348_
timestamp 1669390400
transform 1 0 45360 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2349_
timestamp 1669390400
transform -1 0 48608 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2350_
timestamp 1669390400
transform -1 0 46368 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2351_
timestamp 1669390400
transform 1 0 46144 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2352_
timestamp 1669390400
transform -1 0 46256 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2353_
timestamp 1669390400
transform -1 0 47824 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2354_
timestamp 1669390400
transform -1 0 47040 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2355_
timestamp 1669390400
transform -1 0 46256 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2356_
timestamp 1669390400
transform -1 0 42224 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2357_
timestamp 1669390400
transform -1 0 43120 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2358_
timestamp 1669390400
transform 1 0 42560 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2359_
timestamp 1669390400
transform 1 0 42448 0 -1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2360_
timestamp 1669390400
transform 1 0 35280 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2361_
timestamp 1669390400
transform 1 0 45584 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2362_
timestamp 1669390400
transform -1 0 46928 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2363_
timestamp 1669390400
transform 1 0 45584 0 1 17248
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2364_
timestamp 1669390400
transform -1 0 46480 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2365_
timestamp 1669390400
transform 1 0 44912 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2366_
timestamp 1669390400
transform -1 0 47824 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2367_
timestamp 1669390400
transform 1 0 46032 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2368_
timestamp 1669390400
transform 1 0 46144 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2369_
timestamp 1669390400
transform 1 0 45696 0 -1 21952
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2370_
timestamp 1669390400
transform 1 0 44912 0 -1 20384
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2371_
timestamp 1669390400
transform -1 0 50848 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2372_
timestamp 1669390400
transform -1 0 24640 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2373_
timestamp 1669390400
transform 1 0 23856 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2374_
timestamp 1669390400
transform -1 0 26880 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2375_
timestamp 1669390400
transform 1 0 26320 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2376_
timestamp 1669390400
transform 1 0 27552 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2377_
timestamp 1669390400
transform 1 0 29120 0 1 3136
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2378_
timestamp 1669390400
transform 1 0 30128 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2379_
timestamp 1669390400
transform -1 0 36736 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2380_
timestamp 1669390400
transform -1 0 40992 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2381_
timestamp 1669390400
transform 1 0 41664 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2382_
timestamp 1669390400
transform 1 0 46368 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2383_
timestamp 1669390400
transform -1 0 48160 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2384_
timestamp 1669390400
transform -1 0 36960 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2385_
timestamp 1669390400
transform -1 0 43792 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2386_
timestamp 1669390400
transform -1 0 44576 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2387_
timestamp 1669390400
transform -1 0 44464 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2388_
timestamp 1669390400
transform -1 0 36512 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2389_
timestamp 1669390400
transform 1 0 31360 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2390_
timestamp 1669390400
transform -1 0 31696 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2391_
timestamp 1669390400
transform -1 0 32368 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2392_
timestamp 1669390400
transform -1 0 28000 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2393_
timestamp 1669390400
transform 1 0 23968 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2394_
timestamp 1669390400
transform 1 0 40880 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2395_
timestamp 1669390400
transform 1 0 39872 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2396_
timestamp 1669390400
transform -1 0 40768 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2397_
timestamp 1669390400
transform 1 0 38640 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2398_
timestamp 1669390400
transform 1 0 39088 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2399_
timestamp 1669390400
transform -1 0 41664 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2400_
timestamp 1669390400
transform 1 0 39760 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2401_
timestamp 1669390400
transform -1 0 45920 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2402_
timestamp 1669390400
transform 1 0 40096 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2403_
timestamp 1669390400
transform -1 0 46368 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2404_
timestamp 1669390400
transform -1 0 42336 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2405_
timestamp 1669390400
transform -1 0 42112 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2406_
timestamp 1669390400
transform -1 0 39648 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2407_
timestamp 1669390400
transform -1 0 39536 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2408_
timestamp 1669390400
transform 1 0 39088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2409_
timestamp 1669390400
transform -1 0 24304 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2410_
timestamp 1669390400
transform -1 0 23520 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2411_
timestamp 1669390400
transform 1 0 29456 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2412_
timestamp 1669390400
transform -1 0 42112 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2413_
timestamp 1669390400
transform -1 0 41440 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2414_
timestamp 1669390400
transform -1 0 40656 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2415_
timestamp 1669390400
transform 1 0 39760 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2416_
timestamp 1669390400
transform -1 0 40992 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2417_
timestamp 1669390400
transform -1 0 48384 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2418_
timestamp 1669390400
transform 1 0 29792 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2419_
timestamp 1669390400
transform 1 0 29792 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2420_
timestamp 1669390400
transform -1 0 22960 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2421_
timestamp 1669390400
transform 1 0 21280 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2422_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 23296 0 -1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2423_
timestamp 1669390400
transform 1 0 25648 0 1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2424_
timestamp 1669390400
transform -1 0 26432 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _2425_
timestamp 1669390400
transform -1 0 23520 0 1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2426_
timestamp 1669390400
transform 1 0 28000 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2427_
timestamp 1669390400
transform 1 0 28224 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2428_
timestamp 1669390400
transform 1 0 20944 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2429_
timestamp 1669390400
transform 1 0 21952 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2430_
timestamp 1669390400
transform -1 0 21056 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2431_
timestamp 1669390400
transform 1 0 21504 0 1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2432_
timestamp 1669390400
transform 1 0 24416 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2433_
timestamp 1669390400
transform -1 0 43456 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2434_
timestamp 1669390400
transform 1 0 42224 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2435_
timestamp 1669390400
transform -1 0 38080 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2436_
timestamp 1669390400
transform -1 0 39312 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2437_
timestamp 1669390400
transform -1 0 38304 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2438_
timestamp 1669390400
transform 1 0 38528 0 1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2439_
timestamp 1669390400
transform 1 0 42560 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2440_
timestamp 1669390400
transform 1 0 37744 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2441_
timestamp 1669390400
transform 1 0 38528 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2442_
timestamp 1669390400
transform -1 0 30016 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2443_
timestamp 1669390400
transform 1 0 26544 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2444_
timestamp 1669390400
transform -1 0 25984 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2445_
timestamp 1669390400
transform 1 0 36064 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2446_
timestamp 1669390400
transform 1 0 29680 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2447_
timestamp 1669390400
transform -1 0 32368 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2448_
timestamp 1669390400
transform -1 0 32256 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2449_
timestamp 1669390400
transform 1 0 31248 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2450_
timestamp 1669390400
transform 1 0 36288 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2451_
timestamp 1669390400
transform 1 0 49392 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2452_
timestamp 1669390400
transform -1 0 42560 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2453_
timestamp 1669390400
transform -1 0 44576 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2454_
timestamp 1669390400
transform 1 0 40656 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2455_
timestamp 1669390400
transform 1 0 40656 0 1 17248
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2456_
timestamp 1669390400
transform 1 0 39088 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2457_
timestamp 1669390400
transform 1 0 36288 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2458_
timestamp 1669390400
transform 1 0 37408 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2459_
timestamp 1669390400
transform -1 0 38864 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2460_
timestamp 1669390400
transform -1 0 39088 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2461_
timestamp 1669390400
transform -1 0 37968 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2462_
timestamp 1669390400
transform 1 0 23184 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2463_
timestamp 1669390400
transform 1 0 38864 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2464_
timestamp 1669390400
transform 1 0 36736 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2465_
timestamp 1669390400
transform -1 0 44576 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2466_
timestamp 1669390400
transform -1 0 44576 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2467_
timestamp 1669390400
transform -1 0 36288 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2468_
timestamp 1669390400
transform -1 0 36512 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2469_
timestamp 1669390400
transform -1 0 22960 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_2  _2470_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 21056 0 -1 15680
box -86 -86 3222 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2471_
timestamp 1669390400
transform 1 0 20160 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2472_
timestamp 1669390400
transform -1 0 22400 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2473_
timestamp 1669390400
transform -1 0 20720 0 -1 18816
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2474_
timestamp 1669390400
transform -1 0 2912 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2475_
timestamp 1669390400
transform 1 0 31248 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2476_
timestamp 1669390400
transform 1 0 31248 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2477_
timestamp 1669390400
transform -1 0 36960 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2478_
timestamp 1669390400
transform -1 0 41440 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2479_
timestamp 1669390400
transform -1 0 38864 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2480_
timestamp 1669390400
transform 1 0 36512 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2481_
timestamp 1669390400
transform 1 0 37408 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2482_
timestamp 1669390400
transform 1 0 33600 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2483_
timestamp 1669390400
transform -1 0 44576 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2484_
timestamp 1669390400
transform 1 0 31696 0 -1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2485_
timestamp 1669390400
transform 1 0 33488 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2486_
timestamp 1669390400
transform -1 0 30128 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2487_
timestamp 1669390400
transform -1 0 29008 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2488_
timestamp 1669390400
transform -1 0 29008 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2489_
timestamp 1669390400
transform -1 0 26432 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2490_
timestamp 1669390400
transform -1 0 36288 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2491_
timestamp 1669390400
transform -1 0 34496 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2492_
timestamp 1669390400
transform -1 0 38192 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2493_
timestamp 1669390400
transform -1 0 37968 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2494_
timestamp 1669390400
transform -1 0 35392 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2495_
timestamp 1669390400
transform -1 0 36512 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2496_
timestamp 1669390400
transform 1 0 33936 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2497_
timestamp 1669390400
transform -1 0 36064 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _2498_
timestamp 1669390400
transform 1 0 35056 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2499_
timestamp 1669390400
transform 1 0 36400 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2500_
timestamp 1669390400
transform -1 0 35616 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2501_
timestamp 1669390400
transform 1 0 39872 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2502_
timestamp 1669390400
transform -1 0 41664 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2503_
timestamp 1669390400
transform -1 0 36512 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2504_
timestamp 1669390400
transform -1 0 36288 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2505_
timestamp 1669390400
transform -1 0 43120 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2506_
timestamp 1669390400
transform -1 0 36288 0 -1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2507_
timestamp 1669390400
transform 1 0 34608 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2508_
timestamp 1669390400
transform -1 0 30016 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2509_
timestamp 1669390400
transform 1 0 27888 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2510_
timestamp 1669390400
transform -1 0 28896 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2511_
timestamp 1669390400
transform -1 0 26320 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2512_
timestamp 1669390400
transform -1 0 29680 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2513_
timestamp 1669390400
transform 1 0 34272 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2514_
timestamp 1669390400
transform 1 0 38416 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2515_
timestamp 1669390400
transform 1 0 34384 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2516_
timestamp 1669390400
transform -1 0 40992 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2517_
timestamp 1669390400
transform -1 0 37856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2518_
timestamp 1669390400
transform 1 0 35728 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2519_
timestamp 1669390400
transform 1 0 23520 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2520_
timestamp 1669390400
transform 1 0 13776 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2521_
timestamp 1669390400
transform -1 0 19488 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2522_
timestamp 1669390400
transform 1 0 18816 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2523_
timestamp 1669390400
transform 1 0 18592 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2524_
timestamp 1669390400
transform 1 0 15344 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2525_
timestamp 1669390400
transform 1 0 18256 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _2526_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 19824 0 -1 17248
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2527_
timestamp 1669390400
transform -1 0 18032 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2528_
timestamp 1669390400
transform 1 0 15680 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2529_
timestamp 1669390400
transform -1 0 57680 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2530_
timestamp 1669390400
transform 1 0 14560 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2531_
timestamp 1669390400
transform -1 0 16352 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2532_
timestamp 1669390400
transform -1 0 15120 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2533_
timestamp 1669390400
transform -1 0 31696 0 -1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2534_
timestamp 1669390400
transform -1 0 30128 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2535_
timestamp 1669390400
transform -1 0 28448 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2536_
timestamp 1669390400
transform -1 0 40320 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2537_
timestamp 1669390400
transform 1 0 37968 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2538_
timestamp 1669390400
transform -1 0 39424 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2539_
timestamp 1669390400
transform -1 0 39424 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2540_
timestamp 1669390400
transform 1 0 36848 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2541_
timestamp 1669390400
transform 1 0 37632 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2542_
timestamp 1669390400
transform -1 0 34160 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2543_
timestamp 1669390400
transform 1 0 30688 0 1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2544_
timestamp 1669390400
transform 1 0 32256 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2545_
timestamp 1669390400
transform 1 0 31360 0 1 23520
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2546_
timestamp 1669390400
transform 1 0 28672 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2547_
timestamp 1669390400
transform 1 0 28112 0 -1 14112
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2548_
timestamp 1669390400
transform 1 0 28336 0 -1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2549_
timestamp 1669390400
transform -1 0 38528 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2550_
timestamp 1669390400
transform -1 0 35840 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2551_
timestamp 1669390400
transform -1 0 35056 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2552_
timestamp 1669390400
transform 1 0 34160 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2553_
timestamp 1669390400
transform 1 0 34720 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2554_
timestamp 1669390400
transform 1 0 34160 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2555_
timestamp 1669390400
transform 1 0 34608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2556_
timestamp 1669390400
transform -1 0 36512 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2557_
timestamp 1669390400
transform -1 0 23408 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2558_
timestamp 1669390400
transform 1 0 30464 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2559_
timestamp 1669390400
transform -1 0 36288 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2560_
timestamp 1669390400
transform 1 0 34496 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2561_
timestamp 1669390400
transform -1 0 32368 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2562_
timestamp 1669390400
transform -1 0 32256 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2563_
timestamp 1669390400
transform -1 0 24976 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2564_
timestamp 1669390400
transform -1 0 23632 0 1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2565_
timestamp 1669390400
transform -1 0 23184 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2566_
timestamp 1669390400
transform 1 0 15008 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2567_
timestamp 1669390400
transform 1 0 14896 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2568_
timestamp 1669390400
transform -1 0 17024 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2569_
timestamp 1669390400
transform -1 0 17360 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2570_
timestamp 1669390400
transform 1 0 14560 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2571_
timestamp 1669390400
transform 1 0 15904 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2572_
timestamp 1669390400
transform -1 0 15680 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2573_
timestamp 1669390400
transform -1 0 2912 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2574_
timestamp 1669390400
transform 1 0 27552 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2575_
timestamp 1669390400
transform 1 0 37632 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2576_
timestamp 1669390400
transform -1 0 39536 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2577_
timestamp 1669390400
transform -1 0 39200 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2578_
timestamp 1669390400
transform -1 0 39088 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2579_
timestamp 1669390400
transform 1 0 27440 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2580_
timestamp 1669390400
transform -1 0 27216 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2581_
timestamp 1669390400
transform 1 0 27104 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2582_
timestamp 1669390400
transform -1 0 38304 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2583_
timestamp 1669390400
transform -1 0 36064 0 1 26656
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2584_
timestamp 1669390400
transform -1 0 27664 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2585_
timestamp 1669390400
transform 1 0 26320 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2586_
timestamp 1669390400
transform 1 0 34384 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2587_
timestamp 1669390400
transform -1 0 36960 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2588_
timestamp 1669390400
transform 1 0 34832 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2589_
timestamp 1669390400
transform -1 0 36512 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2590_
timestamp 1669390400
transform 1 0 35728 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2591_
timestamp 1669390400
transform -1 0 37632 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2592_
timestamp 1669390400
transform -1 0 21504 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2593_
timestamp 1669390400
transform -1 0 19936 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2594_
timestamp 1669390400
transform -1 0 18480 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2595_
timestamp 1669390400
transform 1 0 23856 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2596_
timestamp 1669390400
transform -1 0 24528 0 -1 10976
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2597_
timestamp 1669390400
transform -1 0 16800 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2598_
timestamp 1669390400
transform -1 0 16688 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2599_
timestamp 1669390400
transform 1 0 15344 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2600_
timestamp 1669390400
transform 1 0 15120 0 -1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2601_
timestamp 1669390400
transform -1 0 15232 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2602_
timestamp 1669390400
transform -1 0 15120 0 1 9408
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2603_
timestamp 1669390400
transform -1 0 13216 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2604_
timestamp 1669390400
transform -1 0 20160 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2605_
timestamp 1669390400
transform 1 0 18816 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2606_
timestamp 1669390400
transform -1 0 29568 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2607_
timestamp 1669390400
transform -1 0 33936 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2608_
timestamp 1669390400
transform 1 0 33600 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2609_
timestamp 1669390400
transform -1 0 34160 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2610_
timestamp 1669390400
transform 1 0 29456 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2611_
timestamp 1669390400
transform -1 0 30016 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2612_
timestamp 1669390400
transform -1 0 29008 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2613_
timestamp 1669390400
transform -1 0 29120 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2614_
timestamp 1669390400
transform 1 0 28112 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2615_
timestamp 1669390400
transform -1 0 28336 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2616_
timestamp 1669390400
transform -1 0 33824 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2617_
timestamp 1669390400
transform -1 0 34160 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2618_
timestamp 1669390400
transform -1 0 35392 0 -1 15680
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2619_
timestamp 1669390400
transform -1 0 35728 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2620_
timestamp 1669390400
transform -1 0 35616 0 1 7840
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2621_
timestamp 1669390400
transform -1 0 31584 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2622_
timestamp 1669390400
transform -1 0 26096 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2623_
timestamp 1669390400
transform 1 0 23744 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2624_
timestamp 1669390400
transform -1 0 21504 0 -1 9408
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2625_
timestamp 1669390400
transform 1 0 19040 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2626_
timestamp 1669390400
transform -1 0 20160 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2627_
timestamp 1669390400
transform -1 0 18032 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2628_
timestamp 1669390400
transform -1 0 17136 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2629_
timestamp 1669390400
transform -1 0 16352 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2630_
timestamp 1669390400
transform -1 0 16240 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2631_
timestamp 1669390400
transform -1 0 15456 0 1 10976
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2632_
timestamp 1669390400
transform 1 0 2240 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2633_
timestamp 1669390400
transform -1 0 34384 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2634_
timestamp 1669390400
transform -1 0 34160 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _2635_
timestamp 1669390400
transform -1 0 34608 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2636_
timestamp 1669390400
transform -1 0 33488 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2637_
timestamp 1669390400
transform 1 0 25536 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2638_
timestamp 1669390400
transform 1 0 24864 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2639_
timestamp 1669390400
transform -1 0 26320 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2640_
timestamp 1669390400
transform -1 0 25984 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2641_
timestamp 1669390400
transform -1 0 25648 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2642_
timestamp 1669390400
transform -1 0 23968 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2643_
timestamp 1669390400
transform 1 0 29456 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2644_
timestamp 1669390400
transform 1 0 31696 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2645_
timestamp 1669390400
transform 1 0 31808 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2646_
timestamp 1669390400
transform -1 0 30800 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2647_
timestamp 1669390400
transform -1 0 29568 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2648_
timestamp 1669390400
transform -1 0 22624 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2649_
timestamp 1669390400
transform -1 0 22400 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2650_
timestamp 1669390400
transform -1 0 20832 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2651_
timestamp 1669390400
transform -1 0 20832 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2652_
timestamp 1669390400
transform -1 0 20384 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2653_
timestamp 1669390400
transform 1 0 17584 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2654_
timestamp 1669390400
transform 1 0 17584 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2655_
timestamp 1669390400
transform -1 0 17696 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2656_
timestamp 1669390400
transform -1 0 2912 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2657_
timestamp 1669390400
transform -1 0 25088 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2658_
timestamp 1669390400
transform 1 0 22736 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2659_
timestamp 1669390400
transform 1 0 31248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2660_
timestamp 1669390400
transform -1 0 27776 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2661_
timestamp 1669390400
transform 1 0 26544 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2662_
timestamp 1669390400
transform -1 0 26768 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2663_
timestamp 1669390400
transform 1 0 26544 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2664_
timestamp 1669390400
transform -1 0 24192 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2665_
timestamp 1669390400
transform 1 0 20272 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2666_
timestamp 1669390400
transform 1 0 17920 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2667_
timestamp 1669390400
transform 1 0 20384 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2668_
timestamp 1669390400
transform 1 0 21392 0 -1 4704
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2669_
timestamp 1669390400
transform -1 0 58016 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2670_
timestamp 1669390400
transform -1 0 22624 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2671_
timestamp 1669390400
transform 1 0 21504 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2672_
timestamp 1669390400
transform -1 0 28672 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2673_
timestamp 1669390400
transform 1 0 23856 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2674_
timestamp 1669390400
transform -1 0 24528 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2675_
timestamp 1669390400
transform 1 0 24192 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2676_
timestamp 1669390400
transform -1 0 25648 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2677_
timestamp 1669390400
transform 1 0 51520 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2678_
timestamp 1669390400
transform 1 0 53312 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2679_
timestamp 1669390400
transform -1 0 57680 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2680_
timestamp 1669390400
transform 1 0 32480 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2681_
timestamp 1669390400
transform 1 0 33712 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2682_
timestamp 1669390400
transform 1 0 29456 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2683_
timestamp 1669390400
transform 1 0 23072 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2684_
timestamp 1669390400
transform -1 0 15792 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2685_
timestamp 1669390400
transform -1 0 19712 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2686_
timestamp 1669390400
transform -1 0 19264 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2687_
timestamp 1669390400
transform 1 0 26880 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2688_
timestamp 1669390400
transform 1 0 34944 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2689_
timestamp 1669390400
transform 1 0 35728 0 1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2690_
timestamp 1669390400
transform -1 0 35728 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2691_
timestamp 1669390400
transform 1 0 36288 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2692_
timestamp 1669390400
transform -1 0 37968 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2693_
timestamp 1669390400
transform 1 0 30352 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2694_
timestamp 1669390400
transform -1 0 31472 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2695_
timestamp 1669390400
transform 1 0 28000 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2696_
timestamp 1669390400
transform 1 0 27440 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2697_
timestamp 1669390400
transform 1 0 31696 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2698_
timestamp 1669390400
transform -1 0 35392 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2699_
timestamp 1669390400
transform -1 0 32480 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2700_
timestamp 1669390400
transform 1 0 33600 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2701_
timestamp 1669390400
transform 1 0 31360 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2702_
timestamp 1669390400
transform 1 0 32704 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2703_
timestamp 1669390400
transform 1 0 13664 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2704_
timestamp 1669390400
transform -1 0 15904 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2705_
timestamp 1669390400
transform -1 0 20720 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2706_
timestamp 1669390400
transform -1 0 19936 0 1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2707_
timestamp 1669390400
transform -1 0 17360 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2708_
timestamp 1669390400
transform 1 0 14896 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2709_
timestamp 1669390400
transform -1 0 15120 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2710_
timestamp 1669390400
transform -1 0 14896 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2711_
timestamp 1669390400
transform -1 0 12096 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2712_
timestamp 1669390400
transform 1 0 10864 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2713_
timestamp 1669390400
transform -1 0 22960 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2714_
timestamp 1669390400
transform -1 0 23072 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2715_
timestamp 1669390400
transform 1 0 18480 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2716_
timestamp 1669390400
transform 1 0 19376 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2717_
timestamp 1669390400
transform 1 0 22512 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2718_
timestamp 1669390400
transform 1 0 22400 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2719_
timestamp 1669390400
transform 1 0 23184 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2720_
timestamp 1669390400
transform -1 0 37968 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2721_
timestamp 1669390400
transform 1 0 39200 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2722_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 33488 0 -1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2723_
timestamp 1669390400
transform 1 0 33152 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2724_
timestamp 1669390400
transform 1 0 21056 0 -1 28224
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2725_
timestamp 1669390400
transform 1 0 21280 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2726_
timestamp 1669390400
transform 1 0 17248 0 1 25088
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2727_
timestamp 1669390400
transform 1 0 25536 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2728_
timestamp 1669390400
transform 1 0 38192 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _2729_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 22288 0 -1 25088
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2730_
timestamp 1669390400
transform 1 0 17248 0 1 23520
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2731_
timestamp 1669390400
transform 1 0 37408 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2732_
timestamp 1669390400
transform 1 0 37184 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2733_
timestamp 1669390400
transform -1 0 30688 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2734_
timestamp 1669390400
transform 1 0 39872 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2735_
timestamp 1669390400
transform 1 0 39872 0 1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2736_
timestamp 1669390400
transform 1 0 34272 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2737_
timestamp 1669390400
transform 1 0 25200 0 1 32928
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _2738_
timestamp 1669390400
transform 1 0 29792 0 -1 32928
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _2739_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 13776 0 1 28224
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2740_
timestamp 1669390400
transform 1 0 18592 0 -1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2741_
timestamp 1669390400
transform 1 0 13328 0 -1 26656
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _2742_
timestamp 1669390400
transform -1 0 14224 0 -1 28224
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffsnq_1  _2743_
timestamp 1669390400
transform 1 0 18144 0 -1 31360
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2744_
timestamp 1669390400
transform 1 0 23296 0 1 29792
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2745_
timestamp 1669390400
transform 1 0 27552 0 -1 31360
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2746_
timestamp 1669390400
transform 1 0 38192 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2747_
timestamp 1669390400
transform 1 0 37184 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  fanout44 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 29008 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  fanout45 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 26768 0 1 23520
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  fanout46
timestamp 1669390400
transform 1 0 34160 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  fanout47
timestamp 1669390400
transform 1 0 24416 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout48
timestamp 1669390400
transform -1 0 26208 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  fanout49
timestamp 1669390400
transform 1 0 33824 0 -1 34496
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  fanout50
timestamp 1669390400
transform -1 0 24304 0 1 34496
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  fanout51
timestamp 1669390400
transform -1 0 13664 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout52
timestamp 1669390400
transform -1 0 22176 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout53
timestamp 1669390400
transform 1 0 24416 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  fanout54
timestamp 1669390400
transform 1 0 21056 0 -1 23520
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout55
timestamp 1669390400
transform -1 0 15120 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout56
timestamp 1669390400
transform -1 0 36960 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  fanout57
timestamp 1669390400
transform 1 0 42112 0 1 32928
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  fanout58
timestamp 1669390400
transform 1 0 36848 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout59
timestamp 1669390400
transform -1 0 29904 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout60
timestamp 1669390400
transform 1 0 38304 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  fanout61
timestamp 1669390400
transform -1 0 31920 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  fanout62
timestamp 1669390400
transform 1 0 13552 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout63
timestamp 1669390400
transform -1 0 14896 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  fanout64
timestamp 1669390400
transform 1 0 18256 0 -1 25088
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  fanout65
timestamp 1669390400
transform -1 0 40880 0 1 29792
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  fanout66
timestamp 1669390400
transform 1 0 37856 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  fanout67
timestamp 1669390400
transform -1 0 40768 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  fanout68
timestamp 1669390400
transform -1 0 43232 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1
timestamp 1669390400
transform -1 0 30912 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2
timestamp 1669390400
transform 1 0 1680 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input3
timestamp 1669390400
transform -1 0 45472 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input4
timestamp 1669390400
transform -1 0 56560 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input5
timestamp 1669390400
transform 1 0 5600 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output6 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 56336 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output7
timestamp 1669390400
transform -1 0 3248 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output8
timestamp 1669390400
transform -1 0 56112 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output9
timestamp 1669390400
transform 1 0 54768 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output10
timestamp 1669390400
transform -1 0 56336 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output11
timestamp 1669390400
transform -1 0 23856 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output12
timestamp 1669390400
transform 1 0 33712 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output13
timestamp 1669390400
transform 1 0 46480 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output14
timestamp 1669390400
transform -1 0 3248 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output15
timestamp 1669390400
transform -1 0 56336 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output16
timestamp 1669390400
transform -1 0 3248 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output17
timestamp 1669390400
transform -1 0 12432 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output18
timestamp 1669390400
transform -1 0 3248 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output19
timestamp 1669390400
transform -1 0 3248 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output20
timestamp 1669390400
transform -1 0 36512 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output21
timestamp 1669390400
transform 1 0 52640 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output22
timestamp 1669390400
transform 1 0 54768 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output23
timestamp 1669390400
transform 1 0 54768 0 1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output24
timestamp 1669390400
transform -1 0 12992 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output25
timestamp 1669390400
transform -1 0 3248 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output26
timestamp 1669390400
transform -1 0 3248 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output27
timestamp 1669390400
transform 1 0 54768 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output28
timestamp 1669390400
transform 1 0 6832 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output29
timestamp 1669390400
transform -1 0 3248 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output30
timestamp 1669390400
transform 1 0 50512 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output31
timestamp 1669390400
transform -1 0 42448 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output32
timestamp 1669390400
transform -1 0 18928 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output33
timestamp 1669390400
transform -1 0 3248 0 1 50176
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output34
timestamp 1669390400
transform 1 0 54768 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output35
timestamp 1669390400
transform -1 0 28672 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output36
timestamp 1669390400
transform 1 0 54544 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output37
timestamp 1669390400
transform 1 0 54768 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output38
timestamp 1669390400
transform 1 0 18256 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output39
timestamp 1669390400
transform -1 0 24752 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output40
timestamp 1669390400
transform -1 0 40432 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output41
timestamp 1669390400
transform -1 0 3248 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output42
timestamp 1669390400
transform -1 0 3248 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output43
timestamp 1669390400
transform 1 0 54768 0 -1 29792
box -86 -86 1654 870
<< labels >>
flabel metal2 s 28896 59200 29008 59800 0 FreeSans 448 90 0 0 ACK
port 0 nsew signal input
flabel metal2 s 1344 59200 1456 59800 0 FreeSans 448 90 0 0 Bit_In
port 1 nsew signal input
flabel metal2 s 44352 200 44464 800 0 FreeSans 448 90 0 0 EN
port 2 nsew signal input
flabel metal3 s 59200 6720 59800 6832 0 FreeSans 448 0 0 0 I[0]
port 3 nsew signal tristate
flabel metal3 s 200 44352 800 44464 0 FreeSans 448 0 0 0 I[10]
port 4 nsew signal tristate
flabel metal3 s 59200 1344 59800 1456 0 FreeSans 448 0 0 0 I[11]
port 5 nsew signal tristate
flabel metal2 s 55776 200 55888 800 0 FreeSans 448 90 0 0 I[12]
port 6 nsew signal tristate
flabel metal3 s 59200 40320 59800 40432 0 FreeSans 448 0 0 0 I[1]
port 7 nsew signal tristate
flabel metal2 s 22176 200 22288 800 0 FreeSans 448 90 0 0 I[2]
port 8 nsew signal tristate
flabel metal2 s 33600 200 33712 800 0 FreeSans 448 90 0 0 I[3]
port 9 nsew signal tristate
flabel metal2 s 46368 59200 46480 59800 0 FreeSans 448 90 0 0 I[4]
port 10 nsew signal tristate
flabel metal3 s 200 22176 800 22288 0 FreeSans 448 0 0 0 I[5]
port 11 nsew signal tristate
flabel metal3 s 59200 46368 59800 46480 0 FreeSans 448 0 0 0 I[6]
port 12 nsew signal tristate
flabel metal3 s 200 33600 800 33712 0 FreeSans 448 0 0 0 I[7]
port 13 nsew signal tristate
flabel metal2 s 10752 200 10864 800 0 FreeSans 448 90 0 0 I[8]
port 14 nsew signal tristate
flabel metal3 s 200 38976 800 39088 0 FreeSans 448 0 0 0 I[9]
port 15 nsew signal tristate
flabel metal3 s 200 16800 800 16912 0 FreeSans 448 0 0 0 Q[0]
port 16 nsew signal tristate
flabel metal2 s 34944 59200 35056 59800 0 FreeSans 448 90 0 0 Q[10]
port 17 nsew signal tristate
flabel metal2 s 51744 59200 51856 59800 0 FreeSans 448 90 0 0 Q[11]
port 18 nsew signal tristate
flabel metal3 s 59200 18144 59800 18256 0 FreeSans 448 0 0 0 Q[12]
port 19 nsew signal tristate
flabel metal3 s 59200 51744 59800 51856 0 FreeSans 448 0 0 0 Q[1]
port 20 nsew signal tristate
flabel metal2 s 12096 59200 12208 59800 0 FreeSans 448 90 0 0 Q[2]
port 21 nsew signal tristate
flabel metal2 s 0 200 112 800 0 FreeSans 448 90 0 0 Q[3]
port 22 nsew signal tristate
flabel metal3 s 200 10752 800 10864 0 FreeSans 448 0 0 0 Q[4]
port 23 nsew signal tristate
flabel metal3 s 59200 34944 59800 35056 0 FreeSans 448 0 0 0 Q[5]
port 24 nsew signal tristate
flabel metal2 s 6720 59200 6832 59800 0 FreeSans 448 90 0 0 Q[6]
port 25 nsew signal tristate
flabel metal3 s 200 5376 800 5488 0 FreeSans 448 0 0 0 Q[7]
port 26 nsew signal tristate
flabel metal2 s 50400 200 50512 800 0 FreeSans 448 90 0 0 Q[8]
port 27 nsew signal tristate
flabel metal2 s 40320 59200 40432 59800 0 FreeSans 448 90 0 0 Q[9]
port 28 nsew signal tristate
flabel metal3 s 59200 12096 59800 12208 0 FreeSans 448 0 0 0 REQ_SAMPLE
port 29 nsew signal input
flabel metal2 s 5376 200 5488 800 0 FreeSans 448 90 0 0 RST
port 30 nsew signal input
flabel metal2 s 16800 200 16912 800 0 FreeSans 448 90 0 0 addI[0]
port 31 nsew signal tristate
flabel metal3 s 200 50400 800 50512 0 FreeSans 448 0 0 0 addI[1]
port 32 nsew signal tristate
flabel metal3 s 59200 23520 59800 23632 0 FreeSans 448 0 0 0 addI[2]
port 33 nsew signal tristate
flabel metal2 s 27552 200 27664 800 0 FreeSans 448 90 0 0 addI[3]
port 34 nsew signal tristate
flabel metal3 s 59200 57120 59800 57232 0 FreeSans 448 0 0 0 addI[4]
port 35 nsew signal tristate
flabel metal2 s 57120 59200 57232 59800 0 FreeSans 448 90 0 0 addI[5]
port 36 nsew signal tristate
flabel metal2 s 18144 59200 18256 59800 0 FreeSans 448 90 0 0 addQ[0]
port 37 nsew signal tristate
flabel metal2 s 23520 59200 23632 59800 0 FreeSans 448 90 0 0 addQ[1]
port 38 nsew signal tristate
flabel metal2 s 38976 200 39088 800 0 FreeSans 448 90 0 0 addQ[2]
port 39 nsew signal tristate
flabel metal3 s 200 27552 800 27664 0 FreeSans 448 0 0 0 addQ[3]
port 40 nsew signal tristate
flabel metal3 s 200 55776 800 55888 0 FreeSans 448 0 0 0 addQ[4]
port 41 nsew signal tristate
flabel metal3 s 59200 28896 59800 29008 0 FreeSans 448 0 0 0 addQ[5]
port 42 nsew signal tristate
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 43 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 44 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 44 nsew ground bidirectional
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal3 28224 56280 28224 56280 0 ACK
rlabel metal2 1400 58674 1400 58674 0 Bit_In
rlabel metal2 44408 2058 44408 2058 0 EN
rlabel metal2 55384 7056 55384 7056 0 I[0]
rlabel metal3 1358 44408 1358 44408 0 I[10]
rlabel metal3 57274 1400 57274 1400 0 I[11]
rlabel metal2 55832 2478 55832 2478 0 I[12]
rlabel metal2 55384 40824 55384 40824 0 I[1]
rlabel metal2 22568 3388 22568 3388 0 I[2]
rlabel metal3 34104 3640 34104 3640 0 I[3]
rlabel metal2 47320 56056 47320 56056 0 I[4]
rlabel metal3 1358 22232 1358 22232 0 I[5]
rlabel metal2 55384 46480 55384 46480 0 I[6]
rlabel metal3 1358 33656 1358 33656 0 I[7]
rlabel metal2 10808 2086 10808 2086 0 I[8]
rlabel metal3 1358 39032 1358 39032 0 I[9]
rlabel metal3 1358 16856 1358 16856 0 Q[0]
rlabel metal2 35112 56168 35112 56168 0 Q[10]
rlabel metal3 52640 55944 52640 55944 0 Q[11]
rlabel metal2 55944 17976 55944 17976 0 Q[12]
rlabel metal3 57666 51800 57666 51800 0 Q[1]
rlabel metal2 12152 57610 12152 57610 0 Q[2]
rlabel metal2 56 1302 56 1302 0 Q[3]
rlabel metal3 1358 10808 1358 10808 0 Q[4]
rlabel metal2 56056 35280 56056 35280 0 Q[5]
rlabel metal2 7672 56280 7672 56280 0 Q[6]
rlabel metal3 1358 5432 1358 5432 0 Q[7]
rlabel metal3 50904 3640 50904 3640 0 Q[8]
rlabel metal2 41160 56392 41160 56392 0 Q[9]
rlabel metal2 56168 10472 56168 10472 0 REQ_SAMPLE
rlabel metal2 5096 2800 5096 2800 0 RST
rlabel metal2 22904 24416 22904 24416 0 _0000_
rlabel metal3 30688 32648 30688 32648 0 _0002_
rlabel metal3 22568 23688 22568 23688 0 _0004_
rlabel metal3 30128 33096 30128 33096 0 _0005_
rlabel metal2 34216 32144 34216 32144 0 _0006_
rlabel metal2 33936 33320 33936 33320 0 _0007_
rlabel metal3 18312 22232 18312 22232 0 _0008_
rlabel metal2 37968 33320 37968 33320 0 _0009_
rlabel metal2 37744 29624 37744 29624 0 _0010_
rlabel metal3 29232 26264 29232 26264 0 _0011_
rlabel metal2 40488 34776 40488 34776 0 _0012_
rlabel metal2 40488 31304 40488 31304 0 _0013_
rlabel metal2 15400 29064 15400 29064 0 _0014_
rlabel metal2 19376 29400 19376 29400 0 _0015_
rlabel metal2 14392 25816 14392 25816 0 _0016_
rlabel metal3 12432 27384 12432 27384 0 _0017_
rlabel metal2 18872 31248 18872 31248 0 _0018_
rlabel metal2 23688 30184 23688 30184 0 _0019_
rlabel metal2 39200 4088 39200 4088 0 _0020_
rlabel metal2 39480 4368 39480 4368 0 _0021_
rlabel metal3 43064 23912 43064 23912 0 _0022_
rlabel metal2 42616 27160 42616 27160 0 _0023_
rlabel metal2 43624 22512 43624 22512 0 _0024_
rlabel metal2 46760 21616 46760 21616 0 _0025_
rlabel metal2 42728 24248 42728 24248 0 _0026_
rlabel metal4 42056 15848 42056 15848 0 _0027_
rlabel metal2 45416 12264 45416 12264 0 _0028_
rlabel metal2 44072 11872 44072 11872 0 _0029_
rlabel metal2 31416 11984 31416 11984 0 _0030_
rlabel metal2 31640 8456 31640 8456 0 _0031_
rlabel metal3 29568 19992 29568 19992 0 _0032_
rlabel metal2 30520 6104 30520 6104 0 _0033_
rlabel metal3 46480 10808 46480 10808 0 _0034_
rlabel metal3 51296 16744 51296 16744 0 _0035_
rlabel metal2 49560 22848 49560 22848 0 _0036_
rlabel metal2 48720 23912 48720 23912 0 _0037_
rlabel metal2 48888 25872 48888 25872 0 _0038_
rlabel metal2 50232 20720 50232 20720 0 _0039_
rlabel metal2 40208 27048 40208 27048 0 _0040_
rlabel metal3 41944 14896 41944 14896 0 _0041_
rlabel metal2 49896 17528 49896 17528 0 _0042_
rlabel metal2 51800 5712 51800 5712 0 _0043_
rlabel metal2 49728 16744 49728 16744 0 _0044_
rlabel metal2 45976 7168 45976 7168 0 _0045_
rlabel metal3 36904 5768 36904 5768 0 _0046_
rlabel metal2 50344 10584 50344 10584 0 _0047_
rlabel metal2 55944 23016 55944 23016 0 _0048_
rlabel metal2 44744 20944 44744 20944 0 _0049_
rlabel metal3 47040 27608 47040 27608 0 _0050_
rlabel metal2 52136 20328 52136 20328 0 _0051_
rlabel metal3 46704 2520 46704 2520 0 _0052_
rlabel metal2 51688 19096 51688 19096 0 _0053_
rlabel metal3 56112 25480 56112 25480 0 _0054_
rlabel metal2 51016 5600 51016 5600 0 _0055_
rlabel metal2 42504 26152 42504 26152 0 _0056_
rlabel metal3 41888 26936 41888 26936 0 _0057_
rlabel metal2 50008 12488 50008 12488 0 _0058_
rlabel metal2 51240 10136 51240 10136 0 _0059_
rlabel metal2 49448 6832 49448 6832 0 _0060_
rlabel metal3 34776 5768 34776 5768 0 _0061_
rlabel metal2 34216 8176 34216 8176 0 _0062_
rlabel metal2 32200 7056 32200 7056 0 _0063_
rlabel metal3 33152 5992 33152 5992 0 _0064_
rlabel metal3 56448 24472 56448 24472 0 _0065_
rlabel metal2 32536 5600 32536 5600 0 _0066_
rlabel metal3 29288 4312 29288 4312 0 _0067_
rlabel metal2 32424 5880 32424 5880 0 _0068_
rlabel metal3 32368 6664 32368 6664 0 _0069_
rlabel metal2 32984 5768 32984 5768 0 _0070_
rlabel metal2 29400 4424 29400 4424 0 _0071_
rlabel metal2 31304 6104 31304 6104 0 _0072_
rlabel metal2 28392 5152 28392 5152 0 _0073_
rlabel metal2 46872 11200 46872 11200 0 _0074_
rlabel metal2 32088 10640 32088 10640 0 _0075_
rlabel metal3 40040 13832 40040 13832 0 _0076_
rlabel metal2 33208 12880 33208 12880 0 _0077_
rlabel metal2 40320 21784 40320 21784 0 _0078_
rlabel metal2 42000 20104 42000 20104 0 _0079_
rlabel metal2 40376 21000 40376 21000 0 _0080_
rlabel metal2 40768 18424 40768 18424 0 _0081_
rlabel metal2 39592 27944 39592 27944 0 _0082_
rlabel metal2 38752 13720 38752 13720 0 _0083_
rlabel metal3 36008 12936 36008 12936 0 _0084_
rlabel metal3 33992 15848 33992 15848 0 _0085_
rlabel metal2 32536 11704 32536 11704 0 _0086_
rlabel metal2 34216 11704 34216 11704 0 _0087_
rlabel metal2 26152 11760 26152 11760 0 _0088_
rlabel metal3 41160 29512 41160 29512 0 _0089_
rlabel metal2 41328 23912 41328 23912 0 _0090_
rlabel metal2 34216 16464 34216 16464 0 _0091_
rlabel metal2 41776 18648 41776 18648 0 _0092_
rlabel metal2 42840 12544 42840 12544 0 _0093_
rlabel metal2 42840 23016 42840 23016 0 _0094_
rlabel metal2 42616 11928 42616 11928 0 _0095_
rlabel metal2 57176 18760 57176 18760 0 _0096_
rlabel metal2 31080 12096 31080 12096 0 _0097_
rlabel metal3 32088 12824 32088 12824 0 _0098_
rlabel metal3 32200 12152 32200 12152 0 _0099_
rlabel metal2 26376 12320 26376 12320 0 _0100_
rlabel metal3 25536 12936 25536 12936 0 _0101_
rlabel metal2 24528 13944 24528 13944 0 _0102_
rlabel metal2 26488 11704 26488 11704 0 _0103_
rlabel metal2 26544 8232 26544 8232 0 _0104_
rlabel metal2 27048 7896 27048 7896 0 _0105_
rlabel metal2 43848 9464 43848 9464 0 _0106_
rlabel metal3 56056 15960 56056 15960 0 _0107_
rlabel metal2 40880 8232 40880 8232 0 _0108_
rlabel metal2 45752 24584 45752 24584 0 _0109_
rlabel metal2 46088 31472 46088 31472 0 _0110_
rlabel metal2 45416 30912 45416 30912 0 _0111_
rlabel metal2 45808 31192 45808 31192 0 _0112_
rlabel metal2 46368 29624 46368 29624 0 _0113_
rlabel metal3 47600 23800 47600 23800 0 _0114_
rlabel metal2 46424 22960 46424 22960 0 _0115_
rlabel metal2 45640 24080 45640 24080 0 _0116_
rlabel metal2 40488 24920 40488 24920 0 _0117_
rlabel metal2 56840 16856 56840 16856 0 _0118_
rlabel metal2 46872 25144 46872 25144 0 _0119_
rlabel metal2 45528 24976 45528 24976 0 _0120_
rlabel metal3 45696 24584 45696 24584 0 _0121_
rlabel metal3 42168 9800 42168 9800 0 _0122_
rlabel metal2 42952 7672 42952 7672 0 _0123_
rlabel metal2 43624 8736 43624 8736 0 _0124_
rlabel metal2 26712 9464 26712 9464 0 _0125_
rlabel metal3 44632 19992 44632 19992 0 _0126_
rlabel metal2 45864 18032 45864 18032 0 _0127_
rlabel metal2 46648 17920 46648 17920 0 _0128_
rlabel metal2 57848 21616 57848 21616 0 _0129_
rlabel metal3 48608 19992 48608 19992 0 _0130_
rlabel metal3 45360 21560 45360 21560 0 _0131_
rlabel metal3 45696 21672 45696 21672 0 _0132_
rlabel metal2 46368 21560 46368 21560 0 _0133_
rlabel metal2 46312 31808 46312 31808 0 _0134_
rlabel metal2 46872 20552 46872 20552 0 _0135_
rlabel metal3 47432 19992 47432 19992 0 _0136_
rlabel metal3 23744 20552 23744 20552 0 _0137_
rlabel metal3 38808 3080 38808 3080 0 _0138_
rlabel metal2 24136 18760 24136 18760 0 _0139_
rlabel metal2 57568 25704 57568 25704 0 _0140_
rlabel metal2 25032 12264 25032 12264 0 _0141_
rlabel metal2 26320 7448 26320 7448 0 _0142_
rlabel metal2 28392 6608 28392 6608 0 _0143_
rlabel metal2 28896 4200 28896 4200 0 _0144_
rlabel metal2 30296 3976 30296 3976 0 _0145_
rlabel metal3 34776 16856 34776 16856 0 _0146_
rlabel metal2 40544 27832 40544 27832 0 _0147_
rlabel metal3 44352 12936 44352 12936 0 _0148_
rlabel metal2 46648 11816 46648 11816 0 _0149_
rlabel metal3 50120 22120 50120 22120 0 _0150_
rlabel metal2 47712 20552 47712 20552 0 _0151_
rlabel metal2 35784 15148 35784 15148 0 _0152_
rlabel metal3 43120 20776 43120 20776 0 _0153_
rlabel metal2 44184 20272 44184 20272 0 _0154_
rlabel metal3 43176 20552 43176 20552 0 _0155_
rlabel metal2 35336 14560 35336 14560 0 _0156_
rlabel metal2 29736 13608 29736 13608 0 _0157_
rlabel metal2 31416 14280 31416 14280 0 _0158_
rlabel metal3 27608 14392 27608 14392 0 _0159_
rlabel metal2 26264 9968 26264 9968 0 _0160_
rlabel metal3 40936 2856 40936 2856 0 _0161_
rlabel metal3 23464 14504 23464 14504 0 _0162_
rlabel metal3 40096 8232 40096 8232 0 _0163_
rlabel metal2 39256 18368 39256 18368 0 _0164_
rlabel metal2 38920 18984 38920 18984 0 _0165_
rlabel metal4 39480 15624 39480 15624 0 _0166_
rlabel metal2 40040 11648 40040 11648 0 _0167_
rlabel metal3 40600 17864 40600 17864 0 _0168_
rlabel metal2 40152 21000 40152 21000 0 _0169_
rlabel metal2 45416 14672 45416 14672 0 _0170_
rlabel metal3 41272 14504 41272 14504 0 _0171_
rlabel metal2 26544 17080 26544 17080 0 _0172_
rlabel metal3 47656 17080 47656 17080 0 _0173_
rlabel metal2 41832 15344 41832 15344 0 _0174_
rlabel metal2 40264 10808 40264 10808 0 _0175_
rlabel metal2 39256 9800 39256 9800 0 _0176_
rlabel metal3 39480 8344 39480 8344 0 _0177_
rlabel metal2 23464 12656 23464 12656 0 _0178_
rlabel metal2 23520 21784 23520 21784 0 _0179_
rlabel metal3 22736 21560 22736 21560 0 _0180_
rlabel metal2 31416 21896 31416 21896 0 _0181_
rlabel metal3 41552 23128 41552 23128 0 _0182_
rlabel metal2 27216 22344 27216 22344 0 _0183_
rlabel metal3 40600 22232 40600 22232 0 _0184_
rlabel metal2 39928 24416 39928 24416 0 _0185_
rlabel metal3 40320 22456 40320 22456 0 _0186_
rlabel metal2 40488 22512 40488 22512 0 _0187_
rlabel metal3 43848 25144 43848 25144 0 _0188_
rlabel metal2 30352 23352 30352 23352 0 _0189_
rlabel metal3 24080 21672 24080 21672 0 _0190_
rlabel metal3 22680 13944 22680 13944 0 _0191_
rlabel metal2 22568 14224 22568 14224 0 _0192_
rlabel metal3 21504 17640 21504 17640 0 _0193_
rlabel metal3 48496 29400 48496 29400 0 _0194_
rlabel metal2 26376 10696 26376 10696 0 _0195_
rlabel metal3 26040 13384 26040 13384 0 _0196_
rlabel metal2 21672 17192 21672 17192 0 _0197_
rlabel metal2 28504 4984 28504 4984 0 _0198_
rlabel metal2 25536 7672 25536 7672 0 _0199_
rlabel metal2 22064 18424 22064 18424 0 _0200_
rlabel metal3 20944 14616 20944 14616 0 _0201_
rlabel metal3 21616 16856 21616 16856 0 _0202_
rlabel metal2 25648 14280 25648 14280 0 _0203_
rlabel metal2 47208 21056 47208 21056 0 _0204_
rlabel metal2 39088 27720 39088 27720 0 _0205_
rlabel metal2 40880 16968 40880 16968 0 _0206_
rlabel metal3 40320 18984 40320 18984 0 _0207_
rlabel metal2 39704 16520 39704 16520 0 _0208_
rlabel metal3 34104 17080 34104 17080 0 _0209_
rlabel metal2 39368 15568 39368 15568 0 _0210_
rlabel metal2 39592 15344 39592 15344 0 _0211_
rlabel metal2 38920 15904 38920 15904 0 _0212_
rlabel metal2 38808 14616 38808 14616 0 _0213_
rlabel metal3 28448 14504 28448 14504 0 _0214_
rlabel metal2 50232 29792 50232 29792 0 _0215_
rlabel metal3 26320 14504 26320 14504 0 _0216_
rlabel metal3 23128 15064 23128 15064 0 _0217_
rlabel metal3 37128 7560 37128 7560 0 _0218_
rlabel metal2 35224 22512 35224 22512 0 _0219_
rlabel metal2 31808 24696 31808 24696 0 _0220_
rlabel metal2 31696 19432 31696 19432 0 _0221_
rlabel metal2 32648 17304 32648 17304 0 _0222_
rlabel metal2 36792 16576 36792 16576 0 _0223_
rlabel metal2 42392 19040 42392 19040 0 _0224_
rlabel metal2 42728 17976 42728 17976 0 _0225_
rlabel metal2 53816 26152 53816 26152 0 _0226_
rlabel metal2 42168 18088 42168 18088 0 _0227_
rlabel metal2 41272 17528 41272 17528 0 _0228_
rlabel metal2 39928 17024 39928 17024 0 _0229_
rlabel metal2 39144 10640 39144 10640 0 _0230_
rlabel metal2 36568 8848 36568 8848 0 _0231_
rlabel metal2 35224 9184 35224 9184 0 _0232_
rlabel metal2 38416 9240 38416 9240 0 _0233_
rlabel metal2 37856 9912 37856 9912 0 _0234_
rlabel metal2 20216 13720 20216 13720 0 _0235_
rlabel metal3 23016 21448 23016 21448 0 _0236_
rlabel metal2 54040 22456 54040 22456 0 _0237_
rlabel metal2 36904 22680 36904 22680 0 _0238_
rlabel metal2 37016 20384 37016 20384 0 _0239_
rlabel metal2 44352 19432 44352 19432 0 _0240_
rlabel metal2 36120 20272 36120 20272 0 _0241_
rlabel metal2 35784 18592 35784 18592 0 _0242_
rlabel metal2 22232 20384 22232 20384 0 _0243_
rlabel metal2 19152 13720 19152 13720 0 _0244_
rlabel metal2 18424 16520 18424 16520 0 _0245_
rlabel metal2 20888 18480 20888 18480 0 _0246_
rlabel metal2 18984 18704 18984 18704 0 _0247_
rlabel metal2 53984 15288 53984 15288 0 _0248_
rlabel metal2 2744 20608 2744 20608 0 _0249_
rlabel metal2 32872 26096 32872 26096 0 _0250_
rlabel metal2 31528 26040 31528 26040 0 _0251_
rlabel metal2 36456 25480 36456 25480 0 _0252_
rlabel metal2 40936 24640 40936 24640 0 _0253_
rlabel metal2 38920 27160 38920 27160 0 _0254_
rlabel metal2 37464 25704 37464 25704 0 _0255_
rlabel metal3 36120 25368 36120 25368 0 _0256_
rlabel metal2 34160 24920 34160 24920 0 _0257_
rlabel metal2 43848 25872 43848 25872 0 _0258_
rlabel metal2 44072 24360 44072 24360 0 _0259_
rlabel metal2 32760 24808 32760 24808 0 _0260_
rlabel metal2 30072 17920 30072 17920 0 _0261_
rlabel metal3 29120 13048 29120 13048 0 _0262_
rlabel metal3 28840 9800 28840 9800 0 _0263_
rlabel metal2 27832 14168 27832 14168 0 _0264_
rlabel metal2 26152 14112 26152 14112 0 _0265_
rlabel metal3 34440 27608 34440 27608 0 _0266_
rlabel metal2 38920 26656 38920 26656 0 _0267_
rlabel metal2 37688 26992 37688 26992 0 _0268_
rlabel metal2 35560 21560 35560 21560 0 _0269_
rlabel metal3 36232 28392 36232 28392 0 _0270_
rlabel metal3 35504 25704 35504 25704 0 _0271_
rlabel metal2 34104 21504 34104 21504 0 _0272_
rlabel metal3 34888 24472 34888 24472 0 _0273_
rlabel metal2 35168 23912 35168 23912 0 _0274_
rlabel metal2 36568 24416 36568 24416 0 _0275_
rlabel metal2 35448 23688 35448 23688 0 _0276_
rlabel metal3 34888 23912 34888 23912 0 _0277_
rlabel metal2 40320 9688 40320 9688 0 _0278_
rlabel metal2 39928 9576 39928 9576 0 _0279_
rlabel metal2 27440 23240 27440 23240 0 _0280_
rlabel metal3 35448 11256 35448 11256 0 _0281_
rlabel metal3 35112 9688 35112 9688 0 _0282_
rlabel metal2 35504 11928 35504 11928 0 _0283_
rlabel metal2 35280 12376 35280 12376 0 _0284_
rlabel metal2 17976 14000 17976 14000 0 _0285_
rlabel metal2 28504 23800 28504 23800 0 _0286_
rlabel metal2 28504 21224 28504 21224 0 _0287_
rlabel metal2 25984 19432 25984 19432 0 _0288_
rlabel metal2 24640 15960 24640 15960 0 _0289_
rlabel metal3 36456 16856 36456 16856 0 _0290_
rlabel metal3 20272 26152 20272 26152 0 _0291_
rlabel metal2 38864 24136 38864 24136 0 _0292_
rlabel metal2 36120 17080 36120 17080 0 _0293_
rlabel metal2 35504 18536 35504 18536 0 _0294_
rlabel metal2 40488 17304 40488 17304 0 _0295_
rlabel metal3 37184 17080 37184 17080 0 _0296_
rlabel metal2 24920 16128 24920 16128 0 _0297_
rlabel metal3 15568 14728 15568 14728 0 _0298_
rlabel metal3 16632 16072 16632 16072 0 _0299_
rlabel metal2 18760 14112 18760 14112 0 _0300_
rlabel metal2 19488 14504 19488 14504 0 _0301_
rlabel metal2 16408 15904 16408 15904 0 _0302_
rlabel metal2 16576 17864 16576 17864 0 _0303_
rlabel metal3 18088 17416 18088 17416 0 _0304_
rlabel metal2 17864 17304 17864 17304 0 _0305_
rlabel metal3 17136 17864 17136 17864 0 _0306_
rlabel metal2 56672 45640 56672 45640 0 _0307_
rlabel metal3 15008 13720 15008 13720 0 _0308_
rlabel metal2 14952 14000 14952 14000 0 _0309_
rlabel metal3 14840 13160 14840 13160 0 _0310_
rlabel metal2 8792 30856 8792 30856 0 _0311_
rlabel metal3 30240 10696 30240 10696 0 _0312_
rlabel metal2 29400 10528 29400 10528 0 _0313_
rlabel metal4 27944 15400 27944 15400 0 _0314_
rlabel metal2 39816 24304 39816 24304 0 _0315_
rlabel metal3 38920 21728 38920 21728 0 _0316_
rlabel metal3 38360 22120 38360 22120 0 _0317_
rlabel metal2 39032 26320 39032 26320 0 _0318_
rlabel metal2 37352 21952 37352 21952 0 _0319_
rlabel metal3 35616 22456 35616 22456 0 _0320_
rlabel metal2 33936 23352 33936 23352 0 _0321_
rlabel metal2 8008 33488 8008 33488 0 _0322_
rlabel metal3 32144 25368 32144 25368 0 _0323_
rlabel metal2 32760 24080 32760 24080 0 _0324_
rlabel metal3 31136 15512 31136 15512 0 _0325_
rlabel metal2 29176 14336 29176 14336 0 _0326_
rlabel metal2 28952 12040 28952 12040 0 _0327_
rlabel metal2 24136 10976 24136 10976 0 _0328_
rlabel metal3 36792 18984 36792 18984 0 _0329_
rlabel metal2 35336 19320 35336 19320 0 _0330_
rlabel metal2 34496 19208 34496 19208 0 _0331_
rlabel metal2 34888 20552 34888 20552 0 _0332_
rlabel metal2 3080 52808 3080 52808 0 _0333_
rlabel metal2 34832 19880 34832 19880 0 _0334_
rlabel metal2 25368 9800 25368 9800 0 _0335_
rlabel metal3 35224 9912 35224 9912 0 _0336_
rlabel metal2 24920 9520 24920 9520 0 _0337_
rlabel metal2 23128 10640 23128 10640 0 _0338_
rlabel metal3 31472 21672 31472 21672 0 _0339_
rlabel metal2 34664 23072 34664 23072 0 _0340_
rlabel metal2 31696 21560 31696 21560 0 _0341_
rlabel metal2 31416 16688 31416 16688 0 _0342_
rlabel metal3 30632 15232 30632 15232 0 _0343_
rlabel metal2 10248 32088 10248 32088 0 _0344_
rlabel metal2 23240 11648 23240 11648 0 _0345_
rlabel metal2 22904 11816 22904 11816 0 _0346_
rlabel metal2 15512 12656 15512 12656 0 _0347_
rlabel metal2 15512 13440 15512 13440 0 _0348_
rlabel metal2 16520 13160 16520 13160 0 _0349_
rlabel metal3 15960 13944 15960 13944 0 _0350_
rlabel metal3 15960 15848 15960 15848 0 _0351_
rlabel metal2 16072 16912 16072 16912 0 _0352_
rlabel metal3 15736 17752 15736 17752 0 _0353_
rlabel metal2 2744 30016 2744 30016 0 _0354_
rlabel metal3 5488 34888 5488 34888 0 _0355_
rlabel metal3 27496 9128 27496 9128 0 _0356_
rlabel metal2 38304 20776 38304 20776 0 _0357_
rlabel metal2 38920 23016 38920 23016 0 _0358_
rlabel metal2 38024 20384 38024 20384 0 _0359_
rlabel metal2 29848 19152 29848 19152 0 _0360_
rlabel metal3 27104 18536 27104 18536 0 _0361_
rlabel metal2 26992 17640 26992 17640 0 _0362_
rlabel metal2 20552 11704 20552 11704 0 _0363_
rlabel metal3 36456 27048 36456 27048 0 _0364_
rlabel metal3 9520 32536 9520 32536 0 _0365_
rlabel metal2 30744 19096 30744 19096 0 _0366_
rlabel metal2 27272 19992 27272 19992 0 _0367_
rlabel metal2 21560 13104 21560 13104 0 _0368_
rlabel metal2 35224 17304 35224 17304 0 _0369_
rlabel metal2 35784 17640 35784 17640 0 _0370_
rlabel metal2 35728 15624 35728 15624 0 _0371_
rlabel metal3 36736 12152 36736 12152 0 _0372_
rlabel metal3 36792 12264 36792 12264 0 _0373_
rlabel metal2 21224 12376 21224 12376 0 _0374_
rlabel metal2 18984 12432 18984 12432 0 _0375_
rlabel metal2 5656 32256 5656 32256 0 _0376_
rlabel metal2 18312 11816 18312 11816 0 _0377_
rlabel metal3 16576 10696 16576 10696 0 _0378_
rlabel metal2 24360 10864 24360 10864 0 _0379_
rlabel metal3 22092 10696 22092 10696 0 _0380_
rlabel metal2 15624 10248 15624 10248 0 _0381_
rlabel metal2 16408 13440 16408 13440 0 _0382_
rlabel metal2 15904 10696 15904 10696 0 _0383_
rlabel metal2 16184 10528 16184 10528 0 _0384_
rlabel metal2 14616 10136 14616 10136 0 _0385_
rlabel metal3 13440 9128 13440 9128 0 _0386_
rlabel metal2 20888 32704 20888 32704 0 _0387_
rlabel metal2 19880 11480 19880 11480 0 _0388_
rlabel metal2 19264 10696 19264 10696 0 _0389_
rlabel metal2 28616 18032 28616 18032 0 _0390_
rlabel metal3 33712 22232 33712 22232 0 _0391_
rlabel metal2 33880 19880 33880 19880 0 _0392_
rlabel metal3 31248 17416 31248 17416 0 _0393_
rlabel metal3 30072 17528 30072 17528 0 _0394_
rlabel metal3 29008 17528 29008 17528 0 _0395_
rlabel metal2 28000 15176 28000 15176 0 _0396_
rlabel metal2 22624 37912 22624 37912 0 _0397_
rlabel metal2 28728 15960 28728 15960 0 _0398_
rlabel metal2 28336 11368 28336 11368 0 _0399_
rlabel metal2 21728 6776 21728 6776 0 _0400_
rlabel metal2 33320 18144 33320 18144 0 _0401_
rlabel metal2 33656 15960 33656 15960 0 _0402_
rlabel metal2 35000 9240 35000 9240 0 _0403_
rlabel metal3 35112 8344 35112 8344 0 _0404_
rlabel metal2 22400 8120 22400 8120 0 _0405_
rlabel via2 25928 18088 25928 18088 0 _0406_
rlabel metal2 24584 17920 24584 17920 0 _0407_
rlabel metal3 4032 34328 4032 34328 0 _0408_
rlabel metal3 22400 8344 22400 8344 0 _0409_
rlabel metal2 19656 10528 19656 10528 0 _0410_
rlabel metal2 18312 10528 18312 10528 0 _0411_
rlabel metal2 18648 7896 18648 7896 0 _0412_
rlabel metal3 16240 10024 16240 10024 0 _0413_
rlabel metal2 16576 10808 16576 10808 0 _0414_
rlabel metal2 18312 7952 18312 7952 0 _0415_
rlabel metal3 15456 11368 15456 11368 0 _0416_
rlabel metal2 2520 12096 2520 12096 0 _0417_
rlabel metal2 3192 40152 3192 40152 0 _0418_
rlabel metal3 33992 10472 33992 10472 0 _0419_
rlabel metal2 25704 9408 25704 9408 0 _0420_
rlabel metal2 33320 8400 33320 8400 0 _0421_
rlabel metal2 25648 8232 25648 8232 0 _0422_
rlabel metal2 25816 17304 25816 17304 0 _0423_
rlabel metal3 26040 8232 26040 8232 0 _0424_
rlabel metal3 25256 7336 25256 7336 0 _0425_
rlabel metal2 23744 8120 23744 8120 0 _0426_
rlabel metal3 24472 8344 24472 8344 0 _0427_
rlabel metal3 22792 7448 22792 7448 0 _0428_
rlabel metal2 13608 32144 13608 32144 0 _0429_
rlabel metal2 30072 7896 30072 7896 0 _0430_
rlabel metal2 32032 17080 32032 17080 0 _0431_
rlabel metal2 32256 16296 32256 16296 0 _0432_
rlabel metal2 29512 7560 29512 7560 0 _0433_
rlabel metal2 22344 7224 22344 7224 0 _0434_
rlabel metal3 21056 6104 21056 6104 0 _0435_
rlabel metal3 21224 7448 21224 7448 0 _0436_
rlabel metal2 20216 7840 20216 7840 0 _0437_
rlabel metal2 20440 6832 20440 6832 0 _0438_
rlabel metal3 18872 8232 18872 8232 0 _0439_
rlabel metal4 22680 44632 22680 44632 0 _0440_
rlabel metal2 18032 8120 18032 8120 0 _0441_
rlabel metal2 17528 7336 17528 7336 0 _0442_
rlabel metal3 3024 9688 3024 9688 0 _0443_
rlabel metal2 23240 6944 23240 6944 0 _0444_
rlabel metal2 22064 5880 22064 5880 0 _0445_
rlabel metal2 27608 17360 27608 17360 0 _0446_
rlabel metal2 27272 17360 27272 17360 0 _0447_
rlabel metal2 26712 15400 26712 15400 0 _0448_
rlabel metal2 26656 9128 26656 9128 0 _0449_
rlabel metal2 21896 35448 21896 35448 0 _0450_
rlabel metal2 23912 7784 23912 7784 0 _0451_
rlabel via2 22456 4984 22456 4984 0 _0452_
rlabel metal2 20776 5320 20776 5320 0 _0453_
rlabel metal3 21224 5096 21224 5096 0 _0454_
rlabel metal2 20664 4704 20664 4704 0 _0455_
rlabel metal2 23912 3472 23912 3472 0 _0456_
rlabel metal2 22120 5488 22120 5488 0 _0457_
rlabel metal2 25144 4928 25144 4928 0 _0458_
rlabel metal2 24584 6160 24584 6160 0 _0459_
rlabel metal2 1904 32760 1904 32760 0 _0460_
rlabel metal2 24248 5992 24248 5992 0 _0461_
rlabel metal3 24752 4984 24752 4984 0 _0462_
rlabel metal2 24920 5376 24920 5376 0 _0463_
rlabel metal3 52920 8344 52920 8344 0 _0464_
rlabel metal3 57064 39592 57064 39592 0 _0465_
rlabel metal2 33880 31864 33880 31864 0 _0466_
rlabel metal2 24024 29232 24024 29232 0 _0467_
rlabel metal3 3024 31192 3024 31192 0 _0468_
rlabel metal2 15624 25536 15624 25536 0 _0469_
rlabel metal2 17976 23408 17976 23408 0 _0470_
rlabel metal2 18928 22344 18928 22344 0 _0471_
rlabel metal2 19992 29176 19992 29176 0 _0472_
rlabel metal2 35672 30072 35672 30072 0 _0473_
rlabel metal2 35448 29288 35448 29288 0 _0474_
rlabel metal2 36960 29400 36960 29400 0 _0475_
rlabel metal2 19096 36008 19096 36008 0 _0476_
rlabel metal2 30632 29008 30632 29008 0 _0477_
rlabel metal3 29232 27944 29232 27944 0 _0478_
rlabel metal2 28224 25704 28224 25704 0 _0479_
rlabel metal2 32088 29008 32088 29008 0 _0480_
rlabel metal3 33656 28504 33656 28504 0 _0481_
rlabel metal2 31976 30240 31976 30240 0 _0482_
rlabel metal2 32536 29736 32536 29736 0 _0483_
rlabel metal2 21896 47544 21896 47544 0 _0484_
rlabel metal3 15232 29400 15232 29400 0 _0485_
rlabel metal2 19768 30240 19768 30240 0 _0486_
rlabel metal2 14952 29736 14952 29736 0 _0487_
rlabel metal2 15176 30632 15176 30632 0 _0488_
rlabel metal2 14616 26180 14616 26180 0 _0489_
rlabel metal2 10976 27048 10976 27048 0 _0490_
rlabel metal2 23856 33320 23856 33320 0 _0491_
rlabel metal2 22456 31808 22456 31808 0 _0492_
rlabel metal2 22680 32872 22680 32872 0 _0493_
rlabel metal2 19600 31976 19600 31976 0 _0494_
rlabel metal2 23072 33096 23072 33096 0 _0495_
rlabel metal2 23352 32200 23352 32200 0 _0496_
rlabel metal2 37576 4648 37576 4648 0 _0497_
rlabel metal2 24024 34944 24024 34944 0 _0498_
rlabel metal2 22792 34608 22792 34608 0 _0499_
rlabel metal2 2744 32088 2744 32088 0 _0500_
rlabel metal2 11592 34160 11592 34160 0 _0501_
rlabel metal4 24696 47712 24696 47712 0 _0502_
rlabel metal2 27160 52360 27160 52360 0 _0503_
rlabel metal3 25872 45640 25872 45640 0 _0504_
rlabel metal2 24248 34160 24248 34160 0 _0505_
rlabel metal3 33208 35784 33208 35784 0 _0506_
rlabel metal2 25592 49336 25592 49336 0 _0507_
rlabel metal2 26152 23296 26152 23296 0 _0508_
rlabel metal2 24248 19208 24248 19208 0 _0509_
rlabel metal3 25424 28056 25424 28056 0 _0510_
rlabel metal2 44520 8120 44520 8120 0 _0511_
rlabel metal3 29792 15288 29792 15288 0 _0512_
rlabel metal2 23240 24080 23240 24080 0 _0513_
rlabel metal2 26488 25088 26488 25088 0 _0514_
rlabel metal3 25312 20664 25312 20664 0 _0515_
rlabel metal2 24360 21392 24360 21392 0 _0516_
rlabel metal2 26432 24696 26432 24696 0 _0517_
rlabel metal2 24920 23912 24920 23912 0 _0518_
rlabel metal2 24584 23072 24584 23072 0 _0519_
rlabel metal2 31528 41160 31528 41160 0 _0520_
rlabel metal2 32088 52136 32088 52136 0 _0521_
rlabel metal2 30408 48160 30408 48160 0 _0522_
rlabel metal3 30016 49000 30016 49000 0 _0523_
rlabel metal2 31808 33544 31808 33544 0 _0524_
rlabel metal2 29792 33320 29792 33320 0 _0525_
rlabel metal2 30240 33320 30240 33320 0 _0526_
rlabel metal3 18592 27832 18592 27832 0 _0527_
rlabel metal3 18704 26264 18704 26264 0 _0528_
rlabel metal2 26376 26712 26376 26712 0 _0529_
rlabel metal2 28000 50456 28000 50456 0 _0530_
rlabel metal3 37240 48104 37240 48104 0 _0531_
rlabel metal2 31640 52192 31640 52192 0 _0532_
rlabel metal2 20664 35728 20664 35728 0 _0533_
rlabel metal2 13720 43680 13720 43680 0 _0534_
rlabel metal3 7112 33208 7112 33208 0 _0535_
rlabel metal2 11928 32256 11928 32256 0 _0536_
rlabel metal2 20776 41776 20776 41776 0 _0537_
rlabel metal3 17808 39480 17808 39480 0 _0538_
rlabel metal2 22456 40152 22456 40152 0 _0539_
rlabel metal2 20216 39872 20216 39872 0 _0540_
rlabel metal2 1848 37800 1848 37800 0 _0541_
rlabel metal2 3080 30072 3080 30072 0 _0542_
rlabel metal2 17640 48776 17640 48776 0 _0543_
rlabel metal2 20328 40600 20328 40600 0 _0544_
rlabel metal2 2912 31752 2912 31752 0 _0545_
rlabel metal2 3864 35280 3864 35280 0 _0546_
rlabel metal3 4424 41048 4424 41048 0 _0547_
rlabel metal2 2072 48160 2072 48160 0 _0548_
rlabel metal2 9576 42392 9576 42392 0 _0549_
rlabel metal2 9800 42224 9800 42224 0 _0550_
rlabel metal2 6384 35672 6384 35672 0 _0551_
rlabel metal2 4648 45976 4648 45976 0 _0552_
rlabel metal3 12264 25032 12264 25032 0 _0553_
rlabel metal2 16744 33208 16744 33208 0 _0554_
rlabel metal2 18760 34384 18760 34384 0 _0555_
rlabel metal2 17640 32984 17640 32984 0 _0556_
rlabel metal2 18872 34944 18872 34944 0 _0557_
rlabel metal3 19544 40096 19544 40096 0 _0558_
rlabel metal2 14952 35280 14952 35280 0 _0559_
rlabel metal3 10640 38920 10640 38920 0 _0560_
rlabel metal3 22960 38696 22960 38696 0 _0561_
rlabel metal2 3136 35672 3136 35672 0 _0562_
rlabel metal2 2408 42840 2408 42840 0 _0563_
rlabel metal2 3080 31752 3080 31752 0 _0564_
rlabel metal3 2520 29624 2520 29624 0 _0565_
rlabel metal2 2968 34216 2968 34216 0 _0566_
rlabel metal2 2408 40432 2408 40432 0 _0567_
rlabel metal3 2688 31080 2688 31080 0 _0568_
rlabel metal3 22568 41384 22568 41384 0 _0569_
rlabel metal3 22960 41272 22960 41272 0 _0570_
rlabel metal2 8120 44016 8120 44016 0 _0571_
rlabel metal3 2128 53256 2128 53256 0 _0572_
rlabel metal2 22008 47768 22008 47768 0 _0573_
rlabel metal3 24640 49896 24640 49896 0 _0574_
rlabel metal2 24584 41720 24584 41720 0 _0575_
rlabel metal3 25200 41944 25200 41944 0 _0576_
rlabel metal2 25872 42728 25872 42728 0 _0577_
rlabel metal2 28952 40936 28952 40936 0 _0578_
rlabel metal2 16576 39368 16576 39368 0 _0579_
rlabel metal2 17976 40712 17976 40712 0 _0580_
rlabel metal2 17864 35560 17864 35560 0 _0581_
rlabel metal2 18424 41048 18424 41048 0 _0582_
rlabel metal2 6440 38808 6440 38808 0 _0583_
rlabel metal3 17024 34328 17024 34328 0 _0584_
rlabel metal2 9800 36064 9800 36064 0 _0585_
rlabel metal2 12152 41272 12152 41272 0 _0586_
rlabel metal3 7672 35336 7672 35336 0 _0587_
rlabel metal3 17528 48216 17528 48216 0 _0588_
rlabel metal2 18480 37240 18480 37240 0 _0589_
rlabel metal2 11480 34888 11480 34888 0 _0590_
rlabel metal2 2744 35280 2744 35280 0 _0591_
rlabel metal3 9688 47432 9688 47432 0 _0592_
rlabel metal3 8680 32424 8680 32424 0 _0593_
rlabel metal2 14784 48216 14784 48216 0 _0594_
rlabel metal2 18872 36568 18872 36568 0 _0595_
rlabel metal2 19320 32984 19320 32984 0 _0596_
rlabel metal2 21672 36288 21672 36288 0 _0597_
rlabel metal2 19880 47712 19880 47712 0 _0598_
rlabel metal2 40320 51576 40320 51576 0 _0599_
rlabel metal2 1960 41776 1960 41776 0 _0600_
rlabel metal2 7560 41944 7560 41944 0 _0601_
rlabel metal2 3192 43400 3192 43400 0 _0602_
rlabel metal4 8008 45192 8008 45192 0 _0603_
rlabel metal3 1792 52808 1792 52808 0 _0604_
rlabel metal2 15736 38836 15736 38836 0 _0605_
rlabel metal2 19096 37632 19096 37632 0 _0606_
rlabel metal2 40544 44968 40544 44968 0 _0607_
rlabel metal3 37184 40376 37184 40376 0 _0608_
rlabel metal2 38136 39256 38136 39256 0 _0609_
rlabel metal2 31416 36792 31416 36792 0 _0610_
rlabel metal2 29624 37016 29624 37016 0 _0611_
rlabel metal2 23464 46256 23464 46256 0 _0612_
rlabel metal2 16688 41048 16688 41048 0 _0613_
rlabel metal2 4536 36400 4536 36400 0 _0614_
rlabel metal2 2744 45584 2744 45584 0 _0615_
rlabel metal3 14784 36344 14784 36344 0 _0616_
rlabel metal2 12992 41720 12992 41720 0 _0617_
rlabel metal2 15400 43512 15400 43512 0 _0618_
rlabel metal3 14784 47656 14784 47656 0 _0619_
rlabel metal3 21280 37912 21280 37912 0 _0620_
rlabel metal2 2632 40152 2632 40152 0 _0621_
rlabel metal3 15960 36344 15960 36344 0 _0622_
rlabel metal2 21000 39144 21000 39144 0 _0623_
rlabel metal2 16520 44912 16520 44912 0 _0624_
rlabel metal2 3192 53144 3192 53144 0 _0625_
rlabel metal2 1848 45752 1848 45752 0 _0626_
rlabel metal2 24584 49224 24584 49224 0 _0627_
rlabel metal2 19768 43624 19768 43624 0 _0628_
rlabel metal2 18816 40264 18816 40264 0 _0629_
rlabel metal2 20328 38080 20328 38080 0 _0630_
rlabel metal2 15456 49000 15456 49000 0 _0631_
rlabel metal2 24136 40712 24136 40712 0 _0632_
rlabel metal2 25088 39704 25088 39704 0 _0633_
rlabel metal3 25144 38696 25144 38696 0 _0634_
rlabel metal2 26712 37520 26712 37520 0 _0635_
rlabel metal2 29568 36456 29568 36456 0 _0636_
rlabel metal3 5432 17080 5432 17080 0 _0637_
rlabel metal2 28840 36512 28840 36512 0 _0638_
rlabel metal2 39032 35952 39032 35952 0 _0639_
rlabel metal3 36512 50680 36512 50680 0 _0640_
rlabel metal2 32312 42112 32312 42112 0 _0641_
rlabel metal2 32592 37240 32592 37240 0 _0642_
rlabel metal2 22904 36960 22904 36960 0 _0643_
rlabel metal3 1904 52248 1904 52248 0 _0644_
rlabel metal2 29344 51240 29344 51240 0 _0645_
rlabel metal2 17024 34888 17024 34888 0 _0646_
rlabel metal2 23576 36344 23576 36344 0 _0647_
rlabel metal2 24024 43064 24024 43064 0 _0648_
rlabel metal2 23800 37296 23800 37296 0 _0649_
rlabel metal2 2856 30240 2856 30240 0 _0650_
rlabel metal2 2296 42000 2296 42000 0 _0651_
rlabel metal2 2744 43232 2744 43232 0 _0652_
rlabel metal2 3864 43456 3864 43456 0 _0653_
rlabel metal2 12040 44800 12040 44800 0 _0654_
rlabel metal2 6328 36792 6328 36792 0 _0655_
rlabel metal2 10920 36904 10920 36904 0 _0656_
rlabel metal2 14504 37744 14504 37744 0 _0657_
rlabel metal2 11704 39116 11704 39116 0 _0658_
rlabel metal2 29904 39368 29904 39368 0 _0659_
rlabel metal2 31976 37688 31976 37688 0 _0660_
rlabel metal3 33264 36456 33264 36456 0 _0661_
rlabel metal2 34664 36288 34664 36288 0 _0662_
rlabel metal2 3304 26880 3304 26880 0 _0663_
rlabel metal2 2240 27160 2240 27160 0 _0664_
rlabel metal2 2632 46088 2632 46088 0 _0665_
rlabel metal2 2912 47208 2912 47208 0 _0666_
rlabel metal4 14056 47096 14056 47096 0 _0667_
rlabel metal3 19992 44184 19992 44184 0 _0668_
rlabel metal2 3304 43288 3304 43288 0 _0669_
rlabel metal2 12320 43512 12320 43512 0 _0670_
rlabel metal2 2240 40376 2240 40376 0 _0671_
rlabel metal2 11032 43176 11032 43176 0 _0672_
rlabel metal2 15288 47600 15288 47600 0 _0673_
rlabel metal2 14896 47208 14896 47208 0 _0674_
rlabel metal2 22568 43456 22568 43456 0 _0675_
rlabel metal2 18872 45360 18872 45360 0 _0676_
rlabel metal2 18984 44688 18984 44688 0 _0677_
rlabel metal2 3416 41160 3416 41160 0 _0678_
rlabel metal2 22568 42560 22568 42560 0 _0679_
rlabel metal2 22456 44464 22456 44464 0 _0680_
rlabel metal2 2744 51800 2744 51800 0 _0681_
rlabel metal2 23016 43176 23016 43176 0 _0682_
rlabel metal2 25480 40208 25480 40208 0 _0683_
rlabel metal2 27384 36232 27384 36232 0 _0684_
rlabel metal2 33992 36904 33992 36904 0 _0685_
rlabel metal2 28392 42784 28392 42784 0 _0686_
rlabel metal2 28840 42224 28840 42224 0 _0687_
rlabel metal2 28728 53312 28728 53312 0 _0688_
rlabel metal3 22568 44296 22568 44296 0 _0689_
rlabel metal3 5824 50344 5824 50344 0 _0690_
rlabel metal3 19376 50008 19376 50008 0 _0691_
rlabel metal2 38808 48160 38808 48160 0 _0692_
rlabel metal2 19656 49616 19656 49616 0 _0693_
rlabel metal2 16072 54824 16072 54824 0 _0694_
rlabel metal2 19712 46872 19712 46872 0 _0695_
rlabel metal3 20664 45192 20664 45192 0 _0696_
rlabel metal3 6944 48328 6944 48328 0 _0697_
rlabel metal2 33264 53704 33264 53704 0 _0698_
rlabel metal2 1848 52080 1848 52080 0 _0699_
rlabel metal2 32984 56000 32984 56000 0 _0700_
rlabel metal2 15736 45528 15736 45528 0 _0701_
rlabel metal3 18816 45304 18816 45304 0 _0702_
rlabel metal2 10920 44072 10920 44072 0 _0703_
rlabel metal2 27384 51464 27384 51464 0 _0704_
rlabel metal2 18256 49000 18256 49000 0 _0705_
rlabel metal2 17976 42672 17976 42672 0 _0706_
rlabel metal3 19320 42952 19320 42952 0 _0707_
rlabel metal3 20776 44520 20776 44520 0 _0708_
rlabel metal2 21672 44128 21672 44128 0 _0709_
rlabel metal2 29512 42112 29512 42112 0 _0710_
rlabel metal2 35952 37240 35952 37240 0 _0711_
rlabel metal2 39256 36064 39256 36064 0 _0712_
rlabel metal2 39144 36120 39144 36120 0 _0713_
rlabel metal2 35112 36568 35112 36568 0 _0714_
rlabel metal2 35504 37352 35504 37352 0 _0715_
rlabel metal3 40096 36232 40096 36232 0 _0716_
rlabel metal3 33264 35672 33264 35672 0 _0717_
rlabel metal3 34328 40488 34328 40488 0 _0718_
rlabel metal2 25704 49896 25704 49896 0 _0719_
rlabel metal2 32200 51632 32200 51632 0 _0720_
rlabel metal2 9912 41776 9912 41776 0 _0721_
rlabel metal2 12376 39200 12376 39200 0 _0722_
rlabel metal2 8904 42840 8904 42840 0 _0723_
rlabel metal3 13888 39592 13888 39592 0 _0724_
rlabel metal2 21784 41776 21784 41776 0 _0725_
rlabel metal2 16072 42224 16072 42224 0 _0726_
rlabel metal2 16520 38976 16520 38976 0 _0727_
rlabel metal2 24584 40936 24584 40936 0 _0728_
rlabel metal3 20496 39368 20496 39368 0 _0729_
rlabel metal2 7168 45080 7168 45080 0 _0730_
rlabel metal2 19096 40320 19096 40320 0 _0731_
rlabel metal2 23016 40376 23016 40376 0 _0732_
rlabel metal2 23128 40096 23128 40096 0 _0733_
rlabel metal2 34216 39928 34216 39928 0 _0734_
rlabel metal2 33768 39256 33768 39256 0 _0735_
rlabel metal2 36568 38808 36568 38808 0 _0736_
rlabel metal2 37800 38920 37800 38920 0 _0737_
rlabel metal3 18872 38808 18872 38808 0 _0738_
rlabel metal2 6664 47152 6664 47152 0 _0739_
rlabel metal3 17248 38696 17248 38696 0 _0740_
rlabel metal2 11368 39704 11368 39704 0 _0741_
rlabel metal3 16576 48328 16576 48328 0 _0742_
rlabel metal3 17640 24136 17640 24136 0 _0743_
rlabel metal2 11144 39648 11144 39648 0 _0744_
rlabel metal2 19656 39032 19656 39032 0 _0745_
rlabel metal3 23744 38808 23744 38808 0 _0746_
rlabel metal2 27272 37856 27272 37856 0 _0747_
rlabel metal3 26992 38024 26992 38024 0 _0748_
rlabel metal3 39312 38808 39312 38808 0 _0749_
rlabel metal3 26376 42056 26376 42056 0 _0750_
rlabel metal2 26488 42112 26488 42112 0 _0751_
rlabel metal2 29848 41608 29848 41608 0 _0752_
rlabel metal3 17920 41944 17920 41944 0 _0753_
rlabel metal3 18312 41384 18312 41384 0 _0754_
rlabel metal3 11704 42728 11704 42728 0 _0755_
rlabel metal2 25928 49168 25928 49168 0 _0756_
rlabel metal2 7336 42392 7336 42392 0 _0757_
rlabel metal3 8372 23352 8372 23352 0 _0758_
rlabel metal2 32704 54712 32704 54712 0 _0759_
rlabel metal2 12712 42504 12712 42504 0 _0760_
rlabel metal2 33936 55048 33936 55048 0 _0761_
rlabel metal2 16464 42952 16464 42952 0 _0762_
rlabel metal2 16408 43792 16408 43792 0 _0763_
rlabel metal2 17920 41944 17920 41944 0 _0764_
rlabel metal2 25256 42280 25256 42280 0 _0765_
rlabel metal2 29848 40488 29848 40488 0 _0766_
rlabel metal2 39480 38136 39480 38136 0 _0767_
rlabel metal2 40152 37184 40152 37184 0 _0768_
rlabel metal2 42224 53704 42224 53704 0 _0769_
rlabel metal2 41720 36960 41720 36960 0 _0770_
rlabel metal2 41552 36680 41552 36680 0 _0771_
rlabel metal2 42616 38528 42616 38528 0 _0772_
rlabel metal2 38696 37800 38696 37800 0 _0773_
rlabel metal2 39480 39200 39480 39200 0 _0774_
rlabel metal2 38920 39312 38920 39312 0 _0775_
rlabel metal3 39984 39592 39984 39592 0 _0776_
rlabel metal3 2744 46872 2744 46872 0 _0777_
rlabel metal2 2072 44688 2072 44688 0 _0778_
rlabel metal2 12600 47208 12600 47208 0 _0779_
rlabel metal2 13160 44520 13160 44520 0 _0780_
rlabel metal2 12656 43512 12656 43512 0 _0781_
rlabel metal2 13664 45864 13664 45864 0 _0782_
rlabel metal2 2856 52360 2856 52360 0 _0783_
rlabel metal2 18648 46536 18648 46536 0 _0784_
rlabel metal2 12712 45920 12712 45920 0 _0785_
rlabel metal3 13664 45304 13664 45304 0 _0786_
rlabel metal2 39424 53144 39424 53144 0 _0787_
rlabel metal2 13944 45920 13944 45920 0 _0788_
rlabel metal2 9016 47768 9016 47768 0 _0789_
rlabel metal3 6272 45976 6272 45976 0 _0790_
rlabel metal3 40936 52136 40936 52136 0 _0791_
rlabel metal3 4704 48216 4704 48216 0 _0792_
rlabel metal2 3192 49784 3192 49784 0 _0793_
rlabel metal2 38696 47824 38696 47824 0 _0794_
rlabel metal2 39088 50008 39088 50008 0 _0795_
rlabel metal2 3752 49448 3752 49448 0 _0796_
rlabel metal3 4592 48440 4592 48440 0 _0797_
rlabel metal2 5432 46928 5432 46928 0 _0798_
rlabel metal2 25368 44520 25368 44520 0 _0799_
rlabel metal3 13608 41720 13608 41720 0 _0800_
rlabel metal2 14392 42392 14392 42392 0 _0801_
rlabel metal2 6552 42112 6552 42112 0 _0802_
rlabel metal3 22904 42840 22904 42840 0 _0803_
rlabel metal2 26712 43288 26712 43288 0 _0804_
rlabel metal2 28056 44016 28056 44016 0 _0805_
rlabel metal2 28168 43960 28168 43960 0 _0806_
rlabel metal2 40040 40824 40040 40824 0 _0807_
rlabel metal2 39256 41552 39256 41552 0 _0808_
rlabel metal2 3192 50848 3192 50848 0 _0809_
rlabel metal2 38360 56952 38360 56952 0 _0810_
rlabel metal2 40824 52248 40824 52248 0 _0811_
rlabel metal2 2072 53872 2072 53872 0 _0812_
rlabel metal3 15344 21560 15344 21560 0 _0813_
rlabel metal2 24136 41384 24136 41384 0 _0814_
rlabel metal2 31584 38248 31584 38248 0 _0815_
rlabel metal3 31976 55832 31976 55832 0 _0816_
rlabel metal3 15960 49784 15960 49784 0 _0817_
rlabel metal2 18256 44408 18256 44408 0 _0818_
rlabel metal2 22680 43512 22680 43512 0 _0819_
rlabel metal3 9296 46872 9296 46872 0 _0820_
rlabel metal2 8792 46900 8792 46900 0 _0821_
rlabel metal2 9128 45864 9128 45864 0 _0822_
rlabel metal2 10136 45248 10136 45248 0 _0823_
rlabel metal2 10416 41720 10416 41720 0 _0824_
rlabel metal3 31304 42056 31304 42056 0 _0825_
rlabel metal3 33208 42056 33208 42056 0 _0826_
rlabel metal2 34552 43456 34552 43456 0 _0827_
rlabel metal2 35000 42504 35000 42504 0 _0828_
rlabel metal3 34888 42056 34888 42056 0 _0829_
rlabel metal3 33656 51464 33656 51464 0 _0830_
rlabel metal2 37464 42168 37464 42168 0 _0831_
rlabel metal2 38920 42056 38920 42056 0 _0832_
rlabel metal2 36288 44296 36288 44296 0 _0833_
rlabel metal3 34888 50568 34888 50568 0 _0834_
rlabel metal2 34328 45528 34328 45528 0 _0835_
rlabel metal2 34888 43064 34888 43064 0 _0836_
rlabel metal2 35616 43512 35616 43512 0 _0837_
rlabel metal2 39928 43120 39928 43120 0 _0838_
rlabel metal2 27048 50848 27048 50848 0 _0839_
rlabel metal3 27944 38808 27944 38808 0 _0840_
rlabel metal3 9016 40264 9016 40264 0 _0841_
rlabel metal4 6776 42672 6776 42672 0 _0842_
rlabel metal2 20104 46536 20104 46536 0 _0843_
rlabel metal2 9072 44968 9072 44968 0 _0844_
rlabel metal2 1960 43344 1960 43344 0 _0845_
rlabel metal2 9016 40040 9016 40040 0 _0846_
rlabel metal2 9912 40880 9912 40880 0 _0847_
rlabel metal2 25928 40152 25928 40152 0 _0848_
rlabel metal2 38696 40936 38696 40936 0 _0849_
rlabel metal2 40600 41384 40600 41384 0 _0850_
rlabel metal2 38808 44856 38808 44856 0 _0851_
rlabel metal2 40488 40992 40488 40992 0 _0852_
rlabel metal2 41832 40320 41832 40320 0 _0853_
rlabel metal2 42504 39200 42504 39200 0 _0854_
rlabel metal2 2744 4480 2744 4480 0 _0855_
rlabel metal2 26376 43736 26376 43736 0 _0856_
rlabel metal2 27776 50456 27776 50456 0 _0857_
rlabel metal3 27664 45080 27664 45080 0 _0858_
rlabel metal3 17472 47432 17472 47432 0 _0859_
rlabel metal3 11648 48328 11648 48328 0 _0860_
rlabel metal3 13608 47656 13608 47656 0 _0861_
rlabel metal3 15848 47432 15848 47432 0 _0862_
rlabel metal2 10696 40824 10696 40824 0 _0863_
rlabel metal3 15792 40376 15792 40376 0 _0864_
rlabel metal2 16912 49112 16912 49112 0 _0865_
rlabel metal2 20104 48216 20104 48216 0 _0866_
rlabel metal2 17024 48888 17024 48888 0 _0867_
rlabel metal4 15904 46200 15904 46200 0 _0868_
rlabel metal3 16912 46872 16912 46872 0 _0869_
rlabel metal2 16520 47152 16520 47152 0 _0870_
rlabel metal2 26712 44744 26712 44744 0 _0871_
rlabel metal3 27720 45192 27720 45192 0 _0872_
rlabel metal2 42392 44520 42392 44520 0 _0873_
rlabel metal2 32648 43960 32648 43960 0 _0874_
rlabel metal2 34160 47320 34160 47320 0 _0875_
rlabel metal2 20328 55440 20328 55440 0 _0876_
rlabel metal2 18984 51240 18984 51240 0 _0877_
rlabel metal2 13776 48216 13776 48216 0 _0878_
rlabel metal2 14280 52472 14280 52472 0 _0879_
rlabel metal2 25816 54936 25816 54936 0 _0880_
rlabel metal2 10696 53424 10696 53424 0 _0881_
rlabel metal2 11256 53200 11256 53200 0 _0882_
rlabel metal2 30296 52752 30296 52752 0 _0883_
rlabel metal2 41944 52752 41944 52752 0 _0884_
rlabel metal2 31304 56336 31304 56336 0 _0885_
rlabel metal3 28952 54432 28952 54432 0 _0886_
rlabel metal4 33768 51464 33768 51464 0 _0887_
rlabel metal2 11032 54544 11032 54544 0 _0888_
rlabel metal2 12712 53704 12712 53704 0 _0889_
rlabel metal3 32200 21728 32200 21728 0 _0890_
rlabel metal2 35784 45192 35784 45192 0 _0891_
rlabel metal3 35280 45080 35280 45080 0 _0892_
rlabel metal2 38696 43596 38696 43596 0 _0893_
rlabel metal2 29624 43288 29624 43288 0 _0894_
rlabel metal2 29960 44688 29960 44688 0 _0895_
rlabel metal2 21560 49448 21560 49448 0 _0896_
rlabel metal2 11480 50904 11480 50904 0 _0897_
rlabel metal2 10472 48048 10472 48048 0 _0898_
rlabel metal2 11032 50344 11032 50344 0 _0899_
rlabel metal3 6608 52920 6608 52920 0 _0900_
rlabel metal3 8624 51576 8624 51576 0 _0901_
rlabel metal2 10024 50848 10024 50848 0 _0902_
rlabel metal3 11200 51240 11200 51240 0 _0903_
rlabel metal2 16072 47488 16072 47488 0 _0904_
rlabel metal2 39704 43624 39704 43624 0 _0905_
rlabel metal2 42728 44800 42728 44800 0 _0906_
rlabel metal3 41664 53032 41664 53032 0 _0907_
rlabel metal2 42840 43988 42840 43988 0 _0908_
rlabel metal2 44184 43120 44184 43120 0 _0909_
rlabel metal2 44072 44688 44072 44688 0 _0910_
rlabel metal2 44128 41944 44128 41944 0 _0911_
rlabel metal2 40264 42280 40264 42280 0 _0912_
rlabel metal2 44016 41720 44016 41720 0 _0913_
rlabel metal2 43064 41384 43064 41384 0 _0914_
rlabel metal3 44800 41160 44800 41160 0 _0915_
rlabel metal2 44072 39536 44072 39536 0 _0916_
rlabel metal2 41608 39648 41608 39648 0 _0917_
rlabel metal3 44128 40488 44128 40488 0 _0918_
rlabel metal3 43232 40376 43232 40376 0 _0919_
rlabel metal3 44744 40600 44744 40600 0 _0920_
rlabel metal2 2744 10752 2744 10752 0 _0921_
rlabel via2 44184 44408 44184 44408 0 _0922_
rlabel metal2 37016 44744 37016 44744 0 _0923_
rlabel metal2 21336 47992 21336 47992 0 _0924_
rlabel metal3 19824 49672 19824 49672 0 _0925_
rlabel metal3 22568 45080 22568 45080 0 _0926_
rlabel metal2 31080 45416 31080 45416 0 _0927_
rlabel metal3 11984 44968 11984 44968 0 _0928_
rlabel metal2 23688 46536 23688 46536 0 _0929_
rlabel metal2 31864 45360 31864 45360 0 _0930_
rlabel metal2 31976 44352 31976 44352 0 _0931_
rlabel metal3 33264 44520 33264 44520 0 _0932_
rlabel metal2 39480 45696 39480 45696 0 _0933_
rlabel metal2 37352 44576 37352 44576 0 _0934_
rlabel metal2 39480 50736 39480 50736 0 _0935_
rlabel metal2 20328 48216 20328 48216 0 _0936_
rlabel metal2 2016 50008 2016 50008 0 _0937_
rlabel metal2 20216 48440 20216 48440 0 _0938_
rlabel metal3 18984 47432 18984 47432 0 _0939_
rlabel metal2 26152 47040 26152 47040 0 _0940_
rlabel metal3 30072 47544 30072 47544 0 _0941_
rlabel metal2 39256 47432 39256 47432 0 _0942_
rlabel metal2 21784 50456 21784 50456 0 _0943_
rlabel metal2 3752 54768 3752 54768 0 _0944_
rlabel metal3 21840 49896 21840 49896 0 _0945_
rlabel metal2 23912 47824 23912 47824 0 _0946_
rlabel metal2 24472 47768 24472 47768 0 _0947_
rlabel metal2 23576 51632 23576 51632 0 _0948_
rlabel metal3 20832 48216 20832 48216 0 _0949_
rlabel metal2 21672 48608 21672 48608 0 _0950_
rlabel metal3 23968 48776 23968 48776 0 _0951_
rlabel metal2 26712 48160 26712 48160 0 _0952_
rlabel metal2 25704 46256 25704 46256 0 _0953_
rlabel metal2 27160 46816 27160 46816 0 _0954_
rlabel metal2 27664 46872 27664 46872 0 _0955_
rlabel metal3 27720 47432 27720 47432 0 _0956_
rlabel metal2 40600 46984 40600 46984 0 _0957_
rlabel metal2 43960 44688 43960 44688 0 _0958_
rlabel metal3 45416 43512 45416 43512 0 _0959_
rlabel metal3 45136 44296 45136 44296 0 _0960_
rlabel metal2 45416 41832 45416 41832 0 _0961_
rlabel metal3 45248 42728 45248 42728 0 _0962_
rlabel metal2 45752 40656 45752 40656 0 _0963_
rlabel metal2 47544 39928 47544 39928 0 _0964_
rlabel metal2 32760 45948 32760 45948 0 _0965_
rlabel metal3 4760 50344 4760 50344 0 _0966_
rlabel metal2 16072 50344 16072 50344 0 _0967_
rlabel metal2 15736 51016 15736 51016 0 _0968_
rlabel metal2 14504 43008 14504 43008 0 _0969_
rlabel metal3 15232 43624 15232 43624 0 _0970_
rlabel metal3 17304 51352 17304 51352 0 _0971_
rlabel metal3 20664 51016 20664 51016 0 _0972_
rlabel metal3 34552 47432 34552 47432 0 _0973_
rlabel metal2 34888 47432 34888 47432 0 _0974_
rlabel metal2 37240 47040 37240 47040 0 _0975_
rlabel metal2 30072 51744 30072 51744 0 _0976_
rlabel metal2 28056 53032 28056 53032 0 _0977_
rlabel metal2 12824 47992 12824 47992 0 _0978_
rlabel metal2 21112 48048 21112 48048 0 _0979_
rlabel metal2 23352 47600 23352 47600 0 _0980_
rlabel metal3 33432 48440 33432 48440 0 _0981_
rlabel metal2 37800 48384 37800 48384 0 _0982_
rlabel metal2 37912 47992 37912 47992 0 _0983_
rlabel metal2 15288 54376 15288 54376 0 _0984_
rlabel metal2 18312 52528 18312 52528 0 _0985_
rlabel metal3 20160 51912 20160 51912 0 _0986_
rlabel metal3 13104 51352 13104 51352 0 _0987_
rlabel metal2 13888 51240 13888 51240 0 _0988_
rlabel metal3 18144 51240 18144 51240 0 _0989_
rlabel metal2 29848 50904 29848 50904 0 _0990_
rlabel metal3 24920 47320 24920 47320 0 _0991_
rlabel metal2 27496 50484 27496 50484 0 _0992_
rlabel metal3 28784 50680 28784 50680 0 _0993_
rlabel metal2 30800 50456 30800 50456 0 _0994_
rlabel via2 40152 49000 40152 49000 0 _0995_
rlabel metal2 40040 48440 40040 48440 0 _0996_
rlabel metal2 41608 47432 41608 47432 0 _0997_
rlabel metal2 40040 45136 40040 45136 0 _0998_
rlabel metal3 40040 45976 40040 45976 0 _0999_
rlabel metal2 40152 45472 40152 45472 0 _1000_
rlabel metal2 41048 47320 41048 47320 0 _1001_
rlabel metal3 44968 48328 44968 48328 0 _1002_
rlabel metal2 44072 46368 44072 46368 0 _1003_
rlabel metal2 46088 43960 46088 43960 0 _1004_
rlabel metal3 44968 45752 44968 45752 0 _1005_
rlabel metal2 44688 46648 44688 46648 0 _1006_
rlabel metal2 43736 46984 43736 46984 0 _1007_
rlabel metal2 36792 49616 36792 49616 0 _1008_
rlabel metal2 34888 51296 34888 51296 0 _1009_
rlabel metal2 40264 48944 40264 48944 0 _1010_
rlabel metal2 32424 50848 32424 50848 0 _1011_
rlabel metal2 9856 53704 9856 53704 0 _1012_
rlabel metal2 8344 52752 8344 52752 0 _1013_
rlabel metal2 43568 53704 43568 53704 0 _1014_
rlabel metal2 8904 52808 8904 52808 0 _1015_
rlabel metal2 8120 51800 8120 51800 0 _1016_
rlabel metal2 8680 51576 8680 51576 0 _1017_
rlabel metal3 31360 51352 31360 51352 0 _1018_
rlabel metal3 34440 51128 34440 51128 0 _1019_
rlabel metal2 33656 40040 33656 40040 0 _1020_
rlabel metal2 35448 51184 35448 51184 0 _1021_
rlabel metal3 37464 50456 37464 50456 0 _1022_
rlabel metal2 11480 52080 11480 52080 0 _1023_
rlabel metal2 20552 52192 20552 52192 0 _1024_
rlabel metal2 23688 52080 23688 52080 0 _1025_
rlabel metal2 24584 51856 24584 51856 0 _1026_
rlabel metal3 26712 52248 26712 52248 0 _1027_
rlabel metal2 30744 52192 30744 52192 0 _1028_
rlabel metal2 37912 50848 37912 50848 0 _1029_
rlabel metal3 28840 54936 28840 54936 0 _1030_
rlabel metal2 22064 53480 22064 53480 0 _1031_
rlabel metal2 22120 54992 22120 54992 0 _1032_
rlabel metal2 17640 54488 17640 54488 0 _1033_
rlabel metal2 19096 54656 19096 54656 0 _1034_
rlabel metal2 27216 50792 27216 50792 0 _1035_
rlabel metal2 27944 51072 27944 51072 0 _1036_
rlabel metal2 38808 50792 38808 50792 0 _1037_
rlabel metal2 40600 50064 40600 50064 0 _1038_
rlabel metal3 41888 49672 41888 49672 0 _1039_
rlabel metal3 41944 48888 41944 48888 0 _1040_
rlabel metal2 43960 47880 43960 47880 0 _1041_
rlabel metal2 41608 48496 41608 48496 0 _1042_
rlabel metal2 43400 48496 43400 48496 0 _1043_
rlabel metal3 44520 48104 44520 48104 0 _1044_
rlabel metal2 43512 47768 43512 47768 0 _1045_
rlabel metal2 3192 4536 3192 4536 0 _1046_
rlabel metal2 20440 46368 20440 46368 0 _1047_
rlabel metal3 20776 48552 20776 48552 0 _1048_
rlabel metal2 20496 53928 20496 53928 0 _1049_
rlabel metal2 15064 54488 15064 54488 0 _1050_
rlabel metal2 16184 54880 16184 54880 0 _1051_
rlabel metal2 15176 54880 15176 54880 0 _1052_
rlabel metal3 18648 54488 18648 54488 0 _1053_
rlabel metal2 31304 51800 31304 51800 0 _1054_
rlabel metal2 32536 52248 32536 52248 0 _1055_
rlabel metal3 33096 50792 33096 50792 0 _1056_
rlabel metal3 35560 50792 35560 50792 0 _1057_
rlabel metal2 41608 50848 41608 50848 0 _1058_
rlabel metal2 19488 51576 19488 51576 0 _1059_
rlabel metal3 24920 53704 24920 53704 0 _1060_
rlabel metal2 26600 50960 26600 50960 0 _1061_
rlabel metal2 26488 50120 26488 50120 0 _1062_
rlabel metal2 40880 50344 40880 50344 0 _1063_
rlabel metal2 42952 50960 42952 50960 0 _1064_
rlabel metal2 28056 54880 28056 54880 0 _1065_
rlabel metal2 19880 49392 19880 49392 0 _1066_
rlabel metal2 21728 53704 21728 53704 0 _1067_
rlabel metal3 27328 54600 27328 54600 0 _1068_
rlabel metal2 28728 54432 28728 54432 0 _1069_
rlabel metal2 27944 53928 27944 53928 0 _1070_
rlabel metal2 45864 51240 45864 51240 0 _1071_
rlabel metal2 38920 51688 38920 51688 0 _1072_
rlabel metal3 38976 51352 38976 51352 0 _1073_
rlabel metal2 46088 51296 46088 51296 0 _1074_
rlabel metal2 46536 49840 46536 49840 0 _1075_
rlabel metal3 45360 47432 45360 47432 0 _1076_
rlabel metal3 45416 48888 45416 48888 0 _1077_
rlabel metal2 43960 49280 43960 49280 0 _1078_
rlabel metal2 45528 48832 45528 48832 0 _1079_
rlabel metal2 46648 48944 46648 48944 0 _1080_
rlabel metal3 52808 48888 52808 48888 0 _1081_
rlabel metal2 42168 50680 42168 50680 0 _1082_
rlabel metal2 44856 52136 44856 52136 0 _1083_
rlabel metal2 22904 32648 22904 32648 0 _1084_
rlabel metal2 18592 46872 18592 46872 0 _1085_
rlabel metal3 18592 53592 18592 53592 0 _1086_
rlabel metal3 21000 53480 21000 53480 0 _1087_
rlabel metal2 22624 53144 22624 53144 0 _1088_
rlabel metal2 30912 50568 30912 50568 0 _1089_
rlabel metal2 32760 48776 32760 48776 0 _1090_
rlabel metal2 33656 53200 33656 53200 0 _1091_
rlabel metal3 33208 53144 33208 53144 0 _1092_
rlabel metal3 23800 52024 23800 52024 0 _1093_
rlabel metal2 26712 52640 26712 52640 0 _1094_
rlabel metal2 27384 52808 27384 52808 0 _1095_
rlabel metal2 31976 53760 31976 53760 0 _1096_
rlabel metal2 31864 54432 31864 54432 0 _1097_
rlabel metal2 31640 54992 31640 54992 0 _1098_
rlabel metal2 27160 54936 27160 54936 0 _1099_
rlabel metal2 24920 55552 24920 55552 0 _1100_
rlabel metal2 28280 54600 28280 54600 0 _1101_
rlabel metal2 17304 53704 17304 53704 0 _1102_
rlabel metal2 17864 53760 17864 53760 0 _1103_
rlabel metal2 28504 54488 28504 54488 0 _1104_
rlabel metal2 30744 54880 30744 54880 0 _1105_
rlabel metal2 30632 54208 30632 54208 0 _1106_
rlabel metal2 31752 54824 31752 54824 0 _1107_
rlabel metal2 44520 53144 44520 53144 0 _1108_
rlabel metal3 45416 52360 45416 52360 0 _1109_
rlabel metal2 45752 52416 45752 52416 0 _1110_
rlabel metal2 45976 53200 45976 53200 0 _1111_
rlabel metal2 46200 53592 46200 53592 0 _1112_
rlabel metal3 34888 51352 34888 51352 0 _1113_
rlabel metal2 35896 52192 35896 52192 0 _1114_
rlabel metal3 20048 51464 20048 51464 0 _1115_
rlabel metal3 28616 52024 28616 52024 0 _1116_
rlabel metal2 36400 52920 36400 52920 0 _1117_
rlabel metal2 37800 53312 37800 53312 0 _1118_
rlabel metal2 26376 52304 26376 52304 0 _1119_
rlabel metal2 27496 52416 27496 52416 0 _1120_
rlabel metal2 37576 54096 37576 54096 0 _1121_
rlabel metal2 38808 54768 38808 54768 0 _1122_
rlabel metal2 28504 55720 28504 55720 0 _1123_
rlabel metal3 29288 53704 29288 53704 0 _1124_
rlabel metal2 29736 53704 29736 53704 0 _1125_
rlabel metal2 30520 54096 30520 54096 0 _1126_
rlabel metal2 35896 54376 35896 54376 0 _1127_
rlabel metal3 40712 54488 40712 54488 0 _1128_
rlabel metal2 34160 53928 34160 53928 0 _1129_
rlabel metal3 43960 54600 43960 54600 0 _1130_
rlabel metal2 42952 54936 42952 54936 0 _1131_
rlabel metal3 44688 52136 44688 52136 0 _1132_
rlabel metal2 45976 51632 45976 51632 0 _1133_
rlabel metal2 44856 55048 44856 55048 0 _1134_
rlabel metal3 39312 55160 39312 55160 0 _1135_
rlabel metal3 38640 53816 38640 53816 0 _1136_
rlabel metal3 39480 55272 39480 55272 0 _1137_
rlabel metal2 24192 50344 24192 50344 0 _1138_
rlabel metal3 25732 49784 25732 49784 0 _1139_
rlabel metal2 32032 50456 32032 50456 0 _1140_
rlabel metal3 33152 51352 33152 51352 0 _1141_
rlabel metal3 35224 53480 35224 53480 0 _1142_
rlabel metal2 39368 54992 39368 54992 0 _1143_
rlabel metal3 40600 55048 40600 55048 0 _1144_
rlabel metal2 40824 54936 40824 54936 0 _1145_
rlabel metal2 45752 54656 45752 54656 0 _1146_
rlabel metal2 44072 54768 44072 54768 0 _1147_
rlabel metal3 45248 55384 45248 55384 0 _1148_
rlabel metal3 46928 55160 46928 55160 0 _1149_
rlabel metal2 42168 53256 42168 53256 0 _1150_
rlabel metal3 40432 53592 40432 53592 0 _1151_
rlabel metal2 41832 53032 41832 53032 0 _1152_
rlabel metal2 35840 53032 35840 53032 0 _1153_
rlabel metal2 35672 53144 35672 53144 0 _1154_
rlabel metal3 38808 52920 38808 52920 0 _1155_
rlabel metal2 48440 51296 48440 51296 0 _1156_
rlabel metal2 47936 31752 47936 31752 0 _1157_
rlabel metal2 47096 27552 47096 27552 0 _1158_
rlabel metal2 49448 26096 49448 26096 0 _1159_
rlabel metal2 50456 31248 50456 31248 0 _1160_
rlabel metal2 49728 29624 49728 29624 0 _1161_
rlabel metal2 49784 29288 49784 29288 0 _1162_
rlabel metal2 50120 27048 50120 27048 0 _1163_
rlabel metal3 39032 20776 39032 20776 0 _1164_
rlabel metal2 45360 29960 45360 29960 0 _1165_
rlabel metal2 52528 31752 52528 31752 0 _1166_
rlabel metal2 44744 30296 44744 30296 0 _1167_
rlabel metal2 44520 30632 44520 30632 0 _1168_
rlabel metal2 48160 31080 48160 31080 0 _1169_
rlabel metal2 56280 25480 56280 25480 0 _1170_
rlabel metal2 44240 27384 44240 27384 0 _1171_
rlabel metal2 48552 30016 48552 30016 0 _1172_
rlabel metal2 46200 29568 46200 29568 0 _1173_
rlabel metal2 44072 28224 44072 28224 0 _1174_
rlabel metal3 57232 23352 57232 23352 0 _1175_
rlabel metal3 55888 23352 55888 23352 0 _1176_
rlabel metal2 46872 27776 46872 27776 0 _1177_
rlabel metal3 47096 27496 47096 27496 0 _1178_
rlabel metal2 43960 27048 43960 27048 0 _1179_
rlabel metal2 52584 17136 52584 17136 0 _1180_
rlabel metal2 55608 29792 55608 29792 0 _1181_
rlabel metal2 44856 26376 44856 26376 0 _1182_
rlabel metal3 44240 26040 44240 26040 0 _1183_
rlabel metal3 55776 21672 55776 21672 0 _1184_
rlabel metal3 54768 19096 54768 19096 0 _1185_
rlabel metal3 49336 14448 49336 14448 0 _1186_
rlabel metal2 52696 23744 52696 23744 0 _1187_
rlabel metal2 45416 19040 45416 19040 0 _1188_
rlabel metal3 54488 24808 54488 24808 0 _1189_
rlabel metal2 47152 15960 47152 15960 0 _1190_
rlabel metal2 50456 24640 50456 24640 0 _1191_
rlabel metal2 56840 20552 56840 20552 0 _1192_
rlabel metal2 51800 17192 51800 17192 0 _1193_
rlabel metal3 54432 13832 54432 13832 0 _1194_
rlabel metal2 46424 17528 46424 17528 0 _1195_
rlabel metal2 44408 12880 44408 12880 0 _1196_
rlabel metal2 47432 22512 47432 22512 0 _1197_
rlabel metal2 49896 12208 49896 12208 0 _1198_
rlabel metal2 49560 12432 49560 12432 0 _1199_
rlabel metal2 45136 7672 45136 7672 0 _1200_
rlabel metal3 47096 26936 47096 26936 0 _1201_
rlabel metal3 44912 14392 44912 14392 0 _1202_
rlabel metal2 49672 28112 49672 28112 0 _1203_
rlabel metal2 47544 24360 47544 24360 0 _1204_
rlabel metal2 52584 22288 52584 22288 0 _1205_
rlabel metal2 43176 27496 43176 27496 0 _1206_
rlabel metal2 43288 14504 43288 14504 0 _1207_
rlabel metal2 44072 14112 44072 14112 0 _1208_
rlabel metal3 45360 12264 45360 12264 0 _1209_
rlabel metal3 43960 10024 43960 10024 0 _1210_
rlabel metal2 42672 6104 42672 6104 0 _1211_
rlabel metal2 44408 6328 44408 6328 0 _1212_
rlabel metal2 45640 7560 45640 7560 0 _1213_
rlabel metal3 56112 15288 56112 15288 0 _1214_
rlabel metal2 53592 10976 53592 10976 0 _1215_
rlabel metal2 48888 28616 48888 28616 0 _1216_
rlabel metal2 48216 14112 48216 14112 0 _1217_
rlabel metal2 49336 28560 49336 28560 0 _1218_
rlabel metal2 50344 7616 50344 7616 0 _1219_
rlabel metal2 55272 19712 55272 19712 0 _1220_
rlabel metal2 54824 15568 54824 15568 0 _1221_
rlabel metal3 41608 12264 41608 12264 0 _1222_
rlabel metal2 54040 12208 54040 12208 0 _1223_
rlabel metal3 53088 10696 53088 10696 0 _1224_
rlabel metal2 32648 20944 32648 20944 0 _1225_
rlabel metal2 46200 21896 46200 21896 0 _1226_
rlabel metal2 54264 21224 54264 21224 0 _1227_
rlabel metal3 34160 15960 34160 15960 0 _1228_
rlabel metal2 45976 23576 45976 23576 0 _1229_
rlabel metal2 53424 12376 53424 12376 0 _1230_
rlabel metal2 57736 21840 57736 21840 0 _1231_
rlabel metal3 42896 16184 42896 16184 0 _1232_
rlabel metal2 53704 24192 53704 24192 0 _1233_
rlabel metal3 49448 18704 49448 18704 0 _1234_
rlabel metal2 52080 23352 52080 23352 0 _1235_
rlabel metal2 54264 29960 54264 29960 0 _1236_
rlabel metal3 48692 23912 48692 23912 0 _1237_
rlabel metal2 46088 17696 46088 17696 0 _1238_
rlabel metal2 46760 18368 46760 18368 0 _1239_
rlabel metal3 53760 12152 53760 12152 0 _1240_
rlabel metal2 52920 10976 52920 10976 0 _1241_
rlabel metal2 52864 9016 52864 9016 0 _1242_
rlabel metal2 48048 8008 48048 8008 0 _1243_
rlabel metal2 39592 21560 39592 21560 0 _1244_
rlabel metal3 49784 25256 49784 25256 0 _1245_
rlabel metal3 47992 20776 47992 20776 0 _1246_
rlabel metal2 48552 28672 48552 28672 0 _1247_
rlabel metal3 51800 20776 51800 20776 0 _1248_
rlabel metal3 48608 29288 48608 29288 0 _1249_
rlabel metal2 48328 21784 48328 21784 0 _1250_
rlabel metal2 49560 21784 49560 21784 0 _1251_
rlabel metal2 44128 21560 44128 21560 0 _1252_
rlabel metal2 48216 18704 48216 18704 0 _1253_
rlabel metal3 49112 21000 49112 21000 0 _1254_
rlabel metal4 48664 27496 48664 27496 0 _1255_
rlabel metal3 48496 18536 48496 18536 0 _1256_
rlabel metal2 47992 8960 47992 8960 0 _1257_
rlabel metal3 52192 32648 52192 32648 0 _1258_
rlabel metal2 46872 7840 46872 7840 0 _1259_
rlabel metal2 48104 8288 48104 8288 0 _1260_
rlabel metal2 55048 8624 55048 8624 0 _1261_
rlabel metal2 55944 7448 55944 7448 0 _1262_
rlabel metal2 52808 7784 52808 7784 0 _1263_
rlabel metal2 53256 7728 53256 7728 0 _1264_
rlabel metal2 46984 11704 46984 11704 0 _1265_
rlabel metal2 39368 21728 39368 21728 0 _1266_
rlabel metal2 47544 15960 47544 15960 0 _1267_
rlabel metal3 52584 28504 52584 28504 0 _1268_
rlabel metal2 47096 15148 47096 15148 0 _1269_
rlabel metal4 47208 15708 47208 15708 0 _1270_
rlabel metal2 47992 14224 47992 14224 0 _1271_
rlabel metal2 47208 12712 47208 12712 0 _1272_
rlabel metal2 45528 17360 45528 17360 0 _1273_
rlabel metal2 45752 11928 45752 11928 0 _1274_
rlabel metal2 46536 29848 46536 29848 0 _1275_
rlabel metal3 46088 29512 46088 29512 0 _1276_
rlabel metal2 44800 29176 44800 29176 0 _1277_
rlabel metal2 50288 24696 50288 24696 0 _1278_
rlabel metal2 56616 24920 56616 24920 0 _1279_
rlabel metal2 44184 16408 44184 16408 0 _1280_
rlabel metal3 46704 15848 46704 15848 0 _1281_
rlabel metal2 44016 17080 44016 17080 0 _1282_
rlabel metal2 48552 24360 48552 24360 0 _1283_
rlabel metal3 45864 24696 45864 24696 0 _1284_
rlabel metal2 44968 15400 44968 15400 0 _1285_
rlabel metal2 44856 11872 44856 11872 0 _1286_
rlabel metal2 45080 9688 45080 9688 0 _1287_
rlabel metal2 44632 9296 44632 9296 0 _1288_
rlabel metal2 45528 6608 45528 6608 0 _1289_
rlabel metal3 38696 30072 38696 30072 0 _1290_
rlabel metal2 48216 6384 48216 6384 0 _1291_
rlabel metal2 48440 7056 48440 7056 0 _1292_
rlabel metal2 42728 7728 42728 7728 0 _1293_
rlabel metal3 48608 24808 48608 24808 0 _1294_
rlabel metal3 49392 16744 49392 16744 0 _1295_
rlabel metal2 48608 16296 48608 16296 0 _1296_
rlabel metal3 48552 27048 48552 27048 0 _1297_
rlabel metal2 49784 28336 49784 28336 0 _1298_
rlabel metal2 49448 27440 49448 27440 0 _1299_
rlabel metal3 49280 26936 49280 26936 0 _1300_
rlabel metal3 30352 20776 30352 20776 0 _1301_
rlabel metal2 52920 15680 52920 15680 0 _1302_
rlabel metal3 53760 15288 53760 15288 0 _1303_
rlabel metal2 50344 13104 50344 13104 0 _1304_
rlabel metal2 47880 8568 47880 8568 0 _1305_
rlabel metal3 47880 7672 47880 7672 0 _1306_
rlabel metal2 44408 7952 44408 7952 0 _1307_
rlabel metal2 47880 7504 47880 7504 0 _1308_
rlabel metal3 48888 6776 48888 6776 0 _1309_
rlabel metal3 51632 15400 51632 15400 0 _1310_
rlabel metal3 52192 15288 52192 15288 0 _1311_
rlabel metal2 50344 14112 50344 14112 0 _1312_
rlabel metal3 40152 14784 40152 14784 0 _1313_
rlabel metal3 51016 16296 51016 16296 0 _1314_
rlabel metal2 50176 15288 50176 15288 0 _1315_
rlabel metal2 45192 18200 45192 18200 0 _1316_
rlabel metal2 50568 15344 50568 15344 0 _1317_
rlabel metal2 50344 9296 50344 9296 0 _1318_
rlabel metal2 50232 11032 50232 11032 0 _1319_
rlabel metal2 50792 9072 50792 9072 0 _1320_
rlabel metal2 49784 8232 49784 8232 0 _1321_
rlabel metal2 53592 7168 53592 7168 0 _1322_
rlabel metal2 54152 12936 54152 12936 0 _1323_
rlabel metal2 33544 4592 33544 4592 0 _1324_
rlabel metal2 47992 6944 47992 6944 0 _1325_
rlabel metal3 49168 6104 49168 6104 0 _1326_
rlabel metal2 47992 5880 47992 5880 0 _1327_
rlabel metal2 28056 7224 28056 7224 0 _1328_
rlabel metal2 27160 7280 27160 7280 0 _1329_
rlabel metal2 26040 22848 26040 22848 0 _1330_
rlabel metal2 28056 18704 28056 18704 0 _1331_
rlabel metal2 46200 16240 46200 16240 0 _1332_
rlabel metal2 43848 30408 43848 30408 0 _1333_
rlabel metal2 51184 19432 51184 19432 0 _1334_
rlabel metal2 41160 27720 41160 27720 0 _1335_
rlabel metal3 48104 27832 48104 27832 0 _1336_
rlabel metal2 47936 25032 47936 25032 0 _1337_
rlabel metal2 46648 28784 46648 28784 0 _1338_
rlabel metal2 41944 27216 41944 27216 0 _1339_
rlabel metal2 41664 26824 41664 26824 0 _1340_
rlabel metal2 48664 25200 48664 25200 0 _1341_
rlabel metal3 40936 25592 40936 25592 0 _1342_
rlabel metal3 46480 28952 46480 28952 0 _1343_
rlabel metal2 44072 23072 44072 23072 0 _1344_
rlabel metal3 40432 2968 40432 2968 0 _1345_
rlabel metal3 17248 3416 17248 3416 0 addI[0]
rlabel metal3 1358 50456 1358 50456 0 addI[1]
rlabel metal3 57666 23576 57666 23576 0 addI[2]
rlabel metal2 27608 2198 27608 2198 0 addI[3]
rlabel metal2 55832 56672 55832 56672 0 addI[4]
rlabel metal3 56616 55384 56616 55384 0 addI[5]
rlabel metal3 18648 55944 18648 55944 0 addQ[0]
rlabel metal2 23576 57610 23576 57610 0 addQ[1]
rlabel metal2 39032 2058 39032 2058 0 addQ[2]
rlabel metal3 1358 27608 1358 27608 0 addQ[3]
rlabel metal3 1358 55832 1358 55832 0 addQ[4]
rlabel metal2 56056 29120 56056 29120 0 addQ[5]
rlabel metal2 19208 27776 19208 27776 0 gen_sym.Reg_2M.data_in
rlabel metal3 21448 25704 21448 25704 0 gen_sym.Reg_2M.data_out
rlabel metal2 17528 25368 17528 25368 0 gen_sym.Reg_2M.enable
rlabel metal3 25424 27608 25424 27608 0 gen_sym.Reg_Sym.data_out\[0\]
rlabel metal2 25032 26544 25032 26544 0 gen_sym.Reg_Sym.data_out\[1\]
rlabel metal2 25592 28504 25592 28504 0 mapper.bit_Q\[1\]
rlabel metal2 25816 55664 25816 55664 0 net1
rlabel metal3 56672 39480 56672 39480 0 net10
rlabel metal2 23688 3976 23688 3976 0 net11
rlabel metal3 32256 4424 32256 4424 0 net12
rlabel metal2 46760 44156 46760 44156 0 net13
rlabel metal2 2408 21504 2408 21504 0 net14
rlabel metal3 56672 45752 56672 45752 0 net15
rlabel metal2 2408 30240 2408 30240 0 net16
rlabel metal2 12488 3528 12488 3528 0 net17
rlabel metal3 3248 12376 3248 12376 0 net18
rlabel metal2 2408 17360 2408 17360 0 net19
rlabel metal3 2184 55944 2184 55944 0 net2
rlabel metal2 35784 55300 35784 55300 0 net20
rlabel metal3 50176 56056 50176 56056 0 net21
rlabel metal3 47656 52808 47656 52808 0 net22
rlabel metal2 48776 51856 48776 51856 0 net23
rlabel metal3 36568 56280 36568 56280 0 net24
rlabel metal2 2408 3976 2408 3976 0 net25
rlabel metal2 2408 11088 2408 11088 0 net26
rlabel metal2 47880 37632 47880 37632 0 net27
rlabel metal2 7224 55608 7224 55608 0 net28
rlabel metal2 2408 6160 2408 6160 0 net29
rlabel metal3 43400 3304 43400 3304 0 net3
rlabel metal2 50680 3976 50680 3976 0 net30
rlabel metal3 44072 54712 44072 54712 0 net31
rlabel metal2 48104 32480 48104 32480 0 net32
rlabel metal2 46648 32984 46648 32984 0 net33
rlabel metal2 40936 30688 40936 30688 0 net34
rlabel metal3 41328 1624 41328 1624 0 net35
rlabel metal3 51744 53816 51744 53816 0 net36
rlabel metal2 54320 55048 54320 55048 0 net37
rlabel metal2 17640 28448 17640 28448 0 net38
rlabel metal2 24416 39592 24416 39592 0 net39
rlabel metal2 43120 31080 43120 31080 0 net4
rlabel metal2 17080 24360 17080 24360 0 net40
rlabel metal2 3080 27944 3080 27944 0 net41
rlabel metal2 42560 49448 42560 49448 0 net42
rlabel metal3 43680 35616 43680 35616 0 net43
rlabel metal2 26376 38668 26376 38668 0 net44
rlabel metal3 25256 24024 25256 24024 0 net45
rlabel metal3 35560 5208 35560 5208 0 net46
rlabel metal2 26096 23800 26096 23800 0 net47
rlabel metal3 20160 26264 20160 26264 0 net48
rlabel metal2 27552 30968 27552 30968 0 net49
rlabel metal2 7000 8960 7000 8960 0 net5
rlabel metal3 15960 34776 15960 34776 0 net50
rlabel metal3 11592 30856 11592 30856 0 net51
rlabel metal3 21000 25256 21000 25256 0 net52
rlabel metal3 25312 26824 25312 26824 0 net53
rlabel metal2 20496 23688 20496 23688 0 net54
rlabel metal2 21336 23352 21336 23352 0 net55
rlabel metal2 40376 31556 40376 31556 0 net56
rlabel metal2 43064 34048 43064 34048 0 net57
rlabel metal2 42392 33600 42392 33600 0 net58
rlabel metal2 29400 27888 29400 27888 0 net59
rlabel metal2 56224 6552 56224 6552 0 net6
rlabel metal2 41160 4704 41160 4704 0 net60
rlabel metal2 37128 34328 37128 34328 0 net61
rlabel metal2 15176 27272 15176 27272 0 net62
rlabel metal2 14392 25032 14392 25032 0 net63
rlabel metal3 17920 23912 17920 23912 0 net64
rlabel metal2 41104 30184 41104 30184 0 net65
rlabel metal2 40208 31752 40208 31752 0 net66
rlabel metal2 38920 32424 38920 32424 0 net67
rlabel metal3 41048 31416 41048 31416 0 net68
rlabel metal2 2016 29288 2016 29288 0 net7
rlabel metal2 55944 3976 55944 3976 0 net8
rlabel metal2 54320 4536 54320 4536 0 net9
rlabel metal2 24136 15848 24136 15848 0 p_shaping_I.p_shaping_I.bit_in
rlabel metal2 38024 5600 38024 5600 0 p_shaping_I.p_shaping_I.bit_in_1
rlabel metal3 42336 8232 42336 8232 0 p_shaping_I.p_shaping_I.bit_in_2
rlabel metal2 42616 5376 42616 5376 0 p_shaping_I.p_shaping_I.counter\[0\]
rlabel metal3 41888 5992 41888 5992 0 p_shaping_I.p_shaping_I.counter\[1\]
rlabel metal3 25816 24808 25816 24808 0 p_shaping_I.p_shaping_I.ctl_1
rlabel metal2 28616 32984 28616 32984 0 p_shaping_Q.p_shaping_I.bit_in
rlabel metal2 25928 32592 25928 32592 0 p_shaping_Q.p_shaping_I.bit_in_1
rlabel metal2 27720 40992 27720 40992 0 p_shaping_Q.p_shaping_I.bit_in_2
rlabel metal2 37800 34496 37800 34496 0 p_shaping_Q.p_shaping_I.counter\[0\]
rlabel metal3 34104 40936 34104 40936 0 p_shaping_Q.p_shaping_I.counter\[1\]
rlabel metal2 32088 32984 32088 32984 0 p_shaping_Q.p_shaping_I.ctl_1
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
